magic
tech sky130A
magscale 1 2
timestamp 1682239706
<< viali >>
rect 2329 32521 2363 32555
rect 4353 32521 4387 32555
rect 5181 32521 5215 32555
rect 6009 32521 6043 32555
rect 6929 32521 6963 32555
rect 7757 32521 7791 32555
rect 8585 32521 8619 32555
rect 9505 32521 9539 32555
rect 10333 32521 10367 32555
rect 11161 32521 11195 32555
rect 2145 32385 2179 32419
rect 7757 32385 7791 32419
rect 8585 32385 8619 32419
rect 11897 32385 11931 32419
rect 14289 32385 14323 32419
rect 14473 32385 14507 32419
rect 15189 32385 15223 32419
rect 17049 32385 17083 32419
rect 17765 32385 17799 32419
rect 20065 32385 20099 32419
rect 22017 32385 22051 32419
rect 22201 32385 22235 32419
rect 22661 32385 22695 32419
rect 22845 32385 22879 32419
rect 23489 32385 23523 32419
rect 25881 32385 25915 32419
rect 26065 32385 26099 32419
rect 27353 32385 27387 32419
rect 27813 32385 27847 32419
rect 2421 32317 2455 32351
rect 3065 32317 3099 32351
rect 3433 32317 3467 32351
rect 3985 32317 4019 32351
rect 4813 32317 4847 32351
rect 5641 32317 5675 32351
rect 6561 32317 6595 32351
rect 7389 32317 7423 32351
rect 8217 32317 8251 32351
rect 9137 32317 9171 32351
rect 9965 32317 9999 32351
rect 10793 32317 10827 32351
rect 12357 32317 12391 32351
rect 13277 32317 13311 32351
rect 14933 32317 14967 32351
rect 17509 32317 17543 32351
rect 19809 32317 19843 32351
rect 25421 32317 25455 32351
rect 1869 32249 1903 32283
rect 4353 32249 4387 32283
rect 5181 32249 5215 32283
rect 6009 32249 6043 32283
rect 6929 32249 6963 32283
rect 9505 32249 9539 32283
rect 10333 32249 10367 32283
rect 11161 32249 11195 32283
rect 12633 32249 12667 32283
rect 13553 32249 13587 32283
rect 16865 32249 16899 32283
rect 2881 32181 2915 32215
rect 3433 32181 3467 32215
rect 11713 32181 11747 32215
rect 12817 32181 12851 32215
rect 13737 32181 13771 32215
rect 16313 32181 16347 32215
rect 18889 32181 18923 32215
rect 21189 32181 21223 32215
rect 23305 32181 23339 32215
rect 24777 32181 24811 32215
rect 27997 32181 28031 32215
rect 3341 31977 3375 32011
rect 2145 31909 2179 31943
rect 4445 31909 4479 31943
rect 5273 31909 5307 31943
rect 7757 31909 7791 31943
rect 7849 31909 7883 31943
rect 8493 31909 8527 31943
rect 9965 31909 9999 31943
rect 12633 31909 12667 31943
rect 13553 31909 13587 31943
rect 17877 31909 17911 31943
rect 18705 31909 18739 31943
rect 20821 31909 20855 31943
rect 22937 31909 22971 31943
rect 25973 31909 26007 31943
rect 26433 31909 26467 31943
rect 27261 31909 27295 31943
rect 27721 31909 27755 31943
rect 2605 31841 2639 31875
rect 2697 31841 2731 31875
rect 13737 31841 13771 31875
rect 3249 31773 3283 31807
rect 4077 31773 4111 31807
rect 4905 31773 4939 31807
rect 5733 31773 5767 31807
rect 6101 31773 6135 31807
rect 6561 31773 6595 31807
rect 6929 31773 6963 31807
rect 7389 31773 7423 31807
rect 8309 31773 8343 31807
rect 10425 31773 10459 31807
rect 10701 31773 10735 31807
rect 12817 31773 12851 31807
rect 14289 31773 14323 31807
rect 16486 31773 16520 31807
rect 18337 31773 18371 31807
rect 19441 31773 19475 31807
rect 21557 31773 21591 31807
rect 23581 31773 23615 31807
rect 24593 31773 24627 31807
rect 26433 31773 26467 31807
rect 26617 31773 26651 31807
rect 27721 31773 27755 31807
rect 27905 31773 27939 31807
rect 9597 31705 9631 31739
rect 10946 31705 10980 31739
rect 13277 31705 13311 31739
rect 16764 31705 16798 31739
rect 19686 31705 19720 31739
rect 21802 31705 21836 31739
rect 24838 31705 24872 31739
rect 2605 31637 2639 31671
rect 4445 31637 4479 31671
rect 5273 31637 5307 31671
rect 6101 31637 6135 31671
rect 6929 31637 6963 31671
rect 10057 31637 10091 31671
rect 12081 31637 12115 31671
rect 15577 31637 15611 31671
rect 18705 31637 18739 31671
rect 23397 31637 23431 31671
rect 2053 31433 2087 31467
rect 5181 31433 5215 31467
rect 6009 31433 6043 31467
rect 7021 31433 7055 31467
rect 7849 31433 7883 31467
rect 8677 31433 8711 31467
rect 10977 31433 11011 31467
rect 16865 31433 16899 31467
rect 24501 31433 24535 31467
rect 27169 31433 27203 31467
rect 15200 31365 15234 31399
rect 2513 31297 2547 31331
rect 4813 31297 4847 31331
rect 5181 31297 5215 31331
rect 6009 31297 6043 31331
rect 7021 31297 7055 31331
rect 9404 31297 9438 31331
rect 11161 31297 11195 31331
rect 12633 31297 12667 31331
rect 13360 31297 13394 31331
rect 17049 31297 17083 31331
rect 17765 31297 17799 31331
rect 19605 31297 19639 31331
rect 21373 31297 21407 31331
rect 22273 31297 22307 31331
rect 23857 31297 23891 31331
rect 24041 31297 24075 31331
rect 24685 31297 24719 31331
rect 25329 31297 25363 31331
rect 26433 31297 26467 31331
rect 26617 31297 26651 31331
rect 27353 31297 27387 31331
rect 1685 31229 1719 31263
rect 5641 31229 5675 31263
rect 6653 31229 6687 31263
rect 7481 31229 7515 31263
rect 8309 31229 8343 31263
rect 9137 31229 9171 31263
rect 12265 31229 12299 31263
rect 13093 31229 13127 31263
rect 14933 31229 14967 31263
rect 17509 31229 17543 31263
rect 19349 31229 19383 31263
rect 22017 31229 22051 31263
rect 27997 31229 28031 31263
rect 2053 31161 2087 31195
rect 7849 31161 7883 31195
rect 8677 31161 8711 31195
rect 20729 31161 20763 31195
rect 25973 31161 26007 31195
rect 3801 31093 3835 31127
rect 10517 31093 10551 31127
rect 12633 31093 12667 31127
rect 14473 31093 14507 31127
rect 16313 31093 16347 31127
rect 18889 31093 18923 31127
rect 21189 31093 21223 31127
rect 23397 31093 23431 31127
rect 9965 30889 9999 30923
rect 13737 30889 13771 30923
rect 15669 30889 15703 30923
rect 18429 30889 18463 30923
rect 20913 30889 20947 30923
rect 25421 30889 25455 30923
rect 26709 30889 26743 30923
rect 4077 30821 4111 30855
rect 6101 30821 6135 30855
rect 6929 30821 6963 30855
rect 16497 30821 16531 30855
rect 17325 30821 17359 30855
rect 17785 30821 17819 30855
rect 27813 30821 27847 30855
rect 3341 30753 3375 30787
rect 7849 30753 7883 30787
rect 9597 30753 9631 30787
rect 12173 30753 12207 30787
rect 13737 30753 13771 30787
rect 14289 30753 14323 30787
rect 16129 30753 16163 30787
rect 21373 30753 21407 30787
rect 24041 30753 24075 30787
rect 27307 30753 27341 30787
rect 1593 30685 1627 30719
rect 4629 30685 4663 30719
rect 5733 30685 5767 30719
rect 6561 30685 6595 30719
rect 7573 30685 7607 30719
rect 9965 30685 9999 30719
rect 12633 30685 12667 30719
rect 13369 30685 13403 30719
rect 16957 30685 16991 30719
rect 17969 30685 18003 30719
rect 18613 30685 18647 30719
rect 19533 30685 19567 30719
rect 21629 30685 21663 30719
rect 23213 30685 23247 30719
rect 23397 30685 23431 30719
rect 24593 30685 24627 30719
rect 24777 30685 24811 30719
rect 26065 30685 26099 30719
rect 27204 30685 27238 30719
rect 27997 30685 28031 30719
rect 4353 30617 4387 30651
rect 10425 30617 10459 30651
rect 14556 30617 14590 30651
rect 19800 30617 19834 30651
rect 4537 30549 4571 30583
rect 6101 30549 6135 30583
rect 6929 30549 6963 30583
rect 12817 30549 12851 30583
rect 16497 30549 16531 30583
rect 17325 30549 17359 30583
rect 22753 30549 22787 30583
rect 5273 30345 5307 30379
rect 12081 30345 12115 30379
rect 15853 30345 15887 30379
rect 20729 30345 20763 30379
rect 2145 30277 2179 30311
rect 7205 30277 7239 30311
rect 10048 30277 10082 30311
rect 17132 30277 17166 30311
rect 27307 30277 27341 30311
rect 1961 30209 1995 30243
rect 2053 30209 2087 30243
rect 2237 30209 2271 30243
rect 2421 30209 2455 30243
rect 2881 30209 2915 30243
rect 5273 30209 5307 30243
rect 6745 30209 6779 30243
rect 8125 30209 8159 30243
rect 12081 30209 12115 30243
rect 12725 30209 12759 30243
rect 12992 30209 13026 30243
rect 20269 30209 20303 30243
rect 20913 30209 20947 30243
rect 22017 30209 22051 30243
rect 22201 30209 22235 30243
rect 23101 30209 23135 30243
rect 24685 30209 24719 30243
rect 24869 30209 24903 30243
rect 25329 30209 25363 30243
rect 25513 30209 25547 30243
rect 25963 30209 25997 30243
rect 26157 30209 26191 30243
rect 27204 30209 27238 30243
rect 27997 30209 28031 30243
rect 4629 30141 4663 30175
rect 5089 30141 5123 30175
rect 5641 30141 5675 30175
rect 7665 30141 7699 30175
rect 8401 30141 8435 30175
rect 9781 30141 9815 30175
rect 11713 30141 11747 30175
rect 14565 30141 14599 30175
rect 15025 30141 15059 30175
rect 15485 30141 15519 30175
rect 16865 30141 16899 30175
rect 18797 30141 18831 30175
rect 19073 30141 19107 30175
rect 22845 30141 22879 30175
rect 7573 30073 7607 30107
rect 14933 30073 14967 30107
rect 15853 30073 15887 30107
rect 1777 30005 1811 30039
rect 6561 30005 6595 30039
rect 11161 30005 11195 30039
rect 14105 30005 14139 30039
rect 18245 30005 18279 30039
rect 20085 30005 20119 30039
rect 24225 30005 24259 30039
rect 27813 30005 27847 30039
rect 2789 29801 2823 29835
rect 13093 29801 13127 29835
rect 13553 29801 13587 29835
rect 20821 29801 20855 29835
rect 23213 29801 23247 29835
rect 27629 29801 27663 29835
rect 4445 29733 4479 29767
rect 5273 29733 5307 29767
rect 6101 29733 6135 29767
rect 7757 29733 7791 29767
rect 14565 29733 14599 29767
rect 26985 29733 27019 29767
rect 2145 29665 2179 29699
rect 5733 29665 5767 29699
rect 7389 29665 7423 29699
rect 21833 29665 21867 29699
rect 2421 29597 2455 29631
rect 4077 29597 4111 29631
rect 4905 29597 4939 29631
rect 6561 29597 6595 29631
rect 6929 29597 6963 29631
rect 8217 29597 8251 29631
rect 8585 29597 8619 29631
rect 9597 29597 9631 29631
rect 11713 29597 11747 29631
rect 13737 29597 13771 29631
rect 15025 29597 15059 29631
rect 15281 29597 15315 29631
rect 17141 29597 17175 29631
rect 19441 29597 19475 29631
rect 19697 29597 19731 29631
rect 22089 29597 22123 29631
rect 23673 29597 23707 29631
rect 23857 29597 23891 29631
rect 25145 29597 25179 29631
rect 27169 29597 27203 29631
rect 27813 29597 27847 29631
rect 2605 29529 2639 29563
rect 9864 29529 9898 29563
rect 11980 29529 12014 29563
rect 14381 29529 14415 29563
rect 17386 29529 17420 29563
rect 25390 29529 25424 29563
rect 2513 29461 2547 29495
rect 4445 29461 4479 29495
rect 5273 29461 5307 29495
rect 6101 29461 6135 29495
rect 6929 29461 6963 29495
rect 7757 29461 7791 29495
rect 8585 29461 8619 29495
rect 10977 29461 11011 29495
rect 16405 29461 16439 29495
rect 18521 29461 18555 29495
rect 26525 29461 26559 29495
rect 2881 29257 2915 29291
rect 5089 29257 5123 29291
rect 6009 29257 6043 29291
rect 7665 29257 7699 29291
rect 8585 29257 8619 29291
rect 9413 29257 9447 29291
rect 11713 29257 11747 29291
rect 12725 29257 12759 29291
rect 13553 29257 13587 29291
rect 14749 29257 14783 29291
rect 16221 29257 16255 29291
rect 19533 29257 19567 29291
rect 21465 29257 21499 29291
rect 22017 29257 22051 29291
rect 27307 29257 27341 29291
rect 3801 29189 3835 29223
rect 3985 29189 4019 29223
rect 17570 29189 17604 29223
rect 19165 29189 19199 29223
rect 25881 29189 25915 29223
rect 1593 29121 1627 29155
rect 5089 29121 5123 29155
rect 6009 29121 6043 29155
rect 6745 29121 6779 29155
rect 7021 29121 7055 29155
rect 7481 29121 7515 29155
rect 8217 29121 8251 29155
rect 9045 29121 9079 29155
rect 11897 29121 11931 29155
rect 12725 29121 12759 29155
rect 13553 29121 13587 29155
rect 15761 29121 15795 29155
rect 17325 29121 17359 29155
rect 19349 29121 19383 29155
rect 20085 29121 20119 29155
rect 20352 29121 20386 29155
rect 22201 29121 22235 29155
rect 22661 29121 22695 29155
rect 22845 29121 22879 29155
rect 24205 29121 24239 29155
rect 25789 29121 25823 29155
rect 25973 29121 26007 29155
rect 26433 29121 26467 29155
rect 26617 29121 26651 29155
rect 27204 29121 27238 29155
rect 27997 29121 28031 29155
rect 4721 29053 4755 29087
rect 5641 29053 5675 29087
rect 6561 29053 6595 29087
rect 10241 29053 10275 29087
rect 12357 29053 12391 29087
rect 13185 29053 13219 29087
rect 14289 29053 14323 29087
rect 23949 29053 23983 29087
rect 4169 28985 4203 29019
rect 6929 28985 6963 29019
rect 8585 28985 8619 29019
rect 9413 28985 9447 29019
rect 10517 28985 10551 29019
rect 10701 28985 10735 29019
rect 14657 28985 14691 29019
rect 16129 28985 16163 29019
rect 25329 28985 25363 29019
rect 27813 28985 27847 29019
rect 3985 28917 4019 28951
rect 18705 28917 18739 28951
rect 23489 28917 23523 28951
rect 26433 28917 26467 28951
rect 15209 28713 15243 28747
rect 17141 28713 17175 28747
rect 21465 28713 21499 28747
rect 22293 28713 22327 28747
rect 9321 28645 9355 28679
rect 11069 28645 11103 28679
rect 11897 28645 11931 28679
rect 15025 28645 15059 28679
rect 18797 28645 18831 28679
rect 23581 28645 23615 28679
rect 25973 28645 26007 28679
rect 8033 28577 8067 28611
rect 13185 28577 13219 28611
rect 26893 28577 26927 28611
rect 1777 28509 1811 28543
rect 2033 28509 2067 28543
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 5273 28509 5307 28543
rect 6837 28509 6871 28543
rect 7481 28509 7515 28543
rect 7665 28509 7699 28543
rect 9137 28509 9171 28543
rect 9873 28509 9907 28543
rect 10241 28509 10275 28543
rect 10701 28509 10735 28543
rect 11529 28509 11563 28543
rect 12357 28509 12391 28543
rect 12725 28509 12759 28543
rect 13553 28509 13587 28543
rect 15669 28509 15703 28543
rect 19625 28509 19659 28543
rect 19881 28509 19915 28543
rect 21649 28509 21683 28543
rect 22937 28509 22971 28543
rect 24593 28509 24627 28543
rect 24849 28509 24883 28543
rect 14749 28441 14783 28475
rect 18429 28441 18463 28475
rect 27138 28441 27172 28475
rect 3157 28373 3191 28407
rect 4261 28373 4295 28407
rect 7665 28373 7699 28407
rect 10241 28373 10275 28407
rect 11069 28373 11103 28407
rect 11897 28373 11931 28407
rect 12725 28373 12759 28407
rect 13553 28373 13587 28407
rect 18889 28373 18923 28407
rect 21005 28373 21039 28407
rect 28273 28373 28307 28407
rect 4997 28169 5031 28203
rect 7205 28169 7239 28203
rect 8125 28169 8159 28203
rect 9137 28169 9171 28203
rect 11897 28169 11931 28203
rect 14473 28169 14507 28203
rect 16313 28169 16347 28203
rect 24777 28169 24811 28203
rect 25421 28169 25455 28203
rect 26157 28169 26191 28203
rect 27951 28169 27985 28203
rect 8217 28101 8251 28135
rect 11805 28101 11839 28135
rect 1777 28033 1811 28067
rect 1869 28033 1903 28067
rect 2605 28033 2639 28067
rect 2872 28033 2906 28067
rect 4997 28033 5031 28067
rect 5641 28033 5675 28067
rect 7849 28033 7883 28067
rect 8309 28033 8343 28067
rect 9853 28033 9887 28067
rect 12449 28033 12483 28067
rect 14105 28033 14139 28067
rect 14289 28033 14323 28067
rect 14933 28033 14967 28067
rect 15117 28033 15151 28067
rect 15209 28033 15243 28067
rect 15301 28033 15335 28067
rect 17121 28033 17155 28067
rect 18705 28033 18739 28067
rect 18889 28033 18923 28067
rect 18981 28033 19015 28067
rect 19073 28033 19107 28067
rect 20341 28033 20375 28067
rect 22549 28033 22583 28067
rect 24317 28033 24351 28067
rect 24961 28033 24995 28067
rect 25605 28033 25639 28067
rect 26065 28033 26099 28067
rect 27169 28033 27203 28067
rect 27848 28033 27882 28067
rect 2053 27965 2087 27999
rect 4629 27965 4663 27999
rect 5457 27965 5491 27999
rect 6009 27965 6043 27999
rect 6745 27965 6779 27999
rect 8769 27965 8803 27999
rect 9597 27965 9631 27999
rect 12725 27965 12759 27999
rect 15945 27965 15979 27999
rect 16313 27965 16347 27999
rect 16865 27965 16899 27999
rect 20085 27965 20119 27999
rect 22293 27965 22327 27999
rect 5917 27897 5951 27931
rect 7113 27897 7147 27931
rect 9137 27897 9171 27931
rect 18245 27897 18279 27931
rect 3985 27829 4019 27863
rect 10977 27829 11011 27863
rect 15485 27829 15519 27863
rect 19257 27829 19291 27863
rect 21465 27829 21499 27863
rect 23673 27829 23707 27863
rect 27353 27829 27387 27863
rect 4077 27557 4111 27591
rect 5641 27557 5675 27591
rect 7297 27557 7331 27591
rect 12725 27557 12759 27591
rect 14933 27557 14967 27591
rect 18429 27557 18463 27591
rect 20085 27557 20119 27591
rect 6469 27489 6503 27523
rect 6929 27489 6963 27523
rect 7757 27489 7791 27523
rect 9597 27489 9631 27523
rect 15761 27489 15795 27523
rect 17141 27489 17175 27523
rect 19625 27489 19659 27523
rect 2053 27421 2087 27455
rect 3985 27421 4019 27455
rect 4261 27421 4295 27455
rect 4537 27421 4571 27455
rect 4813 27421 4847 27455
rect 5273 27421 5307 27455
rect 6101 27421 6135 27455
rect 6285 27421 6319 27455
rect 8033 27421 8067 27455
rect 9965 27421 9999 27455
rect 10425 27421 10459 27455
rect 12357 27421 12391 27455
rect 13185 27421 13219 27455
rect 13553 27421 13587 27455
rect 14749 27421 14783 27455
rect 15393 27421 15427 27455
rect 16405 27421 16439 27455
rect 17509 27421 17543 27455
rect 18061 27421 18095 27455
rect 20269 27421 20303 27455
rect 20913 27421 20947 27455
rect 21373 27421 21407 27455
rect 22017 27421 22051 27455
rect 22661 27421 22695 27455
rect 24593 27421 24627 27455
rect 26985 27421 27019 27455
rect 2320 27353 2354 27387
rect 10670 27353 10704 27387
rect 14565 27353 14599 27387
rect 22906 27353 22940 27387
rect 24838 27353 24872 27387
rect 27230 27353 27264 27387
rect 3433 27285 3467 27319
rect 5641 27285 5675 27319
rect 7297 27285 7331 27319
rect 9965 27285 9999 27319
rect 11805 27285 11839 27319
rect 12725 27285 12759 27319
rect 13553 27285 13587 27319
rect 15761 27285 15795 27319
rect 16221 27285 16255 27319
rect 17509 27285 17543 27319
rect 18521 27285 18555 27319
rect 20729 27285 20763 27319
rect 21557 27285 21591 27319
rect 22109 27285 22143 27319
rect 24041 27285 24075 27319
rect 25973 27285 26007 27319
rect 28365 27285 28399 27319
rect 9321 27081 9355 27115
rect 9781 27081 9815 27115
rect 10977 27081 11011 27115
rect 12725 27081 12759 27115
rect 13553 27081 13587 27115
rect 15301 27081 15335 27115
rect 16129 27081 16163 27115
rect 17877 27081 17911 27115
rect 19441 27081 19475 27115
rect 2605 27013 2639 27047
rect 7941 27013 7975 27047
rect 14933 27013 14967 27047
rect 15945 27013 15979 27047
rect 17417 27013 17451 27047
rect 22262 27013 22296 27047
rect 1777 26945 1811 26979
rect 2053 26945 2087 26979
rect 4813 26945 4847 26979
rect 4997 26945 5031 26979
rect 5733 26945 5767 26979
rect 5825 26945 5859 26979
rect 6745 26945 6779 26979
rect 7113 26945 7147 26979
rect 7757 26945 7791 26979
rect 8033 26945 8067 26979
rect 10149 26945 10183 26979
rect 11161 26945 11195 26979
rect 12357 26945 12391 26979
rect 13185 26945 13219 26979
rect 14105 26945 14139 26979
rect 14289 26945 14323 26979
rect 15117 26945 15151 26979
rect 15761 26945 15795 26979
rect 17049 26945 17083 26979
rect 17233 26945 17267 26979
rect 18061 26945 18095 26979
rect 19617 26945 19651 26979
rect 20453 26945 20487 26979
rect 21097 26945 21131 26979
rect 24041 26945 24075 26979
rect 24501 26945 24535 26979
rect 25493 26945 25527 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 27813 26945 27847 26979
rect 27997 26945 28031 26979
rect 2145 26877 2179 26911
rect 6561 26877 6595 26911
rect 8953 26877 8987 26911
rect 10241 26877 10275 26911
rect 10333 26877 10367 26911
rect 11713 26877 11747 26911
rect 18521 26877 18555 26911
rect 18981 26877 19015 26911
rect 22017 26877 22051 26911
rect 25237 26877 25271 26911
rect 4077 26809 4111 26843
rect 5089 26809 5123 26843
rect 5917 26809 5951 26843
rect 7021 26809 7055 26843
rect 9321 26809 9355 26843
rect 12725 26809 12759 26843
rect 13553 26809 13587 26843
rect 14473 26809 14507 26843
rect 18797 26809 18831 26843
rect 7573 26741 7607 26775
rect 20269 26741 20303 26775
rect 20913 26741 20947 26775
rect 23397 26741 23431 26775
rect 23857 26741 23891 26775
rect 24593 26741 24627 26775
rect 26617 26741 26651 26775
rect 7573 26537 7607 26571
rect 11989 26537 12023 26571
rect 17877 26537 17911 26571
rect 18889 26537 18923 26571
rect 8585 26469 8619 26503
rect 10701 26469 10735 26503
rect 13645 26469 13679 26503
rect 18797 26469 18831 26503
rect 3433 26401 3467 26435
rect 4169 26401 4203 26435
rect 4813 26401 4847 26435
rect 5641 26401 5675 26435
rect 7113 26401 7147 26435
rect 8217 26401 8251 26435
rect 9137 26401 9171 26435
rect 11989 26401 12023 26435
rect 12817 26401 12851 26435
rect 13277 26401 13311 26435
rect 25145 26401 25179 26435
rect 3985 26333 4019 26367
rect 4537 26333 4571 26367
rect 5273 26333 5307 26367
rect 5457 26333 5491 26367
rect 6837 26333 6871 26367
rect 7021 26333 7055 26367
rect 7757 26333 7791 26367
rect 9505 26333 9539 26367
rect 10149 26333 10183 26367
rect 10425 26333 10459 26367
rect 10517 26333 10551 26367
rect 11621 26333 11655 26367
rect 12633 26333 12667 26367
rect 14841 26333 14875 26367
rect 14934 26333 14968 26367
rect 15209 26333 15243 26367
rect 15347 26333 15381 26367
rect 16497 26333 16531 26367
rect 19441 26333 19475 26367
rect 21281 26333 21315 26367
rect 23121 26333 23155 26367
rect 23305 26333 23339 26367
rect 23765 26333 23799 26367
rect 23949 26333 23983 26367
rect 26985 26333 27019 26367
rect 27241 26333 27275 26367
rect 1685 26265 1719 26299
rect 4077 26265 4111 26299
rect 6653 26265 6687 26299
rect 10333 26265 10367 26299
rect 12449 26265 12483 26299
rect 15117 26265 15151 26299
rect 16742 26265 16776 26299
rect 18429 26265 18463 26299
rect 19686 26265 19720 26299
rect 21526 26265 21560 26299
rect 23213 26265 23247 26299
rect 23857 26265 23891 26299
rect 25390 26265 25424 26299
rect 8585 26197 8619 26231
rect 9505 26197 9539 26231
rect 13645 26197 13679 26231
rect 15485 26197 15519 26231
rect 20821 26197 20855 26231
rect 22661 26197 22695 26231
rect 26525 26197 26559 26231
rect 28365 26197 28399 26231
rect 2421 25993 2455 26027
rect 8125 25993 8159 26027
rect 9413 25993 9447 26027
rect 9781 25993 9815 26027
rect 9873 25993 9907 26027
rect 11069 25993 11103 26027
rect 19625 25993 19659 26027
rect 21189 25993 21223 26027
rect 3433 25925 3467 25959
rect 6929 25925 6963 25959
rect 15178 25925 15212 25959
rect 16865 25925 16899 25959
rect 17233 25925 17267 25959
rect 22273 25925 22307 25959
rect 2421 25857 2455 25891
rect 2605 25857 2639 25891
rect 5641 25857 5675 25891
rect 5917 25857 5951 25891
rect 7113 25857 7147 25891
rect 7757 25857 7791 25891
rect 8769 25857 8803 25891
rect 10701 25857 10735 25891
rect 10885 25857 10919 25891
rect 11805 25857 11839 25891
rect 12716 25857 12750 25891
rect 14473 25857 14507 25891
rect 14933 25857 14967 25891
rect 17049 25857 17083 25891
rect 19165 25857 19199 25891
rect 19809 25857 19843 25891
rect 20453 25857 20487 25891
rect 21373 25857 21407 25891
rect 24113 25857 24147 25891
rect 25697 25857 25731 25891
rect 2145 25789 2179 25823
rect 2973 25789 3007 25823
rect 8585 25789 8619 25823
rect 9965 25789 9999 25823
rect 11989 25789 12023 25823
rect 12449 25789 12483 25823
rect 18061 25789 18095 25823
rect 18521 25789 18555 25823
rect 22017 25789 22051 25823
rect 23857 25789 23891 25823
rect 4721 25721 4755 25755
rect 5917 25721 5951 25755
rect 8125 25721 8159 25755
rect 18429 25721 18463 25755
rect 20269 25721 20303 25755
rect 25881 25721 25915 25755
rect 7297 25653 7331 25687
rect 8953 25653 8987 25687
rect 13829 25653 13863 25687
rect 14289 25653 14323 25687
rect 16313 25653 16347 25687
rect 18981 25653 19015 25687
rect 23397 25653 23431 25687
rect 25237 25653 25271 25687
rect 3341 25449 3375 25483
rect 8401 25449 8435 25483
rect 9873 25449 9907 25483
rect 15025 25449 15059 25483
rect 17877 25449 17911 25483
rect 19809 25449 19843 25483
rect 20269 25449 20303 25483
rect 21189 25449 21223 25483
rect 22017 25449 22051 25483
rect 22753 25449 22787 25483
rect 23305 25449 23339 25483
rect 6009 25381 6043 25415
rect 18705 25381 18739 25415
rect 8033 25313 8067 25347
rect 10517 25313 10551 25347
rect 13645 25313 13679 25347
rect 1961 25245 1995 25279
rect 2217 25245 2251 25279
rect 3985 25245 4019 25279
rect 6193 25245 6227 25279
rect 6285 25245 6319 25279
rect 6495 25245 6529 25279
rect 6653 25245 6687 25279
rect 7205 25245 7239 25279
rect 9229 25245 9263 25279
rect 9413 25245 9447 25279
rect 11437 25245 11471 25279
rect 13461 25245 13495 25279
rect 15853 25245 15887 25279
rect 16129 25245 16163 25279
rect 18429 25245 18463 25279
rect 18521 25245 18555 25279
rect 20453 25245 20487 25279
rect 21373 25245 21407 25279
rect 21925 25245 21959 25279
rect 22569 25245 22603 25279
rect 23489 25245 23523 25279
rect 24593 25245 24627 25279
rect 24777 25245 24811 25279
rect 26065 25245 26099 25279
rect 4230 25177 4264 25211
rect 6377 25177 6411 25211
rect 7573 25177 7607 25211
rect 10333 25177 10367 25211
rect 11682 25177 11716 25211
rect 13277 25177 13311 25211
rect 14841 25177 14875 25211
rect 17509 25177 17543 25211
rect 17693 25177 17727 25211
rect 19441 25177 19475 25211
rect 19625 25177 19659 25211
rect 26332 25177 26366 25211
rect 5365 25109 5399 25143
rect 8401 25109 8435 25143
rect 8585 25109 8619 25143
rect 10241 25109 10275 25143
rect 12817 25109 12851 25143
rect 15041 25109 15075 25143
rect 15209 25109 15243 25143
rect 24685 25109 24719 25143
rect 27445 25109 27479 25143
rect 1869 24905 1903 24939
rect 5089 24905 5123 24939
rect 6929 24905 6963 24939
rect 9229 24905 9263 24939
rect 11161 24905 11195 24939
rect 19901 24905 19935 24939
rect 5181 24837 5215 24871
rect 6561 24837 6595 24871
rect 8585 24837 8619 24871
rect 12081 24837 12115 24871
rect 17417 24837 17451 24871
rect 25482 24837 25516 24871
rect 6791 24803 6825 24837
rect 17647 24803 17681 24837
rect 1593 24769 1627 24803
rect 1869 24769 1903 24803
rect 2872 24769 2906 24803
rect 4905 24769 4939 24803
rect 5733 24769 5767 24803
rect 5825 24769 5859 24803
rect 7573 24769 7607 24803
rect 8401 24769 8435 24803
rect 9413 24769 9447 24803
rect 9873 24769 9907 24803
rect 10333 24769 10367 24803
rect 10609 24769 10643 24803
rect 12173 24769 12207 24803
rect 13461 24769 13495 24803
rect 13717 24769 13751 24803
rect 15669 24769 15703 24803
rect 15762 24769 15796 24803
rect 15945 24769 15979 24803
rect 16037 24769 16071 24803
rect 16134 24769 16168 24803
rect 20545 24769 20579 24803
rect 21189 24769 21223 24803
rect 22273 24769 22307 24803
rect 24041 24769 24075 24803
rect 24685 24769 24719 24803
rect 25237 24769 25271 24803
rect 2605 24701 2639 24735
rect 6009 24701 6043 24735
rect 12357 24701 12391 24735
rect 18245 24701 18279 24735
rect 18705 24701 18739 24735
rect 19441 24701 19475 24735
rect 22017 24701 22051 24735
rect 3985 24633 4019 24667
rect 7849 24633 7883 24667
rect 18613 24633 18647 24667
rect 19717 24633 19751 24667
rect 20361 24633 20395 24667
rect 23857 24633 23891 24667
rect 4629 24565 4663 24599
rect 5917 24565 5951 24599
rect 6745 24565 6779 24599
rect 8769 24565 8803 24599
rect 11713 24565 11747 24599
rect 14841 24565 14875 24599
rect 16313 24565 16347 24599
rect 17601 24565 17635 24599
rect 17785 24565 17819 24599
rect 21005 24565 21039 24599
rect 23397 24565 23431 24599
rect 24501 24565 24535 24599
rect 26617 24565 26651 24599
rect 4077 24361 4111 24395
rect 6929 24361 6963 24395
rect 7757 24361 7791 24395
rect 8401 24361 8435 24395
rect 17785 24361 17819 24395
rect 18705 24361 18739 24395
rect 20453 24361 20487 24395
rect 11713 24293 11747 24327
rect 13737 24293 13771 24327
rect 20269 24293 20303 24327
rect 21281 24293 21315 24327
rect 23673 24293 23707 24327
rect 5457 24225 5491 24259
rect 14657 24225 14691 24259
rect 19993 24225 20027 24259
rect 20913 24225 20947 24259
rect 22293 24225 22327 24259
rect 26433 24225 26467 24259
rect 2053 24157 2087 24191
rect 2309 24157 2343 24191
rect 4629 24157 4663 24191
rect 5181 24157 5215 24191
rect 5365 24157 5399 24191
rect 5549 24157 5583 24191
rect 5688 24157 5722 24191
rect 7389 24157 7423 24191
rect 7573 24157 7607 24191
rect 9229 24157 9263 24191
rect 9413 24157 9447 24191
rect 10425 24157 10459 24191
rect 10701 24157 10735 24191
rect 11161 24157 11195 24191
rect 12173 24157 12207 24191
rect 12266 24157 12300 24191
rect 12449 24157 12483 24191
rect 12638 24157 12672 24191
rect 13553 24157 13587 24191
rect 14565 24157 14599 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15025 24157 15059 24191
rect 15669 24157 15703 24191
rect 17877 24157 17911 24191
rect 17969 24157 18003 24191
rect 18061 24157 18095 24191
rect 18245 24157 18279 24191
rect 18889 24157 18923 24191
rect 24593 24157 24627 24191
rect 4353 24089 4387 24123
rect 4537 24089 4571 24123
rect 6561 24089 6595 24123
rect 6745 24089 6779 24123
rect 8309 24089 8343 24123
rect 9597 24089 9631 24123
rect 12541 24089 12575 24123
rect 13369 24089 13403 24123
rect 15914 24089 15948 24123
rect 17509 24089 17543 24123
rect 22560 24089 22594 24123
rect 24860 24089 24894 24123
rect 26678 24089 26712 24123
rect 3433 24021 3467 24055
rect 5917 24021 5951 24055
rect 12817 24021 12851 24055
rect 14289 24021 14323 24055
rect 17049 24021 17083 24055
rect 21373 24021 21407 24055
rect 25973 24021 26007 24055
rect 27813 24021 27847 24055
rect 1869 23817 1903 23851
rect 1961 23817 1995 23851
rect 3893 23817 3927 23851
rect 5089 23817 5123 23851
rect 5181 23817 5215 23851
rect 7849 23817 7883 23851
rect 9597 23817 9631 23851
rect 10993 23817 11027 23851
rect 11713 23817 11747 23851
rect 13369 23817 13403 23851
rect 13829 23817 13863 23851
rect 15025 23817 15059 23851
rect 15853 23817 15887 23851
rect 20453 23817 20487 23851
rect 21097 23817 21131 23851
rect 24593 23817 24627 23851
rect 1777 23749 1811 23783
rect 2605 23749 2639 23783
rect 4813 23749 4847 23783
rect 10793 23749 10827 23783
rect 14657 23749 14691 23783
rect 14873 23749 14907 23783
rect 15485 23749 15519 23783
rect 15690 23749 15724 23783
rect 16957 23749 16991 23783
rect 19165 23749 19199 23783
rect 2145 23681 2179 23715
rect 4997 23681 5031 23715
rect 5365 23681 5399 23715
rect 6009 23681 6043 23715
rect 6653 23681 6687 23715
rect 6929 23681 6963 23715
rect 7481 23681 7515 23715
rect 8879 23681 8913 23715
rect 9965 23681 9999 23715
rect 12081 23681 12115 23715
rect 13001 23681 13035 23715
rect 13185 23681 13219 23715
rect 14013 23681 14047 23715
rect 17785 23681 17819 23715
rect 18797 23681 18831 23715
rect 18981 23681 19015 23715
rect 19625 23681 19659 23715
rect 19809 23681 19843 23715
rect 20637 23681 20671 23715
rect 21281 23681 21315 23715
rect 22293 23681 22327 23715
rect 23213 23681 23247 23715
rect 23480 23681 23514 23715
rect 25493 23681 25527 23715
rect 7573 23613 7607 23647
rect 8401 23613 8435 23647
rect 8585 23613 8619 23647
rect 8978 23613 9012 23647
rect 10057 23613 10091 23647
rect 10241 23613 10275 23647
rect 12173 23613 12207 23647
rect 12357 23613 12391 23647
rect 19993 23613 20027 23647
rect 25237 23613 25271 23647
rect 1593 23545 1627 23579
rect 5825 23545 5859 23579
rect 6929 23545 6963 23579
rect 11161 23545 11195 23579
rect 17601 23545 17635 23579
rect 7665 23477 7699 23511
rect 10977 23477 11011 23511
rect 14841 23477 14875 23511
rect 15669 23477 15703 23511
rect 17049 23477 17083 23511
rect 22109 23477 22143 23511
rect 26617 23477 26651 23511
rect 2513 23273 2547 23307
rect 4077 23273 4111 23307
rect 7849 23273 7883 23307
rect 11345 23273 11379 23307
rect 13553 23273 13587 23307
rect 13737 23273 13771 23307
rect 16037 23273 16071 23307
rect 17049 23273 17083 23307
rect 17877 23273 17911 23307
rect 18889 23273 18923 23307
rect 19901 23273 19935 23307
rect 21925 23273 21959 23307
rect 22937 23273 22971 23307
rect 23489 23273 23523 23307
rect 27445 23273 27479 23307
rect 1685 23205 1719 23239
rect 6469 23205 6503 23239
rect 14657 23205 14691 23239
rect 15209 23205 15243 23239
rect 16221 23205 16255 23239
rect 19717 23205 19751 23239
rect 3065 23137 3099 23171
rect 9689 23137 9723 23171
rect 14749 23137 14783 23171
rect 1685 23069 1719 23103
rect 1961 23069 1995 23103
rect 2789 23069 2823 23103
rect 4353 23069 4387 23103
rect 4445 23069 4479 23103
rect 4537 23069 4571 23103
rect 4721 23069 4755 23103
rect 5365 23069 5399 23103
rect 5549 23069 5583 23103
rect 5641 23069 5675 23103
rect 6285 23069 6319 23103
rect 6561 23069 6595 23103
rect 7481 23069 7515 23103
rect 7849 23069 7883 23103
rect 9505 23069 9539 23103
rect 10333 23069 10367 23103
rect 10517 23069 10551 23103
rect 10701 23069 10735 23103
rect 11529 23069 11563 23103
rect 11989 23069 12023 23103
rect 12137 23069 12171 23103
rect 12454 23069 12488 23103
rect 15393 23069 15427 23103
rect 16681 23069 16715 23103
rect 16865 23069 16899 23103
rect 17509 23069 17543 23103
rect 17693 23069 17727 23103
rect 20545 23069 20579 23103
rect 22845 23069 22879 23103
rect 23673 23069 23707 23103
rect 24777 23069 24811 23103
rect 26065 23069 26099 23103
rect 2973 23001 3007 23035
rect 10609 23001 10643 23035
rect 12265 23001 12299 23035
rect 12357 23001 12391 23035
rect 13369 23001 13403 23035
rect 14289 23001 14323 23035
rect 15853 23001 15887 23035
rect 18521 23001 18555 23035
rect 18705 23001 18739 23035
rect 19441 23001 19475 23035
rect 20790 23001 20824 23035
rect 26332 23001 26366 23035
rect 1869 22933 1903 22967
rect 5181 22933 5215 22967
rect 6101 22933 6135 22967
rect 8033 22933 8067 22967
rect 9137 22933 9171 22967
rect 9597 22933 9631 22967
rect 10885 22933 10919 22967
rect 12633 22933 12667 22967
rect 13569 22933 13603 22967
rect 16053 22933 16087 22967
rect 24593 22933 24627 22967
rect 1970 22729 2004 22763
rect 4537 22729 4571 22763
rect 5089 22729 5123 22763
rect 7297 22729 7331 22763
rect 9137 22729 9171 22763
rect 10977 22729 11011 22763
rect 12909 22729 12943 22763
rect 17233 22729 17267 22763
rect 19717 22729 19751 22763
rect 21005 22729 21039 22763
rect 26617 22729 26651 22763
rect 13645 22661 13679 22695
rect 13861 22661 13895 22695
rect 17693 22661 17727 22695
rect 18705 22661 18739 22695
rect 19533 22661 19567 22695
rect 20177 22661 20211 22695
rect 20545 22661 20579 22695
rect 25482 22661 25516 22695
rect 17923 22627 17957 22661
rect 1593 22593 1627 22627
rect 2237 22593 2271 22627
rect 3525 22593 3559 22627
rect 3617 22593 3651 22627
rect 3709 22593 3743 22627
rect 3893 22593 3927 22627
rect 4353 22593 4387 22627
rect 5457 22593 5491 22627
rect 6837 22593 6871 22627
rect 8677 22593 8711 22627
rect 9597 22593 9631 22627
rect 9864 22593 9898 22627
rect 12633 22593 12667 22627
rect 13001 22593 13035 22627
rect 15577 22593 15611 22627
rect 15761 22593 15795 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 18521 22593 18555 22627
rect 18889 22593 18923 22627
rect 19349 22593 19383 22627
rect 20361 22593 20395 22627
rect 21189 22593 21223 22627
rect 22201 22593 22235 22627
rect 23009 22593 23043 22627
rect 24593 22593 24627 22627
rect 25237 22593 25271 22627
rect 5549 22525 5583 22559
rect 5641 22525 5675 22559
rect 7757 22525 7791 22559
rect 12265 22525 12299 22559
rect 15301 22525 15335 22559
rect 22753 22525 22787 22559
rect 7205 22457 7239 22491
rect 8033 22457 8067 22491
rect 9045 22457 9079 22491
rect 12725 22457 12759 22491
rect 14013 22457 14047 22491
rect 15393 22457 15427 22491
rect 15485 22457 15519 22491
rect 24685 22457 24719 22491
rect 1961 22389 1995 22423
rect 3249 22389 3283 22423
rect 8217 22389 8251 22423
rect 12541 22389 12575 22423
rect 13829 22389 13863 22423
rect 15025 22389 15059 22423
rect 17877 22389 17911 22423
rect 18061 22389 18095 22423
rect 22017 22389 22051 22423
rect 24133 22389 24167 22423
rect 3249 22185 3283 22219
rect 8125 22185 8159 22219
rect 9597 22185 9631 22219
rect 13369 22185 13403 22219
rect 17417 22185 17451 22219
rect 17601 22185 17635 22219
rect 19441 22185 19475 22219
rect 7205 22117 7239 22151
rect 14749 22117 14783 22151
rect 21925 22117 21959 22151
rect 4261 22049 4295 22083
rect 5641 22049 5675 22083
rect 9137 22049 9171 22083
rect 12725 22049 12759 22083
rect 21097 22049 21131 22083
rect 26801 22049 26835 22083
rect 1777 21981 1811 22015
rect 2001 21981 2035 22015
rect 2145 21981 2179 22015
rect 2605 21981 2639 22015
rect 2698 21981 2732 22015
rect 3111 21981 3145 22015
rect 4445 21981 4479 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 5825 21981 5859 22015
rect 6837 21981 6871 22015
rect 8309 21981 8343 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 9505 21981 9539 22015
rect 10425 21981 10459 22015
rect 10609 21981 10643 22015
rect 11069 21981 11103 22015
rect 14565 21981 14599 22015
rect 16221 21981 16255 22015
rect 16405 21981 16439 22015
rect 16497 21981 16531 22015
rect 16589 21981 16623 22015
rect 18245 21981 18279 22015
rect 18889 21981 18923 22015
rect 19625 21981 19659 22015
rect 20269 21981 20303 22015
rect 22661 21981 22695 22015
rect 24961 21981 24995 22015
rect 27057 21981 27091 22015
rect 1593 21913 1627 21947
rect 2881 21913 2915 21947
rect 2973 21913 3007 21947
rect 4629 21913 4663 21947
rect 4721 21913 4755 21947
rect 7021 21913 7055 21947
rect 12357 21913 12391 21947
rect 12541 21913 12575 21947
rect 13185 21913 13219 21947
rect 15393 21913 15427 21947
rect 17233 21913 17267 21947
rect 20729 21913 20763 21947
rect 20913 21913 20947 21947
rect 21649 21913 21683 21947
rect 22906 21913 22940 21947
rect 25206 21913 25240 21947
rect 1869 21845 1903 21879
rect 5365 21845 5399 21879
rect 9321 21845 9355 21879
rect 10609 21845 10643 21879
rect 13385 21845 13419 21879
rect 13553 21845 13587 21879
rect 15485 21845 15519 21879
rect 16773 21845 16807 21879
rect 17433 21845 17467 21879
rect 18061 21845 18095 21879
rect 18705 21845 18739 21879
rect 20085 21845 20119 21879
rect 22109 21845 22143 21879
rect 24041 21845 24075 21879
rect 26341 21845 26375 21879
rect 28181 21845 28215 21879
rect 3801 21641 3835 21675
rect 4997 21641 5031 21675
rect 7941 21641 7975 21675
rect 10425 21641 10459 21675
rect 12725 21641 12759 21675
rect 14749 21641 14783 21675
rect 15853 21641 15887 21675
rect 19717 21641 19751 21675
rect 20637 21641 20671 21675
rect 22477 21641 22511 21675
rect 22937 21641 22971 21675
rect 7849 21573 7883 21607
rect 10057 21573 10091 21607
rect 10257 21573 10291 21607
rect 11989 21573 12023 21607
rect 16865 21573 16899 21607
rect 17065 21573 17099 21607
rect 17693 21573 17727 21607
rect 17893 21573 17927 21607
rect 18521 21573 18555 21607
rect 18721 21573 18755 21607
rect 19533 21573 19567 21607
rect 23940 21573 23974 21607
rect 2053 21505 2087 21539
rect 2237 21505 2271 21539
rect 2513 21505 2547 21539
rect 3065 21505 3099 21539
rect 4169 21505 4203 21539
rect 4261 21505 4295 21539
rect 5273 21505 5307 21539
rect 5365 21505 5399 21539
rect 5457 21505 5491 21539
rect 5641 21505 5675 21539
rect 6929 21505 6963 21539
rect 7113 21505 7147 21539
rect 9045 21505 9079 21539
rect 10885 21505 10919 21539
rect 11713 21505 11747 21539
rect 11897 21505 11931 21539
rect 12081 21505 12115 21539
rect 12909 21505 12943 21539
rect 13625 21505 13659 21539
rect 15945 21505 15979 21539
rect 19349 21505 19383 21539
rect 20269 21505 20303 21539
rect 20453 21505 20487 21539
rect 21281 21505 21315 21539
rect 23121 21505 23155 21539
rect 25697 21505 25731 21539
rect 1593 21437 1627 21471
rect 2697 21437 2731 21471
rect 3985 21437 4019 21471
rect 9505 21437 9539 21471
rect 13369 21437 13403 21471
rect 15577 21437 15611 21471
rect 22017 21437 22051 21471
rect 23673 21437 23707 21471
rect 7297 21369 7331 21403
rect 8769 21369 8803 21403
rect 9413 21369 9447 21403
rect 15485 21369 15519 21403
rect 15669 21369 15703 21403
rect 17233 21369 17267 21403
rect 18061 21369 18095 21403
rect 21097 21369 21131 21403
rect 22293 21369 22327 21403
rect 10241 21301 10275 21335
rect 11069 21301 11103 21335
rect 12265 21301 12299 21335
rect 15209 21301 15243 21335
rect 17049 21301 17083 21335
rect 17877 21301 17911 21335
rect 18705 21301 18739 21335
rect 18889 21301 18923 21335
rect 25053 21301 25087 21335
rect 25513 21301 25547 21335
rect 2237 21097 2271 21131
rect 3433 21097 3467 21131
rect 5457 21097 5491 21131
rect 6009 21097 6043 21131
rect 7757 21097 7791 21131
rect 9597 21097 9631 21131
rect 10793 21097 10827 21131
rect 13369 21097 13403 21131
rect 14565 21097 14599 21131
rect 16497 21097 16531 21131
rect 17601 21097 17635 21131
rect 18705 21097 18739 21131
rect 21741 21097 21775 21131
rect 22201 21097 22235 21131
rect 23305 21097 23339 21131
rect 4353 21029 4387 21063
rect 6561 21029 6595 21063
rect 7113 21029 7147 21063
rect 11805 21029 11839 21063
rect 12633 21029 12667 21063
rect 15485 21029 15519 21063
rect 23121 21029 23155 21063
rect 3985 20961 4019 20995
rect 6653 20961 6687 20995
rect 10149 20961 10183 20995
rect 20913 20961 20947 20995
rect 24593 20961 24627 20995
rect 1593 20893 1627 20927
rect 1686 20893 1720 20927
rect 1869 20893 1903 20927
rect 2058 20893 2092 20927
rect 2789 20893 2823 20927
rect 2937 20893 2971 20927
rect 3254 20893 3288 20927
rect 4169 20893 4203 20927
rect 4445 20893 4479 20927
rect 5273 20893 5307 20927
rect 6134 20893 6168 20927
rect 7297 20893 7331 20927
rect 7941 20893 7975 20927
rect 8585 20893 8619 20927
rect 10977 20893 11011 20927
rect 11621 20893 11655 20927
rect 12357 20893 12391 20927
rect 12449 20893 12483 20927
rect 16129 20893 16163 20927
rect 16313 20893 16347 20927
rect 19441 20893 19475 20927
rect 19589 20893 19623 20927
rect 19809 20893 19843 20927
rect 19906 20893 19940 20927
rect 21373 20893 21407 20927
rect 22385 20893 22419 20927
rect 24860 20893 24894 20927
rect 26801 20893 26835 20927
rect 1961 20825 1995 20859
rect 3065 20825 3099 20859
rect 3157 20825 3191 20859
rect 9965 20825 9999 20859
rect 11437 20825 11471 20859
rect 13277 20825 13311 20859
rect 14381 20825 14415 20859
rect 14581 20825 14615 20859
rect 15301 20825 15335 20859
rect 17417 20825 17451 20859
rect 17633 20825 17667 20859
rect 18521 20825 18555 20859
rect 18721 20825 18755 20859
rect 19717 20825 19751 20859
rect 20545 20825 20579 20859
rect 20729 20825 20763 20859
rect 21557 20825 21591 20859
rect 22845 20825 22879 20859
rect 27046 20825 27080 20859
rect 6193 20757 6227 20791
rect 8401 20757 8435 20791
rect 10057 20757 10091 20791
rect 14749 20757 14783 20791
rect 17785 20757 17819 20791
rect 18889 20757 18923 20791
rect 20085 20757 20119 20791
rect 25973 20757 26007 20791
rect 28181 20757 28215 20791
rect 4997 20553 5031 20587
rect 5825 20553 5859 20587
rect 8677 20553 8711 20587
rect 12541 20553 12575 20587
rect 14381 20553 14415 20587
rect 17233 20553 17267 20587
rect 21281 20553 21315 20587
rect 26617 20553 26651 20587
rect 4629 20485 4663 20519
rect 4721 20485 4755 20519
rect 5641 20485 5675 20519
rect 7665 20485 7699 20519
rect 11805 20485 11839 20519
rect 15301 20485 15335 20519
rect 1593 20417 1627 20451
rect 1777 20417 1811 20451
rect 2329 20417 2363 20451
rect 3065 20417 3099 20451
rect 3249 20417 3283 20451
rect 3341 20417 3375 20451
rect 3617 20417 3651 20451
rect 4445 20417 4479 20451
rect 4813 20417 4847 20451
rect 5733 20417 5767 20451
rect 6929 20417 6963 20451
rect 7113 20417 7147 20451
rect 10057 20417 10091 20451
rect 10149 20417 10183 20451
rect 10333 20417 10367 20451
rect 13185 20417 13219 20451
rect 14197 20417 14231 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 16865 20417 16899 20451
rect 17049 20417 17083 20451
rect 17877 20417 17911 20451
rect 18889 20417 18923 20451
rect 19037 20417 19071 20451
rect 19165 20417 19199 20451
rect 19257 20417 19291 20451
rect 19354 20417 19388 20451
rect 20453 20417 20487 20451
rect 20637 20417 20671 20451
rect 20821 20417 20855 20451
rect 21465 20417 21499 20451
rect 22457 20417 22491 20451
rect 24225 20417 24259 20451
rect 25237 20417 25271 20451
rect 25504 20417 25538 20451
rect 3433 20349 3467 20383
rect 5457 20349 5491 20383
rect 8769 20349 8803 20383
rect 8861 20349 8895 20383
rect 12265 20349 12299 20383
rect 12357 20349 12391 20383
rect 13093 20349 13127 20383
rect 14013 20349 14047 20383
rect 17693 20349 17727 20383
rect 18061 20349 18095 20383
rect 22201 20349 22235 20383
rect 1593 20281 1627 20315
rect 7021 20281 7055 20315
rect 11805 20281 11839 20315
rect 2513 20213 2547 20247
rect 3801 20213 3835 20247
rect 6009 20213 6043 20247
rect 7757 20213 7791 20247
rect 8309 20213 8343 20247
rect 10149 20213 10183 20247
rect 13461 20213 13495 20247
rect 15577 20213 15611 20247
rect 15761 20213 15795 20247
rect 19533 20213 19567 20247
rect 23581 20213 23615 20247
rect 24041 20213 24075 20247
rect 2421 20009 2455 20043
rect 4353 20009 4387 20043
rect 4997 20009 5031 20043
rect 8309 20009 8343 20043
rect 9505 20009 9539 20043
rect 12081 20009 12115 20043
rect 12265 20009 12299 20043
rect 13001 20009 13035 20043
rect 13645 20009 13679 20043
rect 14933 20009 14967 20043
rect 15577 20009 15611 20043
rect 16037 20009 16071 20043
rect 17325 20009 17359 20043
rect 18337 20009 18371 20043
rect 19901 20009 19935 20043
rect 21189 20009 21223 20043
rect 22937 20009 22971 20043
rect 5089 19941 5123 19975
rect 8217 19941 8251 19975
rect 17417 19941 17451 19975
rect 19717 19941 19751 19975
rect 22293 19941 22327 19975
rect 5181 19873 5215 19907
rect 6745 19873 6779 19907
rect 9965 19873 9999 19907
rect 15761 19873 15795 19907
rect 26985 19873 27019 19907
rect 1961 19805 1995 19839
rect 2597 19815 2631 19849
rect 2697 19805 2731 19839
rect 2881 19805 2915 19839
rect 2973 19805 3007 19839
rect 4077 19805 4111 19839
rect 4905 19805 4939 19839
rect 5825 19805 5859 19839
rect 6009 19805 6043 19839
rect 6101 19805 6135 19839
rect 6929 19805 6963 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 9137 19805 9171 19839
rect 12817 19805 12851 19839
rect 13553 19805 13587 19839
rect 15577 19805 15611 19839
rect 15853 19805 15887 19839
rect 17233 19805 17267 19839
rect 17509 19805 17543 19839
rect 17693 19805 17727 19839
rect 18153 19805 18187 19839
rect 19441 19805 19475 19839
rect 21833 19805 21867 19839
rect 22477 19805 22511 19839
rect 23121 19805 23155 19839
rect 24041 19805 24075 19839
rect 7849 19737 7883 19771
rect 9321 19737 9355 19771
rect 10232 19737 10266 19771
rect 11897 19737 11931 19771
rect 14749 19737 14783 19771
rect 16957 19737 16991 19771
rect 20821 19737 20855 19771
rect 21005 19737 21039 19771
rect 27230 19737 27264 19771
rect 1777 19669 1811 19703
rect 5641 19669 5675 19703
rect 11345 19669 11379 19703
rect 12097 19669 12131 19703
rect 14949 19669 14983 19703
rect 15117 19669 15151 19703
rect 21649 19669 21683 19703
rect 23857 19669 23891 19703
rect 28365 19669 28399 19703
rect 2789 19465 2823 19499
rect 2973 19465 3007 19499
rect 4175 19465 4209 19499
rect 4261 19465 4295 19499
rect 9051 19465 9085 19499
rect 9965 19465 9999 19499
rect 12541 19465 12575 19499
rect 15117 19465 15151 19499
rect 16221 19465 16255 19499
rect 17601 19465 17635 19499
rect 19257 19465 19291 19499
rect 20361 19465 20395 19499
rect 22477 19465 22511 19499
rect 23397 19465 23431 19499
rect 5733 19397 5767 19431
rect 9873 19397 9907 19431
rect 13093 19397 13127 19431
rect 13293 19397 13327 19431
rect 13921 19397 13955 19431
rect 14126 19397 14160 19431
rect 14749 19397 14783 19431
rect 14965 19397 14999 19431
rect 17233 19397 17267 19431
rect 17449 19397 17483 19431
rect 18889 19397 18923 19431
rect 19089 19397 19123 19431
rect 19901 19397 19935 19431
rect 22017 19397 22051 19431
rect 22937 19397 22971 19431
rect 1961 19329 1995 19363
rect 2053 19329 2087 19363
rect 2237 19329 2271 19363
rect 2329 19329 2363 19363
rect 2914 19329 2948 19363
rect 4077 19329 4111 19363
rect 4353 19329 4387 19363
rect 4997 19329 5031 19363
rect 5181 19329 5215 19363
rect 5273 19329 5307 19363
rect 5917 19329 5951 19363
rect 6009 19329 6043 19363
rect 7021 19329 7055 19363
rect 7849 19329 7883 19363
rect 8953 19329 8987 19363
rect 9137 19329 9171 19363
rect 9229 19329 9263 19363
rect 10517 19329 10551 19363
rect 10701 19329 10735 19363
rect 10977 19329 11011 19363
rect 12265 19329 12299 19363
rect 16313 19329 16347 19363
rect 18061 19329 18095 19363
rect 18243 19329 18277 19363
rect 20821 19329 20855 19363
rect 21005 19329 21039 19363
rect 24297 19329 24331 19363
rect 1777 19261 1811 19295
rect 3433 19261 3467 19295
rect 8125 19261 8159 19295
rect 10793 19261 10827 19295
rect 11897 19261 11931 19295
rect 12173 19261 12207 19295
rect 12382 19261 12416 19295
rect 15945 19261 15979 19295
rect 18429 19261 18463 19295
rect 21189 19261 21223 19295
rect 24041 19261 24075 19295
rect 3341 19193 3375 19227
rect 4997 19193 5031 19227
rect 7205 19193 7239 19227
rect 14289 19193 14323 19227
rect 16037 19193 16071 19227
rect 20177 19193 20211 19227
rect 22293 19193 22327 19227
rect 23305 19193 23339 19227
rect 5733 19125 5767 19159
rect 13277 19125 13311 19159
rect 13461 19125 13495 19159
rect 14105 19125 14139 19159
rect 14933 19125 14967 19159
rect 15577 19125 15611 19159
rect 15853 19125 15887 19159
rect 17417 19125 17451 19159
rect 19073 19125 19107 19159
rect 25421 19125 25455 19159
rect 2881 18921 2915 18955
rect 5365 18921 5399 18955
rect 7757 18921 7791 18955
rect 9689 18921 9723 18955
rect 13093 18921 13127 18955
rect 14657 18921 14691 18955
rect 21649 18921 21683 18955
rect 26801 18921 26835 18955
rect 1593 18853 1627 18887
rect 4353 18853 4387 18887
rect 11345 18853 11379 18887
rect 12081 18853 12115 18887
rect 16589 18853 16623 18887
rect 4629 18785 4663 18819
rect 4813 18785 4847 18819
rect 10701 18785 10735 18819
rect 11186 18785 11220 18819
rect 11805 18785 11839 18819
rect 18889 18785 18923 18819
rect 25421 18785 25455 18819
rect 1777 18717 1811 18751
rect 1869 18717 1903 18751
rect 2053 18717 2087 18751
rect 2145 18717 2179 18751
rect 3065 18717 3099 18751
rect 3157 18717 3191 18751
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 5549 18717 5583 18751
rect 5825 18717 5859 18751
rect 6837 18717 6871 18751
rect 7941 18717 7975 18751
rect 8217 18717 8251 18751
rect 14565 18717 14599 18751
rect 14657 18717 14691 18751
rect 15301 18717 15335 18751
rect 16405 18717 16439 18751
rect 17141 18717 17175 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 19717 18717 19751 18751
rect 19809 18717 19843 18751
rect 19901 18717 19935 18751
rect 20177 18717 20211 18751
rect 22293 18717 22327 18751
rect 24777 18717 24811 18751
rect 7113 18649 7147 18683
rect 9321 18649 9355 18683
rect 9505 18649 9539 18683
rect 12909 18649 12943 18683
rect 14381 18649 14415 18683
rect 17417 18649 17451 18683
rect 21465 18649 21499 18683
rect 21681 18649 21715 18683
rect 22538 18649 22572 18683
rect 25666 18649 25700 18683
rect 5733 18581 5767 18615
rect 8125 18581 8159 18615
rect 10977 18581 11011 18615
rect 11069 18581 11103 18615
rect 12265 18581 12299 18615
rect 13109 18581 13143 18615
rect 13277 18581 13311 18615
rect 14841 18581 14875 18615
rect 15485 18581 15519 18615
rect 17693 18581 17727 18615
rect 19441 18581 19475 18615
rect 20085 18581 20119 18615
rect 21833 18581 21867 18615
rect 23673 18581 23707 18615
rect 24593 18581 24627 18615
rect 2145 18377 2179 18411
rect 10517 18377 10551 18411
rect 18245 18377 18279 18411
rect 20085 18377 20119 18411
rect 23949 18377 23983 18411
rect 26249 18377 26283 18411
rect 3065 18309 3099 18343
rect 4629 18309 4663 18343
rect 4721 18309 4755 18343
rect 5825 18309 5859 18343
rect 12265 18309 12299 18343
rect 12357 18309 12391 18343
rect 12449 18309 12483 18343
rect 14657 18309 14691 18343
rect 20821 18309 20855 18343
rect 2053 18241 2087 18275
rect 2697 18241 2731 18275
rect 2845 18241 2879 18275
rect 2973 18241 3007 18275
rect 3203 18241 3237 18275
rect 4353 18241 4387 18275
rect 4501 18241 4535 18275
rect 4857 18241 4891 18275
rect 5641 18241 5675 18275
rect 5917 18241 5951 18275
rect 6929 18241 6963 18275
rect 8125 18241 8159 18275
rect 8493 18241 8527 18275
rect 8861 18241 8895 18275
rect 9597 18241 9631 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 11161 18241 11195 18275
rect 13645 18241 13679 18275
rect 14013 18241 14047 18275
rect 14841 18241 14875 18275
rect 14933 18241 14967 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 17121 18241 17155 18275
rect 18961 18241 18995 18275
rect 22201 18241 22235 18275
rect 22845 18241 22879 18275
rect 23489 18241 23523 18275
rect 24676 18241 24710 18275
rect 26433 18241 26467 18275
rect 7113 18173 7147 18207
rect 11713 18173 11747 18207
rect 11897 18173 11931 18207
rect 16865 18173 16899 18207
rect 18705 18173 18739 18207
rect 21281 18173 21315 18207
rect 24409 18173 24443 18207
rect 5457 18105 5491 18139
rect 9229 18105 9263 18139
rect 10977 18105 11011 18139
rect 15117 18105 15151 18139
rect 21097 18105 21131 18139
rect 22017 18105 22051 18139
rect 23857 18105 23891 18139
rect 3341 18037 3375 18071
rect 4997 18037 5031 18071
rect 14933 18037 14967 18071
rect 15945 18037 15979 18071
rect 22661 18037 22695 18071
rect 25789 18037 25823 18071
rect 3341 17833 3375 17867
rect 5641 17833 5675 17867
rect 6469 17833 6503 17867
rect 12173 17833 12207 17867
rect 12817 17833 12851 17867
rect 14473 17833 14507 17867
rect 16405 17833 16439 17867
rect 17233 17833 17267 17867
rect 18061 17833 18095 17867
rect 19809 17833 19843 17867
rect 20453 17833 20487 17867
rect 21649 17833 21683 17867
rect 2697 17765 2731 17799
rect 10241 17765 10275 17799
rect 14657 17765 14691 17799
rect 15669 17765 15703 17799
rect 27813 17765 27847 17799
rect 3433 17697 3467 17731
rect 4261 17697 4295 17731
rect 9965 17697 9999 17731
rect 11529 17697 11563 17731
rect 11989 17697 12023 17731
rect 13369 17697 13403 17731
rect 18153 17697 18187 17731
rect 18245 17697 18279 17731
rect 26433 17697 26467 17731
rect 2145 17629 2179 17663
rect 2513 17629 2547 17663
rect 3157 17629 3191 17663
rect 3249 17629 3283 17663
rect 3985 17629 4019 17663
rect 5457 17629 5491 17663
rect 6469 17629 6503 17663
rect 6745 17629 6779 17663
rect 7849 17629 7883 17663
rect 9229 17629 9263 17663
rect 9505 17629 9539 17663
rect 9873 17629 9907 17663
rect 10793 17629 10827 17663
rect 10885 17629 10919 17663
rect 11805 17629 11839 17663
rect 12725 17629 12759 17663
rect 13553 17629 13587 17663
rect 18337 17629 18371 17663
rect 18521 17629 18555 17663
rect 19441 17629 19475 17663
rect 21833 17629 21867 17663
rect 24593 17629 24627 17663
rect 26689 17629 26723 17663
rect 14519 17595 14553 17629
rect 2329 17561 2363 17595
rect 2421 17561 2455 17595
rect 7389 17561 7423 17595
rect 7481 17561 7515 17595
rect 7941 17561 7975 17595
rect 8033 17561 8067 17595
rect 11897 17561 11931 17595
rect 14289 17561 14323 17595
rect 15301 17561 15335 17595
rect 16221 17561 16255 17595
rect 17141 17561 17175 17595
rect 19625 17561 19659 17595
rect 20269 17561 20303 17595
rect 22753 17561 22787 17595
rect 23489 17561 23523 17595
rect 24838 17561 24872 17595
rect 6653 17493 6687 17527
rect 11069 17493 11103 17527
rect 13737 17493 13771 17527
rect 15761 17493 15795 17527
rect 16421 17493 16455 17527
rect 16589 17493 16623 17527
rect 17785 17493 17819 17527
rect 20469 17493 20503 17527
rect 20637 17493 20671 17527
rect 22845 17493 22879 17527
rect 23581 17493 23615 17527
rect 25973 17493 26007 17527
rect 2605 17289 2639 17323
rect 4445 17289 4479 17323
rect 5917 17289 5951 17323
rect 6653 17289 6687 17323
rect 7849 17289 7883 17323
rect 10885 17289 10919 17323
rect 12817 17289 12851 17323
rect 14933 17289 14967 17323
rect 19165 17289 19199 17323
rect 20453 17289 20487 17323
rect 21373 17289 21407 17323
rect 26617 17289 26651 17323
rect 1685 17221 1719 17255
rect 7665 17221 7699 17255
rect 8033 17221 8067 17255
rect 12449 17221 12483 17255
rect 12665 17221 12699 17255
rect 13277 17221 13311 17255
rect 13493 17221 13527 17255
rect 17141 17221 17175 17255
rect 18797 17221 18831 17255
rect 20085 17221 20119 17255
rect 20177 17221 20211 17255
rect 17371 17187 17405 17221
rect 1593 17153 1627 17187
rect 1777 17153 1811 17187
rect 2237 17153 2271 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 3801 17153 3835 17187
rect 3949 17153 3983 17187
rect 4077 17153 4111 17187
rect 4169 17153 4203 17187
rect 4307 17153 4341 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 5273 17153 5307 17187
rect 5365 17153 5399 17187
rect 5825 17153 5859 17187
rect 6561 17153 6595 17187
rect 7757 17153 7791 17187
rect 8585 17153 8619 17187
rect 8769 17153 8803 17187
rect 9597 17153 9631 17187
rect 9965 17153 9999 17187
rect 10333 17153 10367 17187
rect 11069 17153 11103 17187
rect 11713 17153 11747 17187
rect 14105 17153 14139 17187
rect 14289 17153 14323 17187
rect 14473 17153 14507 17187
rect 15117 17153 15151 17187
rect 16221 17153 16255 17187
rect 18521 17153 18555 17187
rect 18669 17153 18703 17187
rect 18889 17153 18923 17187
rect 18986 17153 19020 17187
rect 19809 17153 19843 17187
rect 19957 17153 19991 17187
rect 20315 17153 20349 17187
rect 22017 17153 22051 17187
rect 23469 17153 23503 17187
rect 25493 17153 25527 17187
rect 27353 17153 27387 17187
rect 2789 17085 2823 17119
rect 2881 17085 2915 17119
rect 6929 17085 6963 17119
rect 7021 17085 7055 17119
rect 20913 17085 20947 17119
rect 23213 17085 23247 17119
rect 25237 17085 25271 17119
rect 27905 17085 27939 17119
rect 5181 17017 5215 17051
rect 6837 17017 6871 17051
rect 7481 17017 7515 17051
rect 8953 17017 8987 17051
rect 21189 17017 21223 17051
rect 22385 17017 22419 17051
rect 22477 17017 22511 17051
rect 24593 17017 24627 17051
rect 28181 17017 28215 17051
rect 11897 16949 11931 16983
rect 12633 16949 12667 16983
rect 13461 16949 13495 16983
rect 13645 16949 13679 16983
rect 16037 16949 16071 16983
rect 17325 16949 17359 16983
rect 17509 16949 17543 16983
rect 27169 16949 27203 16983
rect 28365 16949 28399 16983
rect 1777 16745 1811 16779
rect 5181 16745 5215 16779
rect 5641 16745 5675 16779
rect 7573 16745 7607 16779
rect 13553 16745 13587 16779
rect 20821 16745 20855 16779
rect 5089 16677 5123 16711
rect 19809 16677 19843 16711
rect 22293 16677 22327 16711
rect 23581 16677 23615 16711
rect 26157 16677 26191 16711
rect 6653 16609 6687 16643
rect 9321 16609 9355 16643
rect 10793 16609 10827 16643
rect 10977 16609 11011 16643
rect 17141 16609 17175 16643
rect 17509 16609 17543 16643
rect 17969 16609 18003 16643
rect 18337 16609 18371 16643
rect 19441 16609 19475 16643
rect 21465 16609 21499 16643
rect 24777 16609 24811 16643
rect 26617 16609 26651 16643
rect 1961 16541 1995 16575
rect 2237 16541 2271 16575
rect 3065 16541 3099 16575
rect 3433 16541 3467 16575
rect 4077 16541 4111 16575
rect 4261 16541 4295 16575
rect 5825 16541 5859 16575
rect 6101 16541 6135 16575
rect 6837 16541 6871 16575
rect 7113 16541 7147 16575
rect 7849 16541 7883 16575
rect 8309 16541 8343 16575
rect 9137 16541 9171 16575
rect 9689 16541 9723 16575
rect 11345 16541 11379 16575
rect 12081 16541 12115 16575
rect 12633 16541 12667 16575
rect 12725 16541 12759 16575
rect 14289 16541 14323 16575
rect 16129 16541 16163 16575
rect 16405 16541 16439 16575
rect 16497 16541 16531 16575
rect 17325 16541 17359 16575
rect 18153 16541 18187 16575
rect 19625 16541 19659 16575
rect 21005 16541 21039 16575
rect 21097 16541 21131 16575
rect 2145 16473 2179 16507
rect 4721 16473 4755 16507
rect 6009 16473 6043 16507
rect 7573 16473 7607 16507
rect 7757 16473 7791 16507
rect 9873 16473 9907 16507
rect 11437 16473 11471 16507
rect 11529 16473 11563 16507
rect 12265 16473 12299 16507
rect 12817 16473 12851 16507
rect 13369 16473 13403 16507
rect 14534 16473 14568 16507
rect 16313 16473 16347 16507
rect 21189 16473 21223 16507
rect 21307 16473 21341 16507
rect 21925 16473 21959 16507
rect 23213 16473 23247 16507
rect 25022 16473 25056 16507
rect 26862 16473 26896 16507
rect 4261 16405 4295 16439
rect 7021 16405 7055 16439
rect 8493 16405 8527 16439
rect 9781 16405 9815 16439
rect 13569 16405 13603 16439
rect 13737 16405 13771 16439
rect 15669 16405 15703 16439
rect 16681 16405 16715 16439
rect 22385 16405 22419 16439
rect 23673 16405 23707 16439
rect 27997 16405 28031 16439
rect 1869 16201 1903 16235
rect 3893 16201 3927 16235
rect 6009 16201 6043 16235
rect 8861 16201 8895 16235
rect 8953 16201 8987 16235
rect 10425 16201 10459 16235
rect 10977 16201 11011 16235
rect 15577 16201 15611 16235
rect 18061 16201 18095 16235
rect 19349 16201 19383 16235
rect 20545 16201 20579 16235
rect 21189 16201 21223 16235
rect 23765 16201 23799 16235
rect 27353 16201 27387 16235
rect 27997 16201 28031 16235
rect 4997 16133 5031 16167
rect 6561 16133 6595 16167
rect 6761 16133 6795 16167
rect 13553 16133 13587 16167
rect 17417 16133 17451 16167
rect 19947 16133 19981 16167
rect 23305 16133 23339 16167
rect 24492 16133 24526 16167
rect 13783 16099 13817 16133
rect 1685 16065 1719 16099
rect 1961 16065 1995 16099
rect 2605 16065 2639 16099
rect 4813 16065 4847 16099
rect 5089 16065 5123 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 7389 16065 7423 16099
rect 8309 16065 8343 16099
rect 8493 16065 8527 16099
rect 9045 16065 9079 16099
rect 9965 16065 9999 16099
rect 10241 16065 10275 16099
rect 11161 16065 11195 16099
rect 11713 16065 11747 16099
rect 12633 16065 12667 16099
rect 12725 16065 12759 16099
rect 12909 16065 12943 16099
rect 13001 16065 13035 16099
rect 15577 16065 15611 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 16221 16065 16255 16099
rect 17785 16065 17819 16099
rect 18153 16065 18187 16099
rect 18705 16065 18739 16099
rect 18889 16065 18923 16099
rect 20085 16065 20119 16099
rect 21281 16065 21315 16099
rect 27537 16065 27571 16099
rect 28181 16065 28215 16099
rect 7573 15997 7607 16031
rect 10149 15997 10183 16031
rect 19809 15997 19843 16031
rect 20821 15997 20855 16031
rect 22017 15997 22051 16031
rect 24225 15997 24259 16031
rect 19717 15929 19751 15963
rect 22385 15929 22419 15963
rect 23673 15929 23707 15963
rect 1685 15861 1719 15895
rect 4813 15861 4847 15895
rect 6745 15861 6779 15895
rect 6929 15861 6963 15895
rect 10241 15861 10275 15895
rect 11897 15861 11931 15895
rect 12449 15861 12483 15895
rect 13737 15861 13771 15895
rect 13921 15861 13955 15895
rect 17693 15861 17727 15895
rect 17877 15861 17911 15895
rect 19625 15861 19659 15895
rect 20913 15861 20947 15895
rect 21005 15861 21039 15895
rect 22477 15861 22511 15895
rect 25605 15861 25639 15895
rect 2513 15657 2547 15691
rect 5089 15657 5123 15691
rect 17049 15657 17083 15691
rect 18613 15657 18647 15691
rect 20453 15657 20487 15691
rect 21649 15657 21683 15691
rect 23213 15657 23247 15691
rect 28181 15657 28215 15691
rect 4353 15589 4387 15623
rect 5641 15589 5675 15623
rect 8125 15589 8159 15623
rect 14565 15589 14599 15623
rect 14657 15589 14691 15623
rect 18797 15589 18831 15623
rect 20637 15589 20671 15623
rect 21833 15589 21867 15623
rect 23121 15589 23155 15623
rect 25973 15589 26007 15623
rect 4261 15521 4295 15555
rect 6837 15521 6871 15555
rect 9965 15521 9999 15555
rect 11897 15521 11931 15555
rect 14289 15521 14323 15555
rect 14749 15521 14783 15555
rect 17877 15521 17911 15555
rect 1685 15453 1719 15487
rect 1869 15453 1903 15487
rect 2697 15453 2731 15487
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 5003 15453 5037 15487
rect 5181 15453 5215 15487
rect 5825 15453 5859 15487
rect 5917 15453 5951 15487
rect 6101 15453 6135 15487
rect 6193 15453 6227 15487
rect 7113 15453 7147 15487
rect 8401 15453 8435 15487
rect 9781 15453 9815 15487
rect 11161 15453 11195 15487
rect 11253 15453 11287 15487
rect 11437 15453 11471 15487
rect 15025 15453 15059 15487
rect 15669 15453 15703 15487
rect 16681 15453 16715 15487
rect 16865 15453 16899 15487
rect 17509 15453 17543 15487
rect 17693 15453 17727 15487
rect 19441 15453 19475 15487
rect 24593 15453 24627 15487
rect 26801 15453 26835 15487
rect 27068 15453 27102 15487
rect 18659 15419 18693 15453
rect 20499 15419 20533 15453
rect 2973 15385 3007 15419
rect 8125 15385 8159 15419
rect 12153 15385 12187 15419
rect 18429 15385 18463 15419
rect 19625 15385 19659 15419
rect 20269 15385 20303 15419
rect 21465 15385 21499 15419
rect 22753 15385 22787 15419
rect 23765 15385 23799 15419
rect 24860 15385 24894 15419
rect 2881 15317 2915 15351
rect 3985 15317 4019 15351
rect 8309 15317 8343 15351
rect 9413 15317 9447 15351
rect 9873 15317 9907 15351
rect 13277 15317 13311 15351
rect 14933 15317 14967 15351
rect 15485 15317 15519 15351
rect 19809 15317 19843 15351
rect 21665 15317 21699 15351
rect 23857 15317 23891 15351
rect 1777 15113 1811 15147
rect 7389 15113 7423 15147
rect 7573 15113 7607 15147
rect 8217 15113 8251 15147
rect 8953 15113 8987 15147
rect 9321 15113 9355 15147
rect 10701 15113 10735 15147
rect 12541 15113 12575 15147
rect 16037 15113 16071 15147
rect 17509 15113 17543 15147
rect 18061 15113 18095 15147
rect 22017 15113 22051 15147
rect 23121 15113 23155 15147
rect 28089 15113 28123 15147
rect 11713 15045 11747 15079
rect 11929 15045 11963 15079
rect 21005 15045 21039 15079
rect 22293 15045 22327 15079
rect 1961 14977 1995 15011
rect 2053 14977 2087 15011
rect 2237 14977 2271 15011
rect 2329 14977 2363 15011
rect 2881 14977 2915 15011
rect 5549 14977 5583 15011
rect 8309 14977 8343 15011
rect 8493 14977 8527 15011
rect 10149 14977 10183 15011
rect 10425 14977 10459 15011
rect 10701 14977 10735 15011
rect 12725 14977 12759 15011
rect 13461 14977 13495 15011
rect 13737 14977 13771 15011
rect 14013 14977 14047 15011
rect 14197 14977 14231 15011
rect 15117 14977 15151 15011
rect 15393 14977 15427 15011
rect 16221 14977 16255 15011
rect 17141 14977 17175 15011
rect 17233 14977 17267 15011
rect 17601 14977 17635 15011
rect 18245 14977 18279 15011
rect 18961 14977 18995 15011
rect 20637 14977 20671 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 21123 14977 21157 15011
rect 22202 14977 22236 15011
rect 22385 14977 22419 15011
rect 22503 14977 22537 15011
rect 23305 14977 23339 15011
rect 24205 14977 24239 15011
rect 9413 14909 9447 14943
rect 9505 14909 9539 14943
rect 15301 14909 15335 14943
rect 16865 14909 16899 14943
rect 18705 14909 18739 14943
rect 21281 14909 21315 14943
rect 22661 14909 22695 14943
rect 23949 14909 23983 14943
rect 27629 14909 27663 14943
rect 7021 14841 7055 14875
rect 11161 14841 11195 14875
rect 12081 14841 12115 14875
rect 13829 14841 13863 14875
rect 13921 14841 13955 14875
rect 17325 14841 17359 14875
rect 27905 14841 27939 14875
rect 4169 14773 4203 14807
rect 5641 14773 5675 14807
rect 7389 14773 7423 14807
rect 8033 14773 8067 14807
rect 11897 14773 11931 14807
rect 15209 14773 15243 14807
rect 15577 14773 15611 14807
rect 20085 14773 20119 14807
rect 25329 14773 25363 14807
rect 1685 14569 1719 14603
rect 3249 14569 3283 14603
rect 3433 14569 3467 14603
rect 4997 14569 5031 14603
rect 8493 14569 8527 14603
rect 9505 14569 9539 14603
rect 11345 14569 11379 14603
rect 13277 14569 13311 14603
rect 14749 14569 14783 14603
rect 15669 14569 15703 14603
rect 16129 14569 16163 14603
rect 17325 14569 17359 14603
rect 17601 14569 17635 14603
rect 18705 14569 18739 14603
rect 20453 14569 20487 14603
rect 20637 14569 20671 14603
rect 21465 14569 21499 14603
rect 27629 14569 27663 14603
rect 12081 14501 12115 14535
rect 14565 14501 14599 14535
rect 15577 14501 15611 14535
rect 18889 14501 18923 14535
rect 22569 14501 22603 14535
rect 23397 14501 23431 14535
rect 5457 14433 5491 14467
rect 9137 14433 9171 14467
rect 14289 14433 14323 14467
rect 16497 14433 16531 14467
rect 22661 14433 22695 14467
rect 1869 14365 1903 14399
rect 2145 14365 2179 14399
rect 4169 14365 4203 14399
rect 4261 14365 4295 14399
rect 4445 14365 4479 14399
rect 4537 14365 4571 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 5365 14365 5399 14399
rect 6377 14365 6411 14399
rect 6653 14365 6687 14399
rect 7573 14365 7607 14399
rect 8309 14365 8343 14399
rect 9321 14365 9355 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 11989 14365 12023 14399
rect 12173 14365 12207 14399
rect 13093 14365 13127 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 16405 14365 16439 14399
rect 16589 14365 16623 14399
rect 16681 14365 16715 14399
rect 16865 14365 16899 14399
rect 17693 14365 17727 14399
rect 17785 14365 17819 14399
rect 17877 14365 17911 14399
rect 18061 14365 18095 14399
rect 24777 14365 24811 14399
rect 25421 14365 25455 14399
rect 26249 14365 26283 14399
rect 3295 14331 3329 14365
rect 20499 14331 20533 14365
rect 21511 14331 21545 14365
rect 3065 14297 3099 14331
rect 11161 14297 11195 14331
rect 11361 14297 11395 14331
rect 15209 14297 15243 14331
rect 18521 14297 18555 14331
rect 18737 14297 18771 14331
rect 20269 14297 20303 14331
rect 21281 14297 21315 14331
rect 22201 14297 22235 14331
rect 23121 14297 23155 14331
rect 26494 14297 26528 14331
rect 2053 14229 2087 14263
rect 3985 14229 4019 14263
rect 6193 14229 6227 14263
rect 6561 14229 6595 14263
rect 7757 14229 7791 14263
rect 10517 14229 10551 14263
rect 11529 14229 11563 14263
rect 12817 14229 12851 14263
rect 21649 14229 21683 14263
rect 23581 14229 23615 14263
rect 24593 14229 24627 14263
rect 25237 14229 25271 14263
rect 1593 14025 1627 14059
rect 5641 14025 5675 14059
rect 6561 14025 6595 14059
rect 9321 14025 9355 14059
rect 13553 14025 13587 14059
rect 14289 14025 14323 14059
rect 15853 14025 15887 14059
rect 18613 14025 18647 14059
rect 20545 14025 20579 14059
rect 21281 14025 21315 14059
rect 24041 14025 24075 14059
rect 26617 14025 26651 14059
rect 28089 14025 28123 14059
rect 9873 13957 9907 13991
rect 10057 13957 10091 13991
rect 15485 13957 15519 13991
rect 15685 13957 15719 13991
rect 17417 13957 17451 13991
rect 17617 13957 17651 13991
rect 18245 13957 18279 13991
rect 19441 13957 19475 13991
rect 20177 13957 20211 13991
rect 20269 13957 20303 13991
rect 22503 13957 22537 13991
rect 25504 13957 25538 13991
rect 18475 13923 18509 13957
rect 1777 13889 1811 13923
rect 1961 13889 1995 13923
rect 2237 13889 2271 13923
rect 3249 13889 3283 13923
rect 3801 13889 3835 13923
rect 4721 13889 4755 13923
rect 4813 13889 4847 13923
rect 4997 13889 5031 13923
rect 5273 13889 5307 13923
rect 5549 13889 5583 13923
rect 6745 13889 6779 13923
rect 6837 13889 6871 13923
rect 7095 13889 7129 13923
rect 7941 13889 7975 13923
rect 8217 13889 8251 13923
rect 8493 13889 8527 13923
rect 8677 13889 8711 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 11969 13889 12003 13923
rect 13737 13889 13771 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14657 13889 14691 13923
rect 14933 13889 14967 13923
rect 19257 13889 19291 13923
rect 19901 13889 19935 13923
rect 19994 13889 20028 13923
rect 20366 13889 20400 13923
rect 21465 13889 21499 13923
rect 22201 13889 22235 13923
rect 22293 13889 22327 13923
rect 22386 13889 22420 13923
rect 22661 13889 22695 13923
rect 24225 13889 24259 13923
rect 28273 13889 28307 13923
rect 2053 13821 2087 13855
rect 3433 13821 3467 13855
rect 3525 13821 3559 13855
rect 8401 13821 8435 13855
rect 10241 13821 10275 13855
rect 11713 13821 11747 13855
rect 19073 13821 19107 13855
rect 22017 13821 22051 13855
rect 23121 13821 23155 13855
rect 25237 13821 25271 13855
rect 27169 13821 27203 13855
rect 1869 13753 1903 13787
rect 3341 13753 3375 13787
rect 7021 13753 7055 13787
rect 11069 13753 11103 13787
rect 23397 13753 23431 13787
rect 27445 13753 27479 13787
rect 3617 13685 3651 13719
rect 13093 13685 13127 13719
rect 15669 13685 15703 13719
rect 17601 13685 17635 13719
rect 17785 13685 17819 13719
rect 18429 13685 18463 13719
rect 23581 13685 23615 13719
rect 27629 13685 27663 13719
rect 5457 13481 5491 13515
rect 9137 13481 9171 13515
rect 10149 13481 10183 13515
rect 13369 13481 13403 13515
rect 14565 13481 14599 13515
rect 21281 13481 21315 13515
rect 24041 13481 24075 13515
rect 25973 13481 26007 13515
rect 3065 13413 3099 13447
rect 5641 13413 5675 13447
rect 8493 13413 8527 13447
rect 9597 13413 9631 13447
rect 11069 13413 11103 13447
rect 17785 13413 17819 13447
rect 21465 13413 21499 13447
rect 22753 13413 22787 13447
rect 23857 13413 23891 13447
rect 10793 13345 10827 13379
rect 13001 13345 13035 13379
rect 14381 13345 14415 13379
rect 1685 13277 1719 13311
rect 1952 13277 1986 13311
rect 4261 13277 4295 13311
rect 5089 13277 5123 13311
rect 6653 13277 6687 13311
rect 7113 13277 7147 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 8033 13277 8067 13311
rect 8217 13277 8251 13311
rect 8585 13277 8619 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 9689 13277 9723 13311
rect 10333 13277 10367 13311
rect 13093 13277 13127 13311
rect 14565 13277 14599 13311
rect 15945 13277 15979 13311
rect 16037 13277 16071 13311
rect 17141 13277 17175 13311
rect 17289 13277 17323 13311
rect 17606 13277 17640 13311
rect 18429 13277 18463 13311
rect 18613 13277 18647 13311
rect 19993 13277 20027 13311
rect 20086 13277 20120 13311
rect 20269 13277 20303 13311
rect 20499 13277 20533 13311
rect 24593 13277 24627 13311
rect 26433 13277 26467 13311
rect 26700 13277 26734 13311
rect 6285 13209 6319 13243
rect 6469 13209 6503 13243
rect 11713 13209 11747 13243
rect 11897 13209 11931 13243
rect 14289 13209 14323 13243
rect 17417 13209 17451 13243
rect 17509 13209 17543 13243
rect 20361 13209 20395 13243
rect 21097 13209 21131 13243
rect 22385 13209 22419 13243
rect 23581 13209 23615 13243
rect 24860 13209 24894 13243
rect 4445 13141 4479 13175
rect 5457 13141 5491 13175
rect 7297 13141 7331 13175
rect 11253 13141 11287 13175
rect 12081 13141 12115 13175
rect 14749 13141 14783 13175
rect 16221 13141 16255 13175
rect 18797 13141 18831 13175
rect 20637 13141 20671 13175
rect 21297 13141 21331 13175
rect 22845 13141 22879 13175
rect 27813 13141 27847 13175
rect 2145 12937 2179 12971
rect 3449 12937 3483 12971
rect 3617 12937 3651 12971
rect 5181 12937 5215 12971
rect 5917 12937 5951 12971
rect 7481 12937 7515 12971
rect 8493 12937 8527 12971
rect 12081 12937 12115 12971
rect 13921 12937 13955 12971
rect 15025 12937 15059 12971
rect 18337 12937 18371 12971
rect 18889 12937 18923 12971
rect 19901 12937 19935 12971
rect 22661 12937 22695 12971
rect 28089 12937 28123 12971
rect 3249 12869 3283 12903
rect 10609 12869 10643 12903
rect 11759 12869 11793 12903
rect 11913 12869 11947 12903
rect 17141 12869 17175 12903
rect 17969 12869 18003 12903
rect 18169 12869 18203 12903
rect 21465 12869 21499 12903
rect 24317 12869 24351 12903
rect 27169 12869 27203 12903
rect 2421 12801 2455 12835
rect 2513 12801 2547 12835
rect 2605 12801 2639 12835
rect 2789 12801 2823 12835
rect 4445 12801 4479 12835
rect 5089 12801 5123 12835
rect 5733 12801 5767 12835
rect 6837 12801 6871 12835
rect 7389 12801 7423 12835
rect 8309 12801 8343 12835
rect 8585 12801 8619 12835
rect 9045 12801 9079 12835
rect 9229 12801 9263 12835
rect 9689 12801 9723 12835
rect 10793 12801 10827 12835
rect 12541 12801 12575 12835
rect 12808 12801 12842 12835
rect 14565 12801 14599 12835
rect 15485 12801 15519 12835
rect 15577 12801 15611 12835
rect 15761 12801 15795 12835
rect 16872 12801 16906 12835
rect 16958 12801 16992 12835
rect 17233 12801 17267 12835
rect 17371 12801 17405 12835
rect 19257 12801 19291 12835
rect 20085 12801 20119 12835
rect 20177 12801 20211 12835
rect 21281 12801 21315 12835
rect 22293 12801 22327 12835
rect 22753 12801 22787 12835
rect 23581 12801 23615 12835
rect 24133 12801 24167 12835
rect 25237 12801 25271 12835
rect 25493 12801 25527 12835
rect 28273 12801 28307 12835
rect 4537 12733 4571 12767
rect 4721 12733 4755 12767
rect 7481 12733 7515 12767
rect 15393 12733 15427 12767
rect 19073 12733 19107 12767
rect 19165 12733 19199 12767
rect 19349 12733 19383 12767
rect 20269 12733 20303 12767
rect 20361 12733 20395 12767
rect 21097 12733 21131 12767
rect 10149 12665 10183 12699
rect 14381 12665 14415 12699
rect 23397 12665 23431 12699
rect 27445 12665 27479 12699
rect 3433 12597 3467 12631
rect 8125 12597 8159 12631
rect 9137 12597 9171 12631
rect 9965 12597 9999 12631
rect 10977 12597 11011 12631
rect 11897 12597 11931 12631
rect 15301 12597 15335 12631
rect 17509 12597 17543 12631
rect 18153 12597 18187 12631
rect 22017 12597 22051 12631
rect 22385 12597 22419 12631
rect 22477 12597 22511 12631
rect 26617 12597 26651 12631
rect 27629 12597 27663 12631
rect 2329 12393 2363 12427
rect 4445 12393 4479 12427
rect 5733 12393 5767 12427
rect 5917 12393 5951 12427
rect 7941 12393 7975 12427
rect 10701 12393 10735 12427
rect 13001 12393 13035 12427
rect 14933 12393 14967 12427
rect 15945 12393 15979 12427
rect 16681 12393 16715 12427
rect 16865 12393 16899 12427
rect 17509 12393 17543 12427
rect 18429 12393 18463 12427
rect 18613 12393 18647 12427
rect 19625 12393 19659 12427
rect 28365 12393 28399 12427
rect 3341 12325 3375 12359
rect 7297 12325 7331 12359
rect 8217 12325 8251 12359
rect 8309 12325 8343 12359
rect 12357 12325 12391 12359
rect 15117 12325 15151 12359
rect 17693 12325 17727 12359
rect 21741 12325 21775 12359
rect 22753 12325 22787 12359
rect 23673 12325 23707 12359
rect 10609 12257 10643 12291
rect 10793 12257 10827 12291
rect 12081 12257 12115 12291
rect 21925 12257 21959 12291
rect 26985 12257 27019 12291
rect 1777 12189 1811 12223
rect 2145 12189 2179 12223
rect 3249 12189 3283 12223
rect 4629 12189 4663 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 6377 12189 6411 12223
rect 6561 12189 6595 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 8125 12189 8159 12223
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 9321 12189 9355 12223
rect 9873 12189 9907 12223
rect 10517 12189 10551 12223
rect 11437 12189 11471 12223
rect 13185 12189 13219 12223
rect 15577 12189 15611 12223
rect 15761 12189 15795 12223
rect 20821 12189 20855 12223
rect 21005 12189 21039 12223
rect 24777 12189 24811 12223
rect 14979 12155 15013 12189
rect 1961 12121 1995 12155
rect 2053 12121 2087 12155
rect 5549 12121 5583 12155
rect 6469 12121 6503 12155
rect 10057 12121 10091 12155
rect 14749 12121 14783 12155
rect 16497 12121 16531 12155
rect 16702 12121 16736 12155
rect 17325 12121 17359 12155
rect 18245 12121 18279 12155
rect 19441 12121 19475 12155
rect 20637 12121 20671 12155
rect 21465 12121 21499 12155
rect 22385 12121 22419 12155
rect 23305 12121 23339 12155
rect 27230 12121 27264 12155
rect 5759 12053 5793 12087
rect 9137 12053 9171 12087
rect 11253 12053 11287 12087
rect 12541 12053 12575 12087
rect 17525 12053 17559 12087
rect 18445 12053 18479 12087
rect 19641 12053 19675 12087
rect 19809 12053 19843 12087
rect 22845 12053 22879 12087
rect 23765 12053 23799 12087
rect 24593 12053 24627 12087
rect 2973 11849 3007 11883
rect 3801 11849 3835 11883
rect 4629 11849 4663 11883
rect 5549 11849 5583 11883
rect 13093 11849 13127 11883
rect 13645 11849 13679 11883
rect 15577 11849 15611 11883
rect 18889 11849 18923 11883
rect 19441 11849 19475 11883
rect 25053 11849 25087 11883
rect 27905 11849 27939 11883
rect 1777 11781 1811 11815
rect 8125 11781 8159 11815
rect 11969 11781 12003 11815
rect 15117 11781 15151 11815
rect 17141 11781 17175 11815
rect 17357 11781 17391 11815
rect 27445 11781 27479 11815
rect 1961 11713 1995 11747
rect 2605 11713 2639 11747
rect 2789 11713 2823 11747
rect 3709 11713 3743 11747
rect 3893 11713 3927 11747
rect 3985 11713 4019 11747
rect 4629 11713 4663 11747
rect 5365 11713 5399 11747
rect 5641 11713 5675 11747
rect 6653 11713 6687 11747
rect 6929 11713 6963 11747
rect 7757 11713 7791 11747
rect 8953 11713 8987 11747
rect 9045 11713 9079 11747
rect 9321 11713 9355 11747
rect 9781 11713 9815 11747
rect 10057 11713 10091 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 11713 11713 11747 11747
rect 13645 11713 13679 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14289 11713 14323 11747
rect 14933 11713 14967 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 18705 11713 18739 11747
rect 19625 11713 19659 11747
rect 20341 11713 20375 11747
rect 22109 11713 22143 11747
rect 23213 11713 23247 11747
rect 23929 11713 23963 11747
rect 26617 11713 26651 11747
rect 6745 11645 6779 11679
rect 7941 11645 7975 11679
rect 10149 11645 10183 11679
rect 18521 11645 18555 11679
rect 20085 11645 20119 11679
rect 23673 11645 23707 11679
rect 5181 11577 5215 11611
rect 7849 11577 7883 11611
rect 15853 11577 15887 11611
rect 17509 11577 17543 11611
rect 21465 11577 21499 11611
rect 27721 11577 27755 11611
rect 2145 11509 2179 11543
rect 6929 11509 6963 11543
rect 7113 11509 7147 11543
rect 8769 11509 8803 11543
rect 9229 11509 9263 11543
rect 16037 11509 16071 11543
rect 17325 11509 17359 11543
rect 22201 11509 22235 11543
rect 23029 11509 23063 11543
rect 26433 11509 26467 11543
rect 3985 11305 4019 11339
rect 5549 11305 5583 11339
rect 5733 11305 5767 11339
rect 10425 11305 10459 11339
rect 10517 11305 10551 11339
rect 11897 11305 11931 11339
rect 13277 11305 13311 11339
rect 13645 11305 13679 11339
rect 15393 11305 15427 11339
rect 15577 11305 15611 11339
rect 16221 11305 16255 11339
rect 16865 11305 16899 11339
rect 17325 11305 17359 11339
rect 20453 11305 20487 11339
rect 24041 11305 24075 11339
rect 26249 11305 26283 11339
rect 3157 11237 3191 11271
rect 5181 11237 5215 11271
rect 6193 11237 6227 11271
rect 6929 11237 6963 11271
rect 7849 11237 7883 11271
rect 9781 11237 9815 11271
rect 12265 11237 12299 11271
rect 14657 11237 14691 11271
rect 16405 11237 16439 11271
rect 18705 11237 18739 11271
rect 20637 11237 20671 11271
rect 22017 11237 22051 11271
rect 2237 11169 2271 11203
rect 8309 11169 8343 11203
rect 8493 11169 8527 11203
rect 10609 11169 10643 11203
rect 12173 11169 12207 11203
rect 13369 11169 13403 11203
rect 14749 11169 14783 11203
rect 17049 11169 17083 11203
rect 18889 11169 18923 11203
rect 22661 11169 22695 11203
rect 1777 11101 1811 11135
rect 1961 11101 1995 11135
rect 2697 11101 2731 11135
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 4169 11101 4203 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 6469 11101 6503 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 10333 11101 10367 11135
rect 11437 11101 11471 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 12633 11101 12667 11135
rect 13461 11101 13495 11135
rect 14289 11101 14323 11135
rect 17141 11101 17175 11135
rect 17969 11101 18003 11135
rect 19441 11101 19475 11135
rect 22201 11101 22235 11135
rect 24869 11101 24903 11135
rect 26893 11101 26927 11135
rect 27149 11101 27183 11135
rect 20499 11067 20533 11101
rect 1869 11033 1903 11067
rect 2099 11033 2133 11067
rect 5549 11033 5583 11067
rect 6193 11033 6227 11067
rect 8217 11033 8251 11067
rect 9413 11033 9447 11067
rect 13185 11033 13219 11067
rect 15235 11033 15269 11067
rect 15425 11033 15459 11067
rect 16037 11033 16071 11067
rect 16865 11033 16899 11067
rect 18429 11033 18463 11067
rect 19625 11033 19659 11067
rect 20269 11033 20303 11067
rect 21097 11033 21131 11067
rect 21281 11033 21315 11067
rect 21465 11033 21499 11067
rect 22928 11033 22962 11067
rect 25136 11033 25170 11067
rect 1593 10965 1627 10999
rect 6377 10965 6411 10999
rect 9873 10965 9907 10999
rect 11253 10965 11287 10999
rect 16247 10965 16281 10999
rect 17785 10965 17819 10999
rect 19809 10965 19843 10999
rect 28273 10965 28307 10999
rect 1977 10761 2011 10795
rect 2145 10761 2179 10795
rect 5289 10761 5323 10795
rect 14289 10761 14323 10795
rect 16313 10761 16347 10795
rect 17065 10761 17099 10795
rect 17233 10761 17267 10795
rect 18353 10761 18387 10795
rect 18521 10761 18555 10795
rect 20177 10761 20211 10795
rect 22477 10761 22511 10795
rect 25053 10761 25087 10795
rect 1777 10693 1811 10727
rect 2605 10693 2639 10727
rect 5089 10693 5123 10727
rect 7573 10693 7607 10727
rect 8401 10693 8435 10727
rect 12418 10693 12452 10727
rect 15945 10693 15979 10727
rect 16145 10693 16179 10727
rect 16865 10693 16899 10727
rect 18153 10693 18187 10727
rect 18981 10693 19015 10727
rect 19809 10693 19843 10727
rect 20009 10693 20043 10727
rect 19211 10659 19245 10693
rect 6745 10625 6779 10659
rect 7021 10625 7055 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 9413 10625 9447 10659
rect 9873 10625 9907 10659
rect 10977 10625 11011 10659
rect 12173 10625 12207 10659
rect 14197 10625 14231 10659
rect 14841 10625 14875 10659
rect 15117 10625 15151 10659
rect 20637 10625 20671 10659
rect 20821 10625 20855 10659
rect 23029 10625 23063 10659
rect 23929 10625 23963 10659
rect 25697 10625 25731 10659
rect 26341 10625 26375 10659
rect 8769 10557 8803 10591
rect 15025 10557 15059 10591
rect 22017 10557 22051 10591
rect 23213 10557 23247 10591
rect 23673 10557 23707 10591
rect 3893 10489 3927 10523
rect 9229 10489 9263 10523
rect 10793 10489 10827 10523
rect 22385 10489 22419 10523
rect 25513 10489 25547 10523
rect 1961 10421 1995 10455
rect 5273 10421 5307 10455
rect 5457 10421 5491 10455
rect 7573 10421 7607 10455
rect 10057 10421 10091 10455
rect 13553 10421 13587 10455
rect 15117 10421 15151 10455
rect 15301 10421 15335 10455
rect 16129 10421 16163 10455
rect 17049 10421 17083 10455
rect 18337 10421 18371 10455
rect 19165 10421 19199 10455
rect 19349 10421 19383 10455
rect 19993 10421 20027 10455
rect 21005 10421 21039 10455
rect 26157 10421 26191 10455
rect 5641 10217 5675 10251
rect 6101 10217 6135 10251
rect 7849 10217 7883 10251
rect 9505 10217 9539 10251
rect 9965 10217 9999 10251
rect 10241 10217 10275 10251
rect 11621 10217 11655 10251
rect 13001 10217 13035 10251
rect 13185 10217 13219 10251
rect 15669 10217 15703 10251
rect 17325 10217 17359 10251
rect 28365 10217 28399 10251
rect 6561 10149 6595 10183
rect 10333 10149 10367 10183
rect 19625 10149 19659 10183
rect 21005 10149 21039 10183
rect 21925 10149 21959 10183
rect 22109 10149 22143 10183
rect 22937 10149 22971 10183
rect 23029 10149 23063 10183
rect 23857 10149 23891 10183
rect 3065 10081 3099 10115
rect 5825 10081 5859 10115
rect 7941 10081 7975 10115
rect 12909 10081 12943 10115
rect 14289 10081 14323 10115
rect 21649 10081 21683 10115
rect 1593 10013 1627 10047
rect 1869 10013 1903 10047
rect 3249 10013 3283 10047
rect 4629 10013 4663 10047
rect 4721 10013 4755 10047
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 5917 10013 5951 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7665 10013 7699 10047
rect 8585 10013 8619 10047
rect 9321 10013 9355 10047
rect 10425 10013 10459 10047
rect 10701 10013 10735 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 13001 10013 13035 10047
rect 14545 10013 14579 10047
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 18153 10013 18187 10047
rect 19441 10013 19475 10047
rect 25145 10013 25179 10047
rect 26985 10013 27019 10047
rect 5641 9945 5675 9979
rect 9137 9945 9171 9979
rect 11897 9945 11931 9979
rect 12127 9945 12161 9979
rect 12725 9945 12759 9979
rect 17233 9945 17267 9979
rect 20637 9945 20671 9979
rect 22569 9945 22603 9979
rect 23489 9945 23523 9979
rect 25390 9945 25424 9979
rect 27230 9945 27264 9979
rect 3433 9877 3467 9911
rect 4445 9877 4479 9911
rect 6745 9877 6779 9911
rect 7481 9877 7515 9911
rect 8401 9877 8435 9911
rect 10609 9877 10643 9911
rect 16497 9877 16531 9911
rect 18245 9877 18279 9911
rect 21097 9877 21131 9911
rect 23949 9877 23983 9911
rect 26525 9877 26559 9911
rect 4077 9673 4111 9707
rect 8309 9673 8343 9707
rect 9229 9673 9263 9707
rect 1838 9605 1872 9639
rect 4721 9605 4755 9639
rect 6653 9605 6687 9639
rect 7021 9605 7055 9639
rect 10333 9605 10367 9639
rect 12081 9605 12115 9639
rect 12199 9605 12233 9639
rect 12909 9605 12943 9639
rect 14381 9605 14415 9639
rect 14581 9605 14615 9639
rect 15117 9605 15151 9639
rect 15333 9605 15367 9639
rect 17693 9605 17727 9639
rect 19257 9605 19291 9639
rect 20269 9605 20303 9639
rect 1593 9537 1627 9571
rect 3893 9537 3927 9571
rect 4169 9537 4203 9571
rect 4629 9537 4663 9571
rect 4813 9537 4847 9571
rect 5273 9537 5307 9571
rect 5457 9537 5491 9571
rect 7941 9537 7975 9571
rect 8125 9537 8159 9571
rect 9873 9537 9907 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12311 9537 12345 9571
rect 13737 9537 13771 9571
rect 13921 9537 13955 9571
rect 16313 9537 16347 9571
rect 16957 9537 16991 9571
rect 18061 9537 18095 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 19073 9537 19107 9571
rect 21281 9537 21315 9571
rect 22201 9537 22235 9571
rect 22845 9537 22879 9571
rect 23581 9537 23615 9571
rect 24501 9537 24535 9571
rect 24768 9537 24802 9571
rect 26525 9537 26559 9571
rect 8769 9469 8803 9503
rect 10793 9469 10827 9503
rect 9137 9401 9171 9435
rect 10701 9401 10735 9435
rect 11713 9401 11747 9435
rect 14749 9401 14783 9435
rect 15485 9401 15519 9435
rect 18153 9401 18187 9435
rect 20545 9401 20579 9435
rect 22017 9401 22051 9435
rect 23397 9401 23431 9435
rect 26341 9401 26375 9435
rect 2973 9333 3007 9367
rect 3709 9333 3743 9367
rect 5641 9333 5675 9367
rect 9689 9333 9723 9367
rect 13001 9333 13035 9367
rect 13829 9333 13863 9367
rect 14565 9333 14599 9367
rect 15301 9333 15335 9367
rect 15761 9333 15795 9367
rect 16129 9333 16163 9367
rect 17049 9333 17083 9367
rect 17969 9333 18003 9367
rect 19441 9333 19475 9367
rect 20729 9333 20763 9367
rect 21373 9333 21407 9367
rect 22661 9333 22695 9367
rect 25881 9333 25915 9367
rect 1685 9129 1719 9163
rect 2513 9129 2547 9163
rect 3249 9129 3283 9163
rect 4905 9129 4939 9163
rect 6745 9129 6779 9163
rect 8401 9129 8435 9163
rect 9781 9129 9815 9163
rect 11529 9129 11563 9163
rect 11713 9129 11747 9163
rect 12357 9129 12391 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 13461 9129 13495 9163
rect 14565 9129 14599 9163
rect 15485 9129 15519 9163
rect 15669 9129 15703 9163
rect 18153 9129 18187 9163
rect 19625 9129 19659 9163
rect 20637 9129 20671 9163
rect 24041 9129 24075 9163
rect 25973 9129 26007 9163
rect 28089 9129 28123 9163
rect 4353 9061 4387 9095
rect 7481 9061 7515 9095
rect 8309 9061 8343 9095
rect 9965 9061 9999 9095
rect 10701 9061 10735 9095
rect 13277 9061 13311 9095
rect 19809 9061 19843 9095
rect 21097 9061 21131 9095
rect 3985 8993 4019 9027
rect 8493 8993 8527 9027
rect 13369 8993 13403 9027
rect 14381 8993 14415 9027
rect 26709 8993 26743 9027
rect 1685 8925 1719 8959
rect 1869 8925 1903 8959
rect 2421 8925 2455 8959
rect 2605 8925 2639 8959
rect 4169 8925 4203 8959
rect 4813 8925 4847 8959
rect 5457 8925 5491 8959
rect 5641 8925 5675 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 7757 8925 7791 8959
rect 8217 8925 8251 8959
rect 10425 8925 10459 8959
rect 13553 8925 13587 8959
rect 13737 8925 13771 8959
rect 14565 8925 14599 8959
rect 16129 8925 16163 8959
rect 16385 8925 16419 8959
rect 21281 8925 21315 8959
rect 21925 8925 21959 8959
rect 22661 8925 22695 8959
rect 24593 8925 24627 8959
rect 26965 8925 26999 8959
rect 3065 8857 3099 8891
rect 6469 8857 6503 8891
rect 9597 8857 9631 8891
rect 11345 8857 11379 8891
rect 11561 8857 11595 8891
rect 12173 8857 12207 8891
rect 12373 8857 12407 8891
rect 14289 8857 14323 8891
rect 15301 8857 15335 8891
rect 17969 8857 18003 8891
rect 18185 8857 18219 8891
rect 19441 8857 19475 8891
rect 20269 8857 20303 8891
rect 20453 8857 20487 8891
rect 22906 8857 22940 8891
rect 24838 8857 24872 8891
rect 3265 8789 3299 8823
rect 3433 8789 3467 8823
rect 5825 8789 5859 8823
rect 6929 8789 6963 8823
rect 7481 8789 7515 8823
rect 7573 8789 7607 8823
rect 9807 8789 9841 8823
rect 10885 8789 10919 8823
rect 14749 8789 14783 8823
rect 15511 8789 15545 8823
rect 17509 8789 17543 8823
rect 18337 8789 18371 8823
rect 19641 8789 19675 8823
rect 21741 8789 21775 8823
rect 3617 8585 3651 8619
rect 4537 8585 4571 8619
rect 9137 8585 9171 8619
rect 11161 8585 11195 8619
rect 13093 8585 13127 8619
rect 14933 8585 14967 8619
rect 15593 8585 15627 8619
rect 15761 8585 15795 8619
rect 17065 8585 17099 8619
rect 17233 8585 17267 8619
rect 17903 8585 17937 8619
rect 22017 8585 22051 8619
rect 24501 8585 24535 8619
rect 1838 8517 1872 8551
rect 5549 8517 5583 8551
rect 7205 8517 7239 8551
rect 7665 8517 7699 8551
rect 8677 8517 8711 8551
rect 11958 8517 11992 8551
rect 14565 8517 14599 8551
rect 15393 8517 15427 8551
rect 16865 8517 16899 8551
rect 17693 8517 17727 8551
rect 18705 8517 18739 8551
rect 18889 8517 18923 8551
rect 23366 8517 23400 8551
rect 25228 8517 25262 8551
rect 1593 8449 1627 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 4169 8449 4203 8483
rect 4537 8449 4571 8483
rect 5365 8449 5399 8483
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 10048 8449 10082 8483
rect 13553 8449 13587 8483
rect 14289 8449 14323 8483
rect 14437 8449 14471 8483
rect 14657 8449 14691 8483
rect 14795 8449 14829 8483
rect 18521 8449 18555 8483
rect 19349 8449 19383 8483
rect 19533 8449 19567 8483
rect 20361 8449 20395 8483
rect 21005 8449 21039 8483
rect 22201 8449 22235 8483
rect 4445 8381 4479 8415
rect 5733 8381 5767 8415
rect 8125 8381 8159 8415
rect 9781 8381 9815 8415
rect 11713 8381 11747 8415
rect 19717 8381 19751 8415
rect 23121 8381 23155 8415
rect 24961 8381 24995 8415
rect 2973 8313 3007 8347
rect 8033 8313 8067 8347
rect 9045 8313 9079 8347
rect 20177 8313 20211 8347
rect 20821 8313 20855 8347
rect 26341 8313 26375 8347
rect 4261 8245 4295 8279
rect 13737 8245 13771 8279
rect 15577 8245 15611 8279
rect 17049 8245 17083 8279
rect 17877 8245 17911 8279
rect 18061 8245 18095 8279
rect 3065 8041 3099 8075
rect 4445 8041 4479 8075
rect 6929 8041 6963 8075
rect 10425 8041 10459 8075
rect 11897 8041 11931 8075
rect 12081 8041 12115 8075
rect 15669 8041 15703 8075
rect 15945 8041 15979 8075
rect 19625 8041 19659 8075
rect 23305 8041 23339 8075
rect 27169 8041 27203 8075
rect 7849 7973 7883 8007
rect 9873 7973 9907 8007
rect 16129 7973 16163 8007
rect 19809 7973 19843 8007
rect 22753 7973 22787 8007
rect 1685 7905 1719 7939
rect 7481 7905 7515 7939
rect 9965 7905 9999 7939
rect 12817 7905 12851 7939
rect 18889 7905 18923 7939
rect 22385 7905 22419 7939
rect 1952 7837 1986 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6745 7837 6779 7871
rect 8585 7837 8619 7871
rect 10609 7837 10643 7871
rect 11253 7837 11287 7871
rect 13737 7837 13771 7871
rect 14289 7837 14323 7871
rect 14473 7837 14507 7871
rect 16037 7837 16071 7871
rect 16221 7837 16255 7871
rect 16405 7837 16439 7871
rect 17601 7837 17635 7871
rect 18705 7837 18739 7871
rect 20545 7837 20579 7871
rect 23489 7837 23523 7871
rect 24777 7837 24811 7871
rect 25789 7837 25823 7871
rect 6561 7769 6595 7803
rect 9505 7769 9539 7803
rect 11713 7769 11747 7803
rect 11929 7769 11963 7803
rect 12633 7769 12667 7803
rect 17417 7769 17451 7803
rect 18521 7769 18555 7803
rect 19441 7769 19475 7803
rect 20790 7769 20824 7803
rect 26034 7769 26068 7803
rect 4813 7701 4847 7735
rect 6101 7701 6135 7735
rect 7941 7701 7975 7735
rect 8401 7701 8435 7735
rect 11069 7701 11103 7735
rect 13553 7701 13587 7735
rect 14657 7701 14691 7735
rect 17785 7701 17819 7735
rect 19641 7701 19675 7735
rect 21925 7701 21959 7735
rect 22845 7701 22879 7735
rect 24593 7701 24627 7735
rect 3157 7497 3191 7531
rect 5917 7497 5951 7531
rect 7113 7497 7147 7531
rect 13277 7497 13311 7531
rect 17325 7497 17359 7531
rect 19007 7497 19041 7531
rect 20545 7497 20579 7531
rect 22201 7497 22235 7531
rect 22753 7497 22787 7531
rect 25973 7497 26007 7531
rect 12909 7429 12943 7463
rect 13125 7429 13159 7463
rect 18797 7429 18831 7463
rect 24838 7429 24872 7463
rect 1777 7361 1811 7395
rect 2033 7361 2067 7395
rect 3709 7361 3743 7395
rect 3976 7361 4010 7395
rect 5733 7361 5767 7395
rect 6837 7361 6871 7395
rect 7573 7361 7607 7395
rect 7757 7361 7791 7395
rect 9393 7361 9427 7395
rect 11161 7361 11195 7395
rect 11897 7361 11931 7395
rect 14453 7361 14487 7395
rect 16129 7361 16163 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 20729 7361 20763 7395
rect 21373 7361 21407 7395
rect 22109 7361 22143 7395
rect 22937 7361 22971 7395
rect 23581 7361 23615 7395
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 8217 7293 8251 7327
rect 9137 7293 9171 7327
rect 14197 7293 14231 7327
rect 17693 7293 17727 7327
rect 19625 7293 19659 7327
rect 24593 7293 24627 7327
rect 5089 7225 5123 7259
rect 8493 7225 8527 7259
rect 10517 7225 10551 7259
rect 17785 7225 17819 7259
rect 19165 7225 19199 7259
rect 19993 7225 20027 7259
rect 7665 7157 7699 7191
rect 8677 7157 8711 7191
rect 10977 7157 11011 7191
rect 11713 7157 11747 7191
rect 13093 7157 13127 7191
rect 15577 7157 15611 7191
rect 16221 7157 16255 7191
rect 18981 7157 19015 7191
rect 20085 7157 20119 7191
rect 21189 7157 21223 7191
rect 23397 7157 23431 7191
rect 4629 6953 4663 6987
rect 8401 6953 8435 6987
rect 9873 6953 9907 6987
rect 11989 6953 12023 6987
rect 12173 6953 12207 6987
rect 12633 6953 12667 6987
rect 14657 6953 14691 6987
rect 14841 6953 14875 6987
rect 15485 6953 15519 6987
rect 17601 6953 17635 6987
rect 20821 6953 20855 6987
rect 23121 6953 23155 6987
rect 4813 6885 4847 6919
rect 6745 6885 6779 6919
rect 15669 6885 15703 6919
rect 16497 6885 16531 6919
rect 17417 6885 17451 6919
rect 18429 6885 18463 6919
rect 19717 6885 19751 6919
rect 20637 6885 20671 6919
rect 13093 6817 13127 6851
rect 19901 6817 19935 6851
rect 20361 6817 20395 6851
rect 21741 6817 21775 6851
rect 1593 6749 1627 6783
rect 4261 6749 4295 6783
rect 4629 6749 4663 6783
rect 6377 6749 6411 6783
rect 7941 6749 7975 6783
rect 8585 6749 8619 6783
rect 10517 6749 10551 6783
rect 10665 6749 10699 6783
rect 10885 6749 10919 6783
rect 11023 6749 11057 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 13369 6749 13403 6783
rect 18061 6749 18095 6783
rect 21997 6749 22031 6783
rect 23765 6749 23799 6783
rect 24593 6749 24627 6783
rect 26433 6749 26467 6783
rect 26689 6749 26723 6783
rect 1838 6681 1872 6715
rect 5549 6681 5583 6715
rect 5733 6681 5767 6715
rect 9689 6681 9723 6715
rect 10793 6681 10827 6715
rect 11805 6681 11839 6715
rect 12021 6681 12055 6715
rect 14473 6681 14507 6715
rect 15301 6681 15335 6715
rect 15501 6681 15535 6715
rect 16129 6681 16163 6715
rect 17141 6681 17175 6715
rect 19441 6681 19475 6715
rect 24860 6681 24894 6715
rect 2973 6613 3007 6647
rect 5917 6613 5951 6647
rect 6837 6613 6871 6647
rect 7757 6613 7791 6647
rect 9889 6613 9923 6647
rect 10057 6613 10091 6647
rect 11161 6613 11195 6647
rect 13277 6613 13311 6647
rect 14673 6613 14707 6647
rect 16589 6613 16623 6647
rect 18521 6613 18555 6647
rect 23581 6613 23615 6647
rect 25973 6613 26007 6647
rect 27813 6613 27847 6647
rect 4077 6409 4111 6443
rect 4813 6409 4847 6443
rect 5457 6409 5491 6443
rect 9229 6409 9263 6443
rect 15393 6409 15427 6443
rect 17049 6409 17083 6443
rect 18337 6409 18371 6443
rect 26617 6409 26651 6443
rect 3709 6341 3743 6375
rect 3925 6341 3959 6375
rect 4721 6341 4755 6375
rect 8861 6341 8895 6375
rect 9077 6341 9111 6375
rect 10048 6341 10082 6375
rect 14105 6341 14139 6375
rect 15669 6341 15703 6375
rect 15899 6341 15933 6375
rect 17325 6341 17359 6375
rect 18245 6341 18279 6375
rect 23397 6341 23431 6375
rect 1777 6273 1811 6307
rect 2044 6273 2078 6307
rect 5365 6273 5399 6307
rect 5549 6273 5583 6307
rect 6745 6273 6779 6307
rect 7389 6273 7423 6307
rect 7665 6273 7699 6307
rect 11713 6273 11747 6307
rect 11806 6273 11840 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 12219 6273 12253 6307
rect 12909 6273 12943 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 17233 6273 17267 6307
rect 17417 6273 17451 6307
rect 17555 6273 17589 6307
rect 18889 6273 18923 6307
rect 19073 6273 19107 6307
rect 20269 6273 20303 6307
rect 20729 6273 20763 6307
rect 22293 6273 22327 6307
rect 24225 6273 24259 6307
rect 25493 6273 25527 6307
rect 8309 6205 8343 6239
rect 9781 6205 9815 6239
rect 14565 6205 14599 6239
rect 16037 6205 16071 6239
rect 17693 6205 17727 6239
rect 22017 6205 22051 6239
rect 25237 6205 25271 6239
rect 3157 6137 3191 6171
rect 11161 6137 11195 6171
rect 13093 6137 13127 6171
rect 14473 6137 14507 6171
rect 21005 6137 21039 6171
rect 21189 6137 21223 6171
rect 3893 6069 3927 6103
rect 6561 6069 6595 6103
rect 9045 6069 9079 6103
rect 12357 6069 12391 6103
rect 18889 6069 18923 6103
rect 20085 6069 20119 6103
rect 23489 6069 23523 6103
rect 24041 6069 24075 6103
rect 2513 5865 2547 5899
rect 3065 5865 3099 5899
rect 11897 5865 11931 5899
rect 12081 5865 12115 5899
rect 14473 5865 14507 5899
rect 23121 5865 23155 5899
rect 25973 5865 26007 5899
rect 3985 5797 4019 5831
rect 5549 5797 5583 5831
rect 7021 5797 7055 5831
rect 8585 5797 8619 5831
rect 10517 5797 10551 5831
rect 10977 5797 11011 5831
rect 14657 5797 14691 5831
rect 15393 5797 15427 5831
rect 17509 5797 17543 5831
rect 20821 5797 20855 5831
rect 23857 5797 23891 5831
rect 28365 5797 28399 5831
rect 1869 5729 1903 5763
rect 12909 5729 12943 5763
rect 13553 5729 13587 5763
rect 16497 5729 16531 5763
rect 26985 5729 27019 5763
rect 1685 5661 1719 5695
rect 3249 5661 3283 5695
rect 4261 5661 4295 5695
rect 4905 5661 4939 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 7849 5661 7883 5695
rect 8401 5661 8435 5695
rect 9137 5661 9171 5695
rect 11161 5661 11195 5695
rect 13093 5661 13127 5695
rect 15209 5661 15243 5695
rect 16037 5661 16071 5695
rect 16359 5661 16393 5695
rect 18613 5661 18647 5695
rect 19441 5661 19475 5695
rect 21741 5661 21775 5695
rect 24593 5661 24627 5695
rect 2421 5593 2455 5627
rect 3985 5593 4019 5627
rect 4721 5593 4755 5627
rect 6653 5593 6687 5627
rect 9382 5593 9416 5627
rect 11713 5593 11747 5627
rect 13185 5593 13219 5627
rect 13277 5593 13311 5627
rect 13415 5593 13449 5627
rect 14289 5593 14323 5627
rect 16129 5593 16163 5627
rect 16221 5593 16255 5627
rect 17141 5593 17175 5627
rect 18429 5593 18463 5627
rect 19686 5593 19720 5627
rect 21986 5593 22020 5627
rect 23581 5593 23615 5627
rect 24860 5593 24894 5627
rect 27230 5593 27264 5627
rect 4169 5525 4203 5559
rect 5089 5525 5123 5559
rect 5733 5525 5767 5559
rect 7113 5525 7147 5559
rect 7665 5525 7699 5559
rect 11913 5525 11947 5559
rect 14499 5525 14533 5559
rect 15853 5525 15887 5559
rect 17601 5525 17635 5559
rect 18797 5525 18831 5559
rect 24041 5525 24075 5559
rect 3157 5321 3191 5355
rect 3893 5321 3927 5355
rect 4261 5321 4295 5355
rect 9873 5321 9907 5355
rect 13277 5321 13311 5355
rect 15761 5321 15795 5355
rect 16865 5321 16899 5355
rect 18705 5321 18739 5355
rect 19993 5321 20027 5355
rect 22017 5321 22051 5355
rect 24041 5321 24075 5355
rect 24501 5321 24535 5355
rect 27261 5321 27295 5355
rect 2044 5253 2078 5287
rect 7389 5253 7423 5287
rect 8401 5253 8435 5287
rect 10379 5253 10413 5287
rect 12142 5253 12176 5287
rect 14626 5253 14660 5287
rect 17785 5253 17819 5287
rect 17995 5253 18029 5287
rect 22906 5253 22940 5287
rect 25482 5253 25516 5287
rect 1777 5185 1811 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 4997 5185 5031 5219
rect 5641 5185 5675 5219
rect 6653 5185 6687 5219
rect 10057 5185 10091 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 11161 5185 11195 5219
rect 13921 5185 13955 5219
rect 17049 5185 17083 5219
rect 17509 5185 17543 5219
rect 17693 5185 17727 5219
rect 17877 5185 17911 5219
rect 18889 5185 18923 5219
rect 19533 5185 19567 5219
rect 20177 5185 20211 5219
rect 20821 5185 20855 5219
rect 22201 5185 22235 5219
rect 22661 5185 22695 5219
rect 24685 5185 24719 5219
rect 27169 5185 27203 5219
rect 27353 5185 27387 5219
rect 5457 5117 5491 5151
rect 10517 5117 10551 5151
rect 11897 5117 11931 5151
rect 14381 5117 14415 5151
rect 18153 5117 18187 5151
rect 21281 5117 21315 5151
rect 25237 5117 25271 5151
rect 5825 5049 5859 5083
rect 8769 5049 8803 5083
rect 21097 5049 21131 5083
rect 4813 4981 4847 5015
rect 8861 4981 8895 5015
rect 10977 4981 11011 5015
rect 13737 4981 13771 5015
rect 19349 4981 19383 5015
rect 26617 4981 26651 5015
rect 3157 4777 3191 4811
rect 4445 4777 4479 4811
rect 4997 4777 5031 4811
rect 5641 4777 5675 4811
rect 10517 4777 10551 4811
rect 13737 4777 13771 4811
rect 27169 4777 27203 4811
rect 27721 4777 27755 4811
rect 8401 4709 8435 4743
rect 11805 4709 11839 4743
rect 13645 4709 13679 4743
rect 17325 4709 17359 4743
rect 18245 4709 18279 4743
rect 21557 4709 21591 4743
rect 22385 4709 22419 4743
rect 1777 4641 1811 4675
rect 6561 4641 6595 4675
rect 15761 4641 15795 4675
rect 17049 4641 17083 4675
rect 17969 4641 18003 4675
rect 18429 4641 18463 4675
rect 22017 4641 22051 4675
rect 22477 4641 22511 4675
rect 25789 4641 25823 4675
rect 2044 4573 2078 4607
rect 4905 4573 4939 4607
rect 5825 4573 5859 4607
rect 7021 4573 7055 4607
rect 9137 4573 9171 4607
rect 12633 4573 12667 4607
rect 13277 4573 13311 4607
rect 14473 4573 14507 4607
rect 15301 4573 15335 4607
rect 16037 4573 16071 4607
rect 19625 4573 19659 4607
rect 20177 4573 20211 4607
rect 23213 4573 23247 4607
rect 23489 4573 23523 4607
rect 24777 4573 24811 4607
rect 27629 4573 27663 4607
rect 27813 4573 27847 4607
rect 4077 4505 4111 4539
rect 4261 4505 4295 4539
rect 6377 4505 6411 4539
rect 7266 4505 7300 4539
rect 9382 4505 9416 4539
rect 11529 4505 11563 4539
rect 12449 4505 12483 4539
rect 14289 4505 14323 4539
rect 20422 4505 20456 4539
rect 26034 4505 26068 4539
rect 11989 4437 12023 4471
rect 12817 4437 12851 4471
rect 14657 4437 14691 4471
rect 15117 4437 15151 4471
rect 17509 4437 17543 4471
rect 19441 4437 19475 4471
rect 24593 4437 24627 4471
rect 15761 4233 15795 4267
rect 3893 4165 3927 4199
rect 9505 4165 9539 4199
rect 13737 4165 13771 4199
rect 14648 4165 14682 4199
rect 16865 4165 16899 4199
rect 17049 4165 17083 4199
rect 1777 4097 1811 4131
rect 2033 4097 2067 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 7093 4097 7127 4131
rect 8861 4097 8895 4131
rect 9321 4097 9355 4131
rect 18501 4097 18535 4131
rect 21189 4097 21223 4131
rect 22017 4097 22051 4131
rect 23204 4097 23238 4131
rect 24777 4097 24811 4131
rect 25033 4097 25067 4131
rect 27353 4097 27387 4131
rect 6837 4029 6871 4063
rect 10149 4029 10183 4063
rect 12173 4029 12207 4063
rect 12633 4029 12667 4063
rect 14381 4029 14415 4063
rect 18245 4029 18279 4063
rect 20085 4029 20119 4063
rect 20545 4029 20579 4063
rect 22937 4029 22971 4063
rect 3157 3961 3191 3995
rect 4813 3961 4847 3995
rect 5457 3961 5491 3995
rect 10517 3961 10551 3995
rect 12541 3961 12575 3995
rect 20453 3961 20487 3995
rect 21005 3961 21039 3995
rect 22293 3961 22327 3995
rect 4077 3893 4111 3927
rect 8217 3893 8251 3927
rect 8677 3893 8711 3927
rect 9689 3893 9723 3927
rect 10609 3893 10643 3927
rect 13829 3893 13863 3927
rect 17233 3893 17267 3927
rect 19625 3893 19659 3927
rect 22477 3893 22511 3927
rect 24317 3893 24351 3927
rect 26157 3893 26191 3927
rect 27169 3893 27203 3927
rect 3157 3689 3191 3723
rect 7021 3689 7055 3723
rect 12725 3689 12759 3723
rect 16957 3689 16991 3723
rect 18337 3689 18371 3723
rect 24041 3689 24075 3723
rect 28365 3689 28399 3723
rect 6561 3621 6595 3655
rect 8033 3621 8067 3655
rect 11805 3621 11839 3655
rect 17693 3621 17727 3655
rect 19809 3621 19843 3655
rect 20637 3621 20671 3655
rect 21557 3621 21591 3655
rect 1777 3553 1811 3587
rect 6193 3553 6227 3587
rect 15577 3553 15611 3587
rect 25145 3553 25179 3587
rect 26985 3553 27019 3587
rect 2044 3485 2078 3519
rect 5273 3485 5307 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6377 3485 6411 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7849 3485 7883 3519
rect 9229 3485 9263 3519
rect 10425 3485 10459 3519
rect 10681 3485 10715 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 15833 3485 15867 3519
rect 18521 3485 18555 3519
rect 22661 3485 22695 3519
rect 27241 3485 27275 3519
rect 4077 3417 4111 3451
rect 7665 3417 7699 3451
rect 9413 3417 9447 3451
rect 13369 3417 13403 3451
rect 14473 3417 14507 3451
rect 17417 3417 17451 3451
rect 19441 3417 19475 3451
rect 20361 3417 20395 3451
rect 21281 3417 21315 3451
rect 22906 3417 22940 3451
rect 25390 3417 25424 3451
rect 4169 3349 4203 3383
rect 5457 3349 5491 3383
rect 13737 3349 13771 3383
rect 14657 3349 14691 3383
rect 17877 3349 17911 3383
rect 19901 3349 19935 3383
rect 20821 3349 20855 3383
rect 21741 3349 21775 3383
rect 26525 3349 26559 3383
rect 1777 3145 1811 3179
rect 4353 3145 4387 3179
rect 7573 3145 7607 3179
rect 11989 3145 12023 3179
rect 14013 3145 14047 3179
rect 15853 3145 15887 3179
rect 20361 3145 20395 3179
rect 14718 3077 14752 3111
rect 17141 3077 17175 3111
rect 17325 3077 17359 3111
rect 17509 3077 17543 3111
rect 21005 3077 21039 3111
rect 1593 3009 1627 3043
rect 1777 3009 1811 3043
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 3240 3009 3274 3043
rect 4813 3009 4847 3043
rect 5365 3009 5399 3043
rect 5549 3009 5583 3043
rect 7757 3009 7791 3043
rect 8484 3009 8518 3043
rect 10425 3009 10459 3043
rect 11069 3009 11103 3043
rect 12173 3009 12207 3043
rect 12889 3009 12923 3043
rect 14473 3009 14507 3043
rect 18501 3009 18535 3043
rect 20545 3009 20579 3043
rect 22273 3009 22307 3043
rect 24665 3009 24699 3043
rect 26433 3009 26467 3043
rect 5089 2941 5123 2975
rect 6561 2941 6595 2975
rect 8217 2941 8251 2975
rect 12633 2941 12667 2975
rect 18245 2941 18279 2975
rect 22017 2941 22051 2975
rect 24409 2941 24443 2975
rect 2421 2873 2455 2907
rect 5365 2873 5399 2907
rect 6837 2873 6871 2907
rect 7021 2873 7055 2907
rect 9597 2873 9631 2907
rect 10241 2873 10275 2907
rect 21373 2873 21407 2907
rect 23397 2873 23431 2907
rect 25789 2873 25823 2907
rect 26249 2873 26283 2907
rect 10885 2805 10919 2839
rect 19625 2805 19659 2839
rect 21465 2805 21499 2839
rect 2973 2601 3007 2635
rect 8493 2601 8527 2635
rect 10977 2601 11011 2635
rect 12817 2601 12851 2635
rect 14289 2601 14323 2635
rect 17141 2601 17175 2635
rect 18245 2601 18279 2635
rect 24041 2601 24075 2635
rect 25973 2601 26007 2635
rect 4721 2533 4755 2567
rect 13553 2533 13587 2567
rect 19441 2533 19475 2567
rect 4353 2465 4387 2499
rect 22661 2465 22695 2499
rect 1593 2397 1627 2431
rect 1849 2397 1883 2431
rect 5273 2397 5307 2431
rect 7113 2397 7147 2431
rect 7380 2397 7414 2431
rect 9597 2397 9631 2431
rect 11437 2397 11471 2431
rect 11693 2397 11727 2431
rect 13737 2397 13771 2431
rect 14473 2397 14507 2431
rect 15301 2397 15335 2431
rect 15761 2397 15795 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 19625 2397 19659 2431
rect 20545 2397 20579 2431
rect 24593 2397 24627 2431
rect 26709 2397 26743 2431
rect 26965 2397 26999 2431
rect 5540 2329 5574 2363
rect 9864 2329 9898 2363
rect 16006 2329 16040 2363
rect 20801 2329 20835 2363
rect 22906 2329 22940 2363
rect 24860 2329 24894 2363
rect 4813 2261 4847 2295
rect 6653 2261 6687 2295
rect 15117 2261 15151 2295
rect 17601 2261 17635 2295
rect 21925 2261 21959 2295
rect 28089 2261 28123 2295
rect 3525 2057 3559 2091
rect 5825 2057 5859 2091
rect 9321 2057 9355 2091
rect 11161 2057 11195 2091
rect 26341 2057 26375 2091
rect 2412 1989 2446 2023
rect 4252 1989 4286 2023
rect 8186 1989 8220 2023
rect 12357 1989 12391 2023
rect 13522 1989 13556 2023
rect 15209 1989 15243 2023
rect 17110 1989 17144 2023
rect 18950 1989 18984 2023
rect 22262 1989 22296 2023
rect 2145 1921 2179 1955
rect 3985 1921 4019 1955
rect 6009 1921 6043 1955
rect 7021 1921 7055 1955
rect 7941 1921 7975 1955
rect 9781 1921 9815 1955
rect 10048 1921 10082 1955
rect 11897 1921 11931 1955
rect 13277 1921 13311 1955
rect 16313 1921 16347 1955
rect 16865 1921 16899 1955
rect 18705 1921 18739 1955
rect 20729 1921 20763 1955
rect 21373 1921 21407 1955
rect 24113 1921 24147 1955
rect 25881 1921 25915 1955
rect 26525 1921 26559 1955
rect 12817 1853 12851 1887
rect 15669 1853 15703 1887
rect 22017 1853 22051 1887
rect 23857 1853 23891 1887
rect 7389 1785 7423 1819
rect 12725 1785 12759 1819
rect 14657 1785 14691 1819
rect 15577 1785 15611 1819
rect 20545 1785 20579 1819
rect 23397 1785 23431 1819
rect 25697 1785 25731 1819
rect 5365 1717 5399 1751
rect 7481 1717 7515 1751
rect 11713 1717 11747 1751
rect 16129 1717 16163 1751
rect 18245 1717 18279 1751
rect 20085 1717 20119 1751
rect 21189 1717 21223 1751
rect 25237 1717 25271 1751
rect 5549 1513 5583 1547
rect 9781 1445 9815 1479
rect 14841 1445 14875 1479
rect 1593 1377 1627 1411
rect 4169 1377 4203 1411
rect 11713 1377 11747 1411
rect 14473 1377 14507 1411
rect 15761 1377 15795 1411
rect 24593 1377 24627 1411
rect 1860 1309 1894 1343
rect 6653 1309 6687 1343
rect 10425 1309 10459 1343
rect 10609 1309 10643 1343
rect 10793 1309 10827 1343
rect 13737 1309 13771 1343
rect 15577 1309 15611 1343
rect 17049 1309 17083 1343
rect 17509 1309 17543 1343
rect 19441 1309 19475 1343
rect 21465 1309 21499 1343
rect 22017 1309 22051 1343
rect 24041 1309 24075 1343
rect 24860 1309 24894 1343
rect 26617 1309 26651 1343
rect 27353 1309 27387 1343
rect 27629 1309 27663 1343
rect 4436 1241 4470 1275
rect 6920 1241 6954 1275
rect 9505 1241 9539 1275
rect 11958 1241 11992 1275
rect 15393 1241 15427 1275
rect 17754 1241 17788 1275
rect 19686 1241 19720 1275
rect 22262 1241 22296 1275
rect 2973 1173 3007 1207
rect 5917 1173 5951 1207
rect 8033 1173 8067 1207
rect 9965 1173 9999 1207
rect 13093 1173 13127 1207
rect 13553 1173 13587 1207
rect 14933 1173 14967 1207
rect 16865 1173 16899 1207
rect 18889 1173 18923 1207
rect 20821 1173 20855 1207
rect 21281 1173 21315 1207
rect 23397 1173 23431 1207
rect 23857 1173 23891 1207
rect 25973 1173 26007 1207
rect 26433 1173 26467 1207
rect 27169 1173 27203 1207
<< metal1 >>
rect 13998 33600 14004 33652
rect 14056 33640 14062 33652
rect 21174 33640 21180 33652
rect 14056 33612 21180 33640
rect 14056 33600 14062 33612
rect 21174 33600 21180 33612
rect 21232 33600 21238 33652
rect 12802 33532 12808 33584
rect 12860 33572 12866 33584
rect 19150 33572 19156 33584
rect 12860 33544 19156 33572
rect 12860 33532 12866 33544
rect 19150 33532 19156 33544
rect 19208 33532 19214 33584
rect 9214 33464 9220 33516
rect 9272 33504 9278 33516
rect 16758 33504 16764 33516
rect 9272 33476 16764 33504
rect 9272 33464 9278 33476
rect 16758 33464 16764 33476
rect 16816 33464 16822 33516
rect 17126 33464 17132 33516
rect 17184 33504 17190 33516
rect 25590 33504 25596 33516
rect 17184 33476 25596 33504
rect 17184 33464 17190 33476
rect 25590 33464 25596 33476
rect 25648 33464 25654 33516
rect 14458 33396 14464 33448
rect 14516 33436 14522 33448
rect 24946 33436 24952 33448
rect 14516 33408 24952 33436
rect 14516 33396 14522 33408
rect 24946 33396 24952 33408
rect 25004 33396 25010 33448
rect 7650 33328 7656 33380
rect 7708 33368 7714 33380
rect 16482 33368 16488 33380
rect 7708 33340 16488 33368
rect 7708 33328 7714 33340
rect 16482 33328 16488 33340
rect 16540 33328 16546 33380
rect 16850 33328 16856 33380
rect 16908 33368 16914 33380
rect 23382 33368 23388 33380
rect 16908 33340 23388 33368
rect 16908 33328 16914 33340
rect 23382 33328 23388 33340
rect 23440 33328 23446 33380
rect 4798 33260 4804 33312
rect 4856 33300 4862 33312
rect 6914 33300 6920 33312
rect 4856 33272 6920 33300
rect 4856 33260 4862 33272
rect 6914 33260 6920 33272
rect 6972 33300 6978 33312
rect 27338 33300 27344 33312
rect 6972 33272 27344 33300
rect 6972 33260 6978 33272
rect 27338 33260 27344 33272
rect 27396 33260 27402 33312
rect 10042 33192 10048 33244
rect 10100 33232 10106 33244
rect 10100 33204 17264 33232
rect 10100 33192 10106 33204
rect 10410 33124 10416 33176
rect 10468 33164 10474 33176
rect 17126 33164 17132 33176
rect 10468 33136 17132 33164
rect 10468 33124 10474 33136
rect 17126 33124 17132 33136
rect 17184 33124 17190 33176
rect 17236 33164 17264 33204
rect 17310 33192 17316 33244
rect 17368 33232 17374 33244
rect 27890 33232 27896 33244
rect 17368 33204 27896 33232
rect 17368 33192 17374 33204
rect 27890 33192 27896 33204
rect 27948 33192 27954 33244
rect 26786 33164 26792 33176
rect 17236 33136 26792 33164
rect 26786 33124 26792 33136
rect 26844 33124 26850 33176
rect 8478 33056 8484 33108
rect 8536 33096 8542 33108
rect 13814 33096 13820 33108
rect 8536 33068 13820 33096
rect 8536 33056 8542 33068
rect 13814 33056 13820 33068
rect 13872 33056 13878 33108
rect 14090 33056 14096 33108
rect 14148 33096 14154 33108
rect 19058 33096 19064 33108
rect 14148 33068 19064 33096
rect 14148 33056 14154 33068
rect 19058 33056 19064 33068
rect 19116 33056 19122 33108
rect 19150 33056 19156 33108
rect 19208 33096 19214 33108
rect 23474 33096 23480 33108
rect 19208 33068 23480 33096
rect 19208 33056 19214 33068
rect 23474 33056 23480 33068
rect 23532 33056 23538 33108
rect 13722 32988 13728 33040
rect 13780 33028 13786 33040
rect 23658 33028 23664 33040
rect 13780 33000 23664 33028
rect 13780 32988 13786 33000
rect 23658 32988 23664 33000
rect 23716 32988 23722 33040
rect 12526 32920 12532 32972
rect 12584 32960 12590 32972
rect 16390 32960 16396 32972
rect 12584 32932 16396 32960
rect 12584 32920 12590 32932
rect 16390 32920 16396 32932
rect 16448 32920 16454 32972
rect 16758 32920 16764 32972
rect 16816 32960 16822 32972
rect 27706 32960 27712 32972
rect 16816 32932 27712 32960
rect 16816 32920 16822 32932
rect 27706 32920 27712 32932
rect 27764 32920 27770 32972
rect 2314 32852 2320 32904
rect 2372 32892 2378 32904
rect 9490 32892 9496 32904
rect 2372 32864 9496 32892
rect 2372 32852 2378 32864
rect 9490 32852 9496 32864
rect 9548 32852 9554 32904
rect 13170 32852 13176 32904
rect 13228 32892 13234 32904
rect 16942 32892 16948 32904
rect 13228 32864 16948 32892
rect 13228 32852 13234 32864
rect 16942 32852 16948 32864
rect 17000 32852 17006 32904
rect 17126 32852 17132 32904
rect 17184 32892 17190 32904
rect 17184 32864 17448 32892
rect 17184 32852 17190 32864
rect 8294 32784 8300 32836
rect 8352 32824 8358 32836
rect 17310 32824 17316 32836
rect 8352 32796 17316 32824
rect 8352 32784 8358 32796
rect 17310 32784 17316 32796
rect 17368 32784 17374 32836
rect 17420 32824 17448 32864
rect 19242 32852 19248 32904
rect 19300 32892 19306 32904
rect 22922 32892 22928 32904
rect 19300 32864 22928 32892
rect 19300 32852 19306 32864
rect 22922 32852 22928 32864
rect 22980 32852 22986 32904
rect 21266 32824 21272 32836
rect 17420 32796 21272 32824
rect 21266 32784 21272 32796
rect 21324 32784 21330 32836
rect 26418 32824 26424 32836
rect 22066 32796 26424 32824
rect 11698 32716 11704 32768
rect 11756 32756 11762 32768
rect 14642 32756 14648 32768
rect 11756 32728 14648 32756
rect 11756 32716 11762 32728
rect 14642 32716 14648 32728
rect 14700 32716 14706 32768
rect 16482 32716 16488 32768
rect 16540 32756 16546 32768
rect 22066 32756 22094 32796
rect 26418 32784 26424 32796
rect 26476 32784 26482 32836
rect 16540 32728 22094 32756
rect 16540 32716 16546 32728
rect 22186 32716 22192 32768
rect 22244 32756 22250 32768
rect 25774 32756 25780 32768
rect 22244 32728 25780 32756
rect 22244 32716 22250 32728
rect 25774 32716 25780 32728
rect 25832 32716 25838 32768
rect 1104 32666 29048 32688
rect 1104 32614 7896 32666
rect 7948 32614 7960 32666
rect 8012 32614 8024 32666
rect 8076 32614 8088 32666
rect 8140 32614 8152 32666
rect 8204 32614 14842 32666
rect 14894 32614 14906 32666
rect 14958 32614 14970 32666
rect 15022 32614 15034 32666
rect 15086 32614 15098 32666
rect 15150 32614 21788 32666
rect 21840 32614 21852 32666
rect 21904 32614 21916 32666
rect 21968 32614 21980 32666
rect 22032 32614 22044 32666
rect 22096 32614 28734 32666
rect 28786 32614 28798 32666
rect 28850 32614 28862 32666
rect 28914 32614 28926 32666
rect 28978 32614 28990 32666
rect 29042 32614 29048 32666
rect 1104 32592 29048 32614
rect 2314 32512 2320 32564
rect 2372 32512 2378 32564
rect 4341 32555 4399 32561
rect 4341 32521 4353 32555
rect 4387 32552 4399 32555
rect 5166 32552 5172 32564
rect 4387 32524 5172 32552
rect 4387 32521 4399 32524
rect 4341 32515 4399 32521
rect 5166 32512 5172 32524
rect 5224 32552 5230 32564
rect 5997 32555 6055 32561
rect 5997 32552 6009 32555
rect 5224 32524 6009 32552
rect 5224 32512 5230 32524
rect 5997 32521 6009 32524
rect 6043 32552 6055 32555
rect 6917 32555 6975 32561
rect 6917 32552 6929 32555
rect 6043 32524 6929 32552
rect 6043 32521 6055 32524
rect 5997 32515 6055 32521
rect 6917 32521 6929 32524
rect 6963 32552 6975 32555
rect 7745 32555 7803 32561
rect 7745 32552 7757 32555
rect 6963 32524 7757 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 7745 32521 7757 32524
rect 7791 32552 7803 32555
rect 8573 32555 8631 32561
rect 8573 32552 8585 32555
rect 7791 32524 8585 32552
rect 7791 32521 7803 32524
rect 7745 32515 7803 32521
rect 8573 32521 8585 32524
rect 8619 32552 8631 32555
rect 9493 32555 9551 32561
rect 9493 32552 9505 32555
rect 8619 32524 9505 32552
rect 8619 32521 8631 32524
rect 8573 32515 8631 32521
rect 9493 32521 9505 32524
rect 9539 32552 9551 32555
rect 9950 32552 9956 32564
rect 9539 32524 9956 32552
rect 9539 32521 9551 32524
rect 9493 32515 9551 32521
rect 3326 32444 3332 32496
rect 3384 32484 3390 32496
rect 8386 32484 8392 32496
rect 3384 32456 8392 32484
rect 3384 32444 3390 32456
rect 8386 32444 8392 32456
rect 8444 32444 8450 32496
rect 2133 32419 2191 32425
rect 2133 32385 2145 32419
rect 2179 32416 2191 32419
rect 2866 32416 2872 32428
rect 2179 32388 2872 32416
rect 2179 32385 2191 32388
rect 2133 32379 2191 32385
rect 2866 32376 2872 32388
rect 2924 32376 2930 32428
rect 7006 32416 7012 32428
rect 2976 32388 7012 32416
rect 2406 32308 2412 32360
rect 2464 32308 2470 32360
rect 2682 32308 2688 32360
rect 2740 32348 2746 32360
rect 2976 32348 3004 32388
rect 7006 32376 7012 32388
rect 7064 32376 7070 32428
rect 8588 32425 8616 32515
rect 9950 32512 9956 32524
rect 10008 32552 10014 32564
rect 10321 32555 10379 32561
rect 10321 32552 10333 32555
rect 10008 32524 10333 32552
rect 10008 32512 10014 32524
rect 10321 32521 10333 32524
rect 10367 32552 10379 32555
rect 11149 32555 11207 32561
rect 11149 32552 11161 32555
rect 10367 32524 11161 32552
rect 10367 32521 10379 32524
rect 10321 32515 10379 32521
rect 11149 32521 11161 32524
rect 11195 32521 11207 32555
rect 11149 32515 11207 32521
rect 12406 32524 12664 32552
rect 9582 32444 9588 32496
rect 9640 32484 9646 32496
rect 9640 32456 11284 32484
rect 9640 32444 9646 32456
rect 7745 32419 7803 32425
rect 7745 32385 7757 32419
rect 7791 32416 7803 32419
rect 8573 32419 8631 32425
rect 8573 32416 8585 32419
rect 7791 32388 8585 32416
rect 7791 32385 7803 32388
rect 7745 32379 7803 32385
rect 8573 32385 8585 32388
rect 8619 32385 8631 32419
rect 11146 32416 11152 32428
rect 8573 32379 8631 32385
rect 8956 32388 11152 32416
rect 2740 32320 3004 32348
rect 2740 32308 2746 32320
rect 3050 32308 3056 32360
rect 3108 32308 3114 32360
rect 3234 32308 3240 32360
rect 3292 32348 3298 32360
rect 3421 32351 3479 32357
rect 3421 32348 3433 32351
rect 3292 32320 3433 32348
rect 3292 32308 3298 32320
rect 3421 32317 3433 32320
rect 3467 32348 3479 32351
rect 3973 32351 4031 32357
rect 3467 32320 3924 32348
rect 3467 32317 3479 32320
rect 3421 32311 3479 32317
rect 1857 32283 1915 32289
rect 1857 32249 1869 32283
rect 1903 32280 1915 32283
rect 3896 32280 3924 32320
rect 3973 32317 3985 32351
rect 4019 32348 4031 32351
rect 4798 32348 4804 32360
rect 4019 32320 4804 32348
rect 4019 32317 4031 32320
rect 3973 32311 4031 32317
rect 4798 32308 4804 32320
rect 4856 32308 4862 32360
rect 5629 32351 5687 32357
rect 5629 32317 5641 32351
rect 5675 32348 5687 32351
rect 6549 32351 6607 32357
rect 6549 32348 6561 32351
rect 5675 32320 6561 32348
rect 5675 32317 5687 32320
rect 5629 32311 5687 32317
rect 6549 32317 6561 32320
rect 6595 32348 6607 32351
rect 6638 32348 6644 32360
rect 6595 32320 6644 32348
rect 6595 32317 6607 32320
rect 6549 32311 6607 32317
rect 6638 32308 6644 32320
rect 6696 32308 6702 32360
rect 7377 32351 7435 32357
rect 7377 32317 7389 32351
rect 7423 32348 7435 32351
rect 7466 32348 7472 32360
rect 7423 32320 7472 32348
rect 7423 32317 7435 32320
rect 7377 32311 7435 32317
rect 7466 32308 7472 32320
rect 7524 32348 7530 32360
rect 8205 32351 8263 32357
rect 8205 32348 8217 32351
rect 7524 32320 8217 32348
rect 7524 32308 7530 32320
rect 8205 32317 8217 32320
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 4246 32280 4252 32292
rect 1903 32252 3556 32280
rect 3896 32252 4252 32280
rect 1903 32249 1915 32252
rect 1857 32243 1915 32249
rect 2866 32172 2872 32224
rect 2924 32172 2930 32224
rect 3142 32172 3148 32224
rect 3200 32212 3206 32224
rect 3421 32215 3479 32221
rect 3421 32212 3433 32215
rect 3200 32184 3433 32212
rect 3200 32172 3206 32184
rect 3421 32181 3433 32184
rect 3467 32181 3479 32215
rect 3528 32212 3556 32252
rect 4246 32240 4252 32252
rect 4304 32240 4310 32292
rect 4341 32283 4399 32289
rect 4341 32249 4353 32283
rect 4387 32280 4399 32283
rect 5166 32280 5172 32292
rect 4387 32252 5172 32280
rect 4387 32249 4399 32252
rect 4341 32243 4399 32249
rect 5166 32240 5172 32252
rect 5224 32240 5230 32292
rect 5997 32283 6055 32289
rect 5997 32249 6009 32283
rect 6043 32280 6055 32283
rect 6917 32283 6975 32289
rect 6917 32280 6929 32283
rect 6043 32252 6929 32280
rect 6043 32249 6055 32252
rect 5997 32243 6055 32249
rect 6917 32249 6929 32252
rect 6963 32280 6975 32283
rect 7190 32280 7196 32292
rect 6963 32252 7196 32280
rect 6963 32249 6975 32252
rect 6917 32243 6975 32249
rect 7190 32240 7196 32252
rect 7248 32240 7254 32292
rect 7742 32240 7748 32292
rect 7800 32280 7806 32292
rect 8956 32280 8984 32388
rect 11146 32376 11152 32388
rect 11204 32376 11210 32428
rect 9030 32308 9036 32360
rect 9088 32348 9094 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 9088 32320 9137 32348
rect 9088 32308 9094 32320
rect 9125 32317 9137 32320
rect 9171 32348 9183 32351
rect 9953 32351 10011 32357
rect 9953 32348 9965 32351
rect 9171 32320 9965 32348
rect 9171 32317 9183 32320
rect 9125 32311 9183 32317
rect 9953 32317 9965 32320
rect 9999 32348 10011 32351
rect 10781 32351 10839 32357
rect 10781 32348 10793 32351
rect 9999 32320 10793 32348
rect 9999 32317 10011 32320
rect 9953 32311 10011 32317
rect 10781 32317 10793 32320
rect 10827 32317 10839 32351
rect 11256 32348 11284 32456
rect 11606 32444 11612 32496
rect 11664 32484 11670 32496
rect 12406 32484 12434 32524
rect 11664 32456 12434 32484
rect 12636 32484 12664 32524
rect 14366 32512 14372 32564
rect 14424 32552 14430 32564
rect 22094 32552 22100 32564
rect 14424 32524 22100 32552
rect 14424 32512 14430 32524
rect 22094 32512 22100 32524
rect 22152 32552 22158 32564
rect 25866 32552 25872 32564
rect 22152 32524 22692 32552
rect 22152 32512 22158 32524
rect 12636 32456 20208 32484
rect 11664 32444 11670 32456
rect 11885 32419 11943 32425
rect 11885 32385 11897 32419
rect 11931 32416 11943 32419
rect 11931 32388 13400 32416
rect 11931 32385 11943 32388
rect 11885 32379 11943 32385
rect 12345 32351 12403 32357
rect 12345 32348 12357 32351
rect 11256 32320 12357 32348
rect 10781 32311 10839 32317
rect 12345 32317 12357 32320
rect 12391 32348 12403 32351
rect 13262 32348 13268 32360
rect 12391 32320 13268 32348
rect 12391 32317 12403 32320
rect 12345 32311 12403 32317
rect 13262 32308 13268 32320
rect 13320 32308 13326 32360
rect 13372 32348 13400 32388
rect 13630 32376 13636 32428
rect 13688 32416 13694 32428
rect 14277 32419 14335 32425
rect 14277 32416 14289 32419
rect 13688 32388 14289 32416
rect 13688 32376 13694 32388
rect 14277 32385 14289 32388
rect 14323 32416 14335 32419
rect 14366 32416 14372 32428
rect 14323 32388 14372 32416
rect 14323 32385 14335 32388
rect 14277 32379 14335 32385
rect 14366 32376 14372 32388
rect 14424 32376 14430 32428
rect 14458 32376 14464 32428
rect 14516 32376 14522 32428
rect 14642 32376 14648 32428
rect 14700 32416 14706 32428
rect 15177 32419 15235 32425
rect 15177 32416 15189 32419
rect 14700 32388 15189 32416
rect 14700 32376 14706 32388
rect 15177 32385 15189 32388
rect 15223 32385 15235 32419
rect 15177 32379 15235 32385
rect 16022 32376 16028 32428
rect 16080 32416 16086 32428
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16080 32388 17049 32416
rect 16080 32376 16086 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 17310 32376 17316 32428
rect 17368 32416 17374 32428
rect 17753 32419 17811 32425
rect 17753 32416 17765 32419
rect 17368 32388 17765 32416
rect 17368 32376 17374 32388
rect 17753 32385 17765 32388
rect 17799 32385 17811 32419
rect 17753 32379 17811 32385
rect 18046 32376 18052 32428
rect 18104 32416 18110 32428
rect 20053 32419 20111 32425
rect 20053 32416 20065 32419
rect 18104 32388 20065 32416
rect 18104 32376 18110 32388
rect 20053 32385 20065 32388
rect 20099 32385 20111 32419
rect 20180 32416 20208 32456
rect 20438 32444 20444 32496
rect 20496 32484 20502 32496
rect 20496 32456 22600 32484
rect 20496 32444 20502 32456
rect 22005 32419 22063 32425
rect 20180 32388 21128 32416
rect 20053 32379 20111 32385
rect 14182 32348 14188 32360
rect 13372 32320 14188 32348
rect 14182 32308 14188 32320
rect 14240 32308 14246 32360
rect 14550 32308 14556 32360
rect 14608 32348 14614 32360
rect 14921 32351 14979 32357
rect 14921 32348 14933 32351
rect 14608 32320 14933 32348
rect 14608 32308 14614 32320
rect 14921 32317 14933 32320
rect 14967 32317 14979 32351
rect 14921 32311 14979 32317
rect 16666 32308 16672 32360
rect 16724 32348 16730 32360
rect 17497 32351 17555 32357
rect 17497 32348 17509 32351
rect 16724 32320 17509 32348
rect 16724 32308 16730 32320
rect 17497 32317 17509 32320
rect 17543 32317 17555 32351
rect 17497 32311 17555 32317
rect 19426 32308 19432 32360
rect 19484 32348 19490 32360
rect 19797 32351 19855 32357
rect 19797 32348 19809 32351
rect 19484 32320 19809 32348
rect 19484 32308 19490 32320
rect 19797 32317 19809 32320
rect 19843 32317 19855 32351
rect 19797 32311 19855 32317
rect 7800 32252 8984 32280
rect 9493 32283 9551 32289
rect 7800 32240 7806 32252
rect 9493 32249 9505 32283
rect 9539 32280 9551 32283
rect 10134 32280 10140 32292
rect 9539 32252 10140 32280
rect 9539 32249 9551 32252
rect 9493 32243 9551 32249
rect 10134 32240 10140 32252
rect 10192 32280 10198 32292
rect 10321 32283 10379 32289
rect 10321 32280 10333 32283
rect 10192 32252 10333 32280
rect 10192 32240 10198 32252
rect 10321 32249 10333 32252
rect 10367 32280 10379 32283
rect 11149 32283 11207 32289
rect 11149 32280 11161 32283
rect 10367 32252 11161 32280
rect 10367 32249 10379 32252
rect 10321 32243 10379 32249
rect 11149 32249 11161 32252
rect 11195 32280 11207 32283
rect 12434 32280 12440 32292
rect 11195 32252 12440 32280
rect 11195 32249 11207 32252
rect 11149 32243 11207 32249
rect 12434 32240 12440 32252
rect 12492 32240 12498 32292
rect 12526 32240 12532 32292
rect 12584 32280 12590 32292
rect 12621 32283 12679 32289
rect 12621 32280 12633 32283
rect 12584 32252 12633 32280
rect 12584 32240 12590 32252
rect 12621 32249 12633 32252
rect 12667 32249 12679 32283
rect 12621 32243 12679 32249
rect 12728 32252 12940 32280
rect 11606 32212 11612 32224
rect 3528 32184 11612 32212
rect 3421 32175 3479 32181
rect 11606 32172 11612 32184
rect 11664 32172 11670 32224
rect 11701 32215 11759 32221
rect 11701 32181 11713 32215
rect 11747 32212 11759 32215
rect 12728 32212 12756 32252
rect 11747 32184 12756 32212
rect 11747 32181 11759 32184
rect 11701 32175 11759 32181
rect 12802 32172 12808 32224
rect 12860 32172 12866 32224
rect 12912 32212 12940 32252
rect 13538 32240 13544 32292
rect 13596 32240 13602 32292
rect 14826 32280 14832 32292
rect 13648 32252 14832 32280
rect 13648 32212 13676 32252
rect 14826 32240 14832 32252
rect 14884 32240 14890 32292
rect 16206 32240 16212 32292
rect 16264 32280 16270 32292
rect 16853 32283 16911 32289
rect 16264 32252 16436 32280
rect 16264 32240 16270 32252
rect 12912 32184 13676 32212
rect 13722 32172 13728 32224
rect 13780 32172 13786 32224
rect 13906 32172 13912 32224
rect 13964 32212 13970 32224
rect 16301 32215 16359 32221
rect 16301 32212 16313 32215
rect 13964 32184 16313 32212
rect 13964 32172 13970 32184
rect 16301 32181 16313 32184
rect 16347 32181 16359 32215
rect 16408 32212 16436 32252
rect 16853 32249 16865 32283
rect 16899 32280 16911 32283
rect 17402 32280 17408 32292
rect 16899 32252 17408 32280
rect 16899 32249 16911 32252
rect 16853 32243 16911 32249
rect 17402 32240 17408 32252
rect 17460 32240 17466 32292
rect 21100 32280 21128 32388
rect 22005 32385 22017 32419
rect 22051 32416 22063 32419
rect 22094 32416 22100 32428
rect 22051 32388 22100 32416
rect 22051 32385 22063 32388
rect 22005 32379 22063 32385
rect 22094 32376 22100 32388
rect 22152 32376 22158 32428
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 22572 32348 22600 32456
rect 22664 32425 22692 32524
rect 22756 32524 25872 32552
rect 22649 32419 22707 32425
rect 22649 32385 22661 32419
rect 22695 32385 22707 32419
rect 22649 32379 22707 32385
rect 22756 32348 22784 32524
rect 25866 32512 25872 32524
rect 25924 32512 25930 32564
rect 25130 32484 25136 32496
rect 22848 32456 25136 32484
rect 22848 32425 22876 32456
rect 25130 32444 25136 32456
rect 25188 32444 25194 32496
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 23474 32376 23480 32428
rect 23532 32376 23538 32428
rect 25869 32419 25927 32425
rect 25869 32385 25881 32419
rect 25915 32416 25927 32419
rect 25958 32416 25964 32428
rect 25915 32388 25964 32416
rect 25915 32385 25927 32388
rect 25869 32379 25927 32385
rect 25958 32376 25964 32388
rect 26016 32376 26022 32428
rect 26053 32419 26111 32425
rect 26053 32385 26065 32419
rect 26099 32416 26111 32419
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 26099 32388 27353 32416
rect 26099 32385 26111 32388
rect 26053 32379 26111 32385
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27801 32419 27859 32425
rect 27801 32385 27813 32419
rect 27847 32385 27859 32419
rect 27801 32379 27859 32385
rect 22572 32320 22784 32348
rect 23566 32308 23572 32360
rect 23624 32348 23630 32360
rect 25409 32351 25467 32357
rect 25409 32348 25421 32351
rect 23624 32320 25421 32348
rect 23624 32308 23630 32320
rect 25409 32317 25421 32320
rect 25455 32317 25467 32351
rect 25409 32311 25467 32317
rect 27816 32280 27844 32379
rect 28074 32280 28080 32292
rect 21100 32252 27844 32280
rect 27908 32252 28080 32280
rect 18877 32215 18935 32221
rect 18877 32212 18889 32215
rect 16408 32184 18889 32212
rect 16301 32175 16359 32181
rect 18877 32181 18889 32184
rect 18923 32181 18935 32215
rect 18877 32175 18935 32181
rect 19610 32172 19616 32224
rect 19668 32212 19674 32224
rect 20438 32212 20444 32224
rect 19668 32184 20444 32212
rect 19668 32172 19674 32184
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 21174 32172 21180 32224
rect 21232 32172 21238 32224
rect 21266 32172 21272 32224
rect 21324 32212 21330 32224
rect 23293 32215 23351 32221
rect 23293 32212 23305 32215
rect 21324 32184 23305 32212
rect 21324 32172 21330 32184
rect 23293 32181 23305 32184
rect 23339 32181 23351 32215
rect 23293 32175 23351 32181
rect 24765 32215 24823 32221
rect 24765 32181 24777 32215
rect 24811 32212 24823 32215
rect 27908 32212 27936 32252
rect 28074 32240 28080 32252
rect 28132 32240 28138 32292
rect 24811 32184 27936 32212
rect 24811 32181 24823 32184
rect 24765 32175 24823 32181
rect 27982 32172 27988 32224
rect 28040 32172 28046 32224
rect 1104 32122 28888 32144
rect 1104 32070 4423 32122
rect 4475 32070 4487 32122
rect 4539 32070 4551 32122
rect 4603 32070 4615 32122
rect 4667 32070 4679 32122
rect 4731 32070 11369 32122
rect 11421 32070 11433 32122
rect 11485 32070 11497 32122
rect 11549 32070 11561 32122
rect 11613 32070 11625 32122
rect 11677 32070 18315 32122
rect 18367 32070 18379 32122
rect 18431 32070 18443 32122
rect 18495 32070 18507 32122
rect 18559 32070 18571 32122
rect 18623 32070 25261 32122
rect 25313 32070 25325 32122
rect 25377 32070 25389 32122
rect 25441 32070 25453 32122
rect 25505 32070 25517 32122
rect 25569 32070 28888 32122
rect 1104 32048 28888 32070
rect 3326 31968 3332 32020
rect 3384 31968 3390 32020
rect 3418 31968 3424 32020
rect 3476 32008 3482 32020
rect 27982 32008 27988 32020
rect 3476 31980 27988 32008
rect 3476 31968 3482 31980
rect 27982 31968 27988 31980
rect 28040 31968 28046 32020
rect 2133 31943 2191 31949
rect 2133 31909 2145 31943
rect 2179 31940 2191 31943
rect 4246 31940 4252 31952
rect 2179 31912 4252 31940
rect 2179 31909 2191 31912
rect 2133 31903 2191 31909
rect 4246 31900 4252 31912
rect 4304 31900 4310 31952
rect 4338 31900 4344 31952
rect 4396 31940 4402 31952
rect 4433 31943 4491 31949
rect 4433 31940 4445 31943
rect 4396 31912 4445 31940
rect 4396 31900 4402 31912
rect 4433 31909 4445 31912
rect 4479 31940 4491 31943
rect 5258 31940 5264 31952
rect 4479 31912 5264 31940
rect 4479 31909 4491 31912
rect 4433 31903 4491 31909
rect 5258 31900 5264 31912
rect 5316 31900 5322 31952
rect 7742 31900 7748 31952
rect 7800 31900 7806 31952
rect 7837 31943 7895 31949
rect 7837 31909 7849 31943
rect 7883 31940 7895 31943
rect 8294 31940 8300 31952
rect 7883 31912 8300 31940
rect 7883 31909 7895 31912
rect 7837 31903 7895 31909
rect 8294 31900 8300 31912
rect 8352 31900 8358 31952
rect 8478 31900 8484 31952
rect 8536 31900 8542 31952
rect 9953 31943 10011 31949
rect 9953 31909 9965 31943
rect 9999 31940 10011 31943
rect 10594 31940 10600 31952
rect 9999 31912 10600 31940
rect 9999 31909 10011 31912
rect 9953 31903 10011 31909
rect 10594 31900 10600 31912
rect 10652 31900 10658 31952
rect 12621 31943 12679 31949
rect 12621 31909 12633 31943
rect 12667 31940 12679 31943
rect 13170 31940 13176 31952
rect 12667 31912 13176 31940
rect 12667 31909 12679 31912
rect 12621 31903 12679 31909
rect 13170 31900 13176 31912
rect 13228 31900 13234 31952
rect 13541 31943 13599 31949
rect 13541 31909 13553 31943
rect 13587 31909 13599 31943
rect 13541 31903 13599 31909
rect 2590 31832 2596 31884
rect 2648 31832 2654 31884
rect 2682 31832 2688 31884
rect 2740 31832 2746 31884
rect 2866 31832 2872 31884
rect 2924 31872 2930 31884
rect 10502 31872 10508 31884
rect 2924 31844 10508 31872
rect 2924 31832 2930 31844
rect 10502 31832 10508 31844
rect 10560 31832 10566 31884
rect 3237 31807 3295 31813
rect 3237 31773 3249 31807
rect 3283 31804 3295 31807
rect 3970 31804 3976 31816
rect 3283 31776 3976 31804
rect 3283 31773 3295 31776
rect 3237 31767 3295 31773
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31804 4123 31807
rect 4154 31804 4160 31816
rect 4111 31776 4160 31804
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 3050 31696 3056 31748
rect 3108 31736 3114 31748
rect 4080 31736 4108 31767
rect 4154 31764 4160 31776
rect 4212 31804 4218 31816
rect 4893 31807 4951 31813
rect 4893 31804 4905 31807
rect 4212 31776 4905 31804
rect 4212 31764 4218 31776
rect 4893 31773 4905 31776
rect 4939 31773 4951 31807
rect 4893 31767 4951 31773
rect 5718 31764 5724 31816
rect 5776 31764 5782 31816
rect 6086 31764 6092 31816
rect 6144 31764 6150 31816
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 6917 31807 6975 31813
rect 6917 31773 6929 31807
rect 6963 31773 6975 31807
rect 6917 31767 6975 31773
rect 7377 31807 7435 31813
rect 7377 31773 7389 31807
rect 7423 31804 7435 31807
rect 7558 31804 7564 31816
rect 7423 31776 7564 31804
rect 7423 31773 7435 31776
rect 7377 31767 7435 31773
rect 3108 31708 4108 31736
rect 6104 31736 6132 31764
rect 6932 31736 6960 31767
rect 7558 31764 7564 31776
rect 7616 31804 7622 31816
rect 7616 31776 8248 31804
rect 7616 31764 7622 31776
rect 6104 31708 6960 31736
rect 8220 31736 8248 31776
rect 8294 31764 8300 31816
rect 8352 31764 8358 31816
rect 8404 31776 9536 31804
rect 8404 31736 8432 31776
rect 8220 31708 8432 31736
rect 9508 31736 9536 31776
rect 10042 31764 10048 31816
rect 10100 31764 10106 31816
rect 10410 31764 10416 31816
rect 10468 31804 10474 31816
rect 10468 31776 10640 31804
rect 10468 31764 10474 31776
rect 9582 31736 9588 31748
rect 9508 31708 9588 31736
rect 3108 31696 3114 31708
rect 9582 31696 9588 31708
rect 9640 31696 9646 31748
rect 2593 31671 2651 31677
rect 2593 31637 2605 31671
rect 2639 31668 2651 31671
rect 4338 31668 4344 31680
rect 2639 31640 4344 31668
rect 2639 31637 2651 31640
rect 2593 31631 2651 31637
rect 4338 31628 4344 31640
rect 4396 31628 4402 31680
rect 4433 31671 4491 31677
rect 4433 31637 4445 31671
rect 4479 31668 4491 31671
rect 4522 31668 4528 31680
rect 4479 31640 4528 31668
rect 4479 31637 4491 31640
rect 4433 31631 4491 31637
rect 4522 31628 4528 31640
rect 4580 31628 4586 31680
rect 5166 31628 5172 31680
rect 5224 31668 5230 31680
rect 10060 31677 10088 31764
rect 10612 31736 10640 31776
rect 10686 31764 10692 31816
rect 10744 31764 10750 31816
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31804 12863 31807
rect 13446 31804 13452 31816
rect 12851 31776 13452 31804
rect 12851 31773 12863 31776
rect 12805 31767 12863 31773
rect 13446 31764 13452 31776
rect 13504 31764 13510 31816
rect 10934 31739 10992 31745
rect 10934 31736 10946 31739
rect 10612 31708 10946 31736
rect 10934 31705 10946 31708
rect 10980 31705 10992 31739
rect 10934 31699 10992 31705
rect 13262 31696 13268 31748
rect 13320 31696 13326 31748
rect 13556 31736 13584 31903
rect 17586 31900 17592 31952
rect 17644 31940 17650 31952
rect 17865 31943 17923 31949
rect 17865 31940 17877 31943
rect 17644 31912 17877 31940
rect 17644 31900 17650 31912
rect 17865 31909 17877 31912
rect 17911 31909 17923 31943
rect 17865 31903 17923 31909
rect 18230 31900 18236 31952
rect 18288 31940 18294 31952
rect 18693 31943 18751 31949
rect 18693 31940 18705 31943
rect 18288 31912 18705 31940
rect 18288 31900 18294 31912
rect 18693 31909 18705 31912
rect 18739 31909 18751 31943
rect 18693 31903 18751 31909
rect 20806 31900 20812 31952
rect 20864 31900 20870 31952
rect 22922 31900 22928 31952
rect 22980 31900 22986 31952
rect 23492 31912 23888 31940
rect 13725 31875 13783 31881
rect 13725 31841 13737 31875
rect 13771 31872 13783 31875
rect 14090 31872 14096 31884
rect 13771 31844 14096 31872
rect 13771 31841 13783 31844
rect 13725 31835 13783 31841
rect 14090 31832 14096 31844
rect 14148 31832 14154 31884
rect 23492 31872 23520 31912
rect 23658 31872 23664 31884
rect 17512 31844 19564 31872
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31804 14335 31807
rect 15746 31804 15752 31816
rect 14323 31776 15752 31804
rect 14323 31773 14335 31776
rect 14277 31767 14335 31773
rect 15746 31764 15752 31776
rect 15804 31764 15810 31816
rect 16474 31807 16532 31813
rect 16474 31773 16486 31807
rect 16520 31773 16532 31807
rect 16474 31767 16532 31773
rect 14182 31736 14188 31748
rect 13556 31708 14188 31736
rect 14182 31696 14188 31708
rect 14240 31736 14246 31748
rect 16298 31736 16304 31748
rect 14240 31708 16304 31736
rect 14240 31696 14246 31708
rect 16298 31696 16304 31708
rect 16356 31696 16362 31748
rect 16500 31736 16528 31767
rect 17126 31764 17132 31816
rect 17184 31804 17190 31816
rect 17512 31804 17540 31844
rect 17184 31776 17540 31804
rect 18325 31807 18383 31813
rect 17184 31764 17190 31776
rect 18325 31773 18337 31807
rect 18371 31773 18383 31807
rect 18325 31767 18383 31773
rect 16574 31736 16580 31748
rect 16500 31708 16580 31736
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 16752 31739 16810 31745
rect 16752 31705 16764 31739
rect 16798 31736 16810 31739
rect 16850 31736 16856 31748
rect 16798 31708 16856 31736
rect 16798 31705 16810 31708
rect 16752 31699 16810 31705
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 17678 31696 17684 31748
rect 17736 31736 17742 31748
rect 18340 31736 18368 31767
rect 18414 31764 18420 31816
rect 18472 31804 18478 31816
rect 18472 31776 19380 31804
rect 18472 31764 18478 31776
rect 17736 31708 18368 31736
rect 19352 31736 19380 31776
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 19536 31804 19564 31844
rect 20456 31844 21680 31872
rect 20456 31804 20484 31844
rect 19536 31776 20484 31804
rect 20916 31776 21496 31804
rect 19674 31739 19732 31745
rect 19674 31736 19686 31739
rect 19352 31708 19686 31736
rect 17736 31696 17742 31708
rect 19674 31705 19686 31708
rect 19720 31705 19732 31739
rect 19674 31699 19732 31705
rect 5261 31671 5319 31677
rect 5261 31668 5273 31671
rect 5224 31640 5273 31668
rect 5224 31628 5230 31640
rect 5261 31637 5273 31640
rect 5307 31668 5319 31671
rect 6089 31671 6147 31677
rect 6089 31668 6101 31671
rect 5307 31640 6101 31668
rect 5307 31637 5319 31640
rect 5261 31631 5319 31637
rect 6089 31637 6101 31640
rect 6135 31668 6147 31671
rect 6917 31671 6975 31677
rect 6917 31668 6929 31671
rect 6135 31640 6929 31668
rect 6135 31637 6147 31640
rect 6089 31631 6147 31637
rect 6917 31637 6929 31640
rect 6963 31637 6975 31671
rect 6917 31631 6975 31637
rect 10045 31671 10103 31677
rect 10045 31637 10057 31671
rect 10091 31637 10103 31671
rect 10045 31631 10103 31637
rect 10502 31628 10508 31680
rect 10560 31668 10566 31680
rect 12069 31671 12127 31677
rect 12069 31668 12081 31671
rect 10560 31640 12081 31668
rect 10560 31628 10566 31640
rect 12069 31637 12081 31640
rect 12115 31637 12127 31671
rect 12069 31631 12127 31637
rect 13538 31628 13544 31680
rect 13596 31668 13602 31680
rect 15286 31668 15292 31680
rect 13596 31640 15292 31668
rect 13596 31628 13602 31640
rect 15286 31628 15292 31640
rect 15344 31628 15350 31680
rect 15562 31628 15568 31680
rect 15620 31628 15626 31680
rect 17770 31628 17776 31680
rect 17828 31668 17834 31680
rect 18693 31671 18751 31677
rect 18693 31668 18705 31671
rect 17828 31640 18705 31668
rect 17828 31628 17834 31640
rect 18693 31637 18705 31640
rect 18739 31637 18751 31671
rect 18693 31631 18751 31637
rect 18782 31628 18788 31680
rect 18840 31668 18846 31680
rect 20916 31668 20944 31776
rect 21468 31736 21496 31776
rect 21542 31764 21548 31816
rect 21600 31764 21606 31816
rect 21652 31804 21680 31844
rect 22572 31844 23520 31872
rect 23584 31844 23664 31872
rect 22572 31804 22600 31844
rect 23584 31813 23612 31844
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 23860 31872 23888 31912
rect 25866 31900 25872 31952
rect 25924 31940 25930 31952
rect 25961 31943 26019 31949
rect 25961 31940 25973 31943
rect 25924 31912 25973 31940
rect 25924 31900 25930 31912
rect 25961 31909 25973 31912
rect 26007 31909 26019 31943
rect 25961 31903 26019 31909
rect 26418 31900 26424 31952
rect 26476 31900 26482 31952
rect 26510 31900 26516 31952
rect 26568 31940 26574 31952
rect 27249 31943 27307 31949
rect 27249 31940 27261 31943
rect 26568 31912 27261 31940
rect 26568 31900 26574 31912
rect 27249 31909 27261 31912
rect 27295 31909 27307 31943
rect 27249 31903 27307 31909
rect 27706 31900 27712 31952
rect 27764 31900 27770 31952
rect 23860 31844 24716 31872
rect 23569 31807 23627 31813
rect 21652 31776 22600 31804
rect 22664 31776 23336 31804
rect 21790 31739 21848 31745
rect 21790 31736 21802 31739
rect 21468 31708 21802 31736
rect 21790 31705 21802 31708
rect 21836 31705 21848 31739
rect 22664 31736 22692 31776
rect 21790 31699 21848 31705
rect 22066 31708 22692 31736
rect 23308 31736 23336 31776
rect 23569 31773 23581 31807
rect 23615 31773 23627 31807
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 23860 31780 24593 31804
rect 23569 31767 23627 31773
rect 23676 31776 24593 31780
rect 23676 31752 23888 31776
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 24688 31804 24716 31844
rect 26326 31804 26332 31816
rect 24688 31776 26332 31804
rect 24581 31767 24639 31773
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 26418 31764 26424 31816
rect 26476 31764 26482 31816
rect 26602 31764 26608 31816
rect 26660 31804 26666 31816
rect 26660 31776 27292 31804
rect 26660 31764 26666 31776
rect 23676 31736 23704 31752
rect 23308 31708 23704 31736
rect 18840 31640 20944 31668
rect 18840 31628 18846 31640
rect 21542 31628 21548 31680
rect 21600 31668 21606 31680
rect 22066 31668 22094 31708
rect 23934 31696 23940 31748
rect 23992 31736 23998 31748
rect 24826 31739 24884 31745
rect 24826 31736 24838 31739
rect 23992 31708 24838 31736
rect 23992 31696 23998 31708
rect 24826 31705 24838 31708
rect 24872 31705 24884 31739
rect 27264 31736 27292 31776
rect 27338 31764 27344 31816
rect 27396 31804 27402 31816
rect 27709 31807 27767 31813
rect 27709 31804 27721 31807
rect 27396 31776 27721 31804
rect 27396 31764 27402 31776
rect 27709 31773 27721 31776
rect 27755 31773 27767 31807
rect 27893 31807 27951 31813
rect 27893 31804 27905 31807
rect 27709 31767 27767 31773
rect 27816 31776 27905 31804
rect 27816 31736 27844 31776
rect 27893 31773 27905 31776
rect 27939 31773 27951 31807
rect 27893 31767 27951 31773
rect 27264 31708 27844 31736
rect 24826 31699 24884 31705
rect 21600 31640 22094 31668
rect 21600 31628 21606 31640
rect 23382 31628 23388 31680
rect 23440 31628 23446 31680
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 2041 31467 2099 31473
rect 2041 31433 2053 31467
rect 2087 31464 2099 31467
rect 3142 31464 3148 31476
rect 2087 31436 3148 31464
rect 2087 31433 2099 31436
rect 2041 31427 2099 31433
rect 3142 31424 3148 31436
rect 3200 31464 3206 31476
rect 4522 31464 4528 31476
rect 3200 31436 4528 31464
rect 3200 31424 3206 31436
rect 4522 31424 4528 31436
rect 4580 31464 4586 31476
rect 5166 31464 5172 31476
rect 4580 31436 5172 31464
rect 4580 31424 4586 31436
rect 5166 31424 5172 31436
rect 5224 31464 5230 31476
rect 5997 31467 6055 31473
rect 5997 31464 6009 31467
rect 5224 31436 6009 31464
rect 5224 31424 5230 31436
rect 5997 31433 6009 31436
rect 6043 31464 6055 31467
rect 7009 31467 7067 31473
rect 7009 31464 7021 31467
rect 6043 31436 7021 31464
rect 6043 31433 6055 31436
rect 5997 31427 6055 31433
rect 7009 31433 7021 31436
rect 7055 31464 7067 31467
rect 7834 31464 7840 31476
rect 7055 31436 7840 31464
rect 7055 31433 7067 31436
rect 7009 31427 7067 31433
rect 7834 31424 7840 31436
rect 7892 31464 7898 31476
rect 8665 31467 8723 31473
rect 8665 31464 8677 31467
rect 7892 31436 8677 31464
rect 7892 31424 7898 31436
rect 8665 31433 8677 31436
rect 8711 31433 8723 31467
rect 8665 31427 8723 31433
rect 9030 31424 9036 31476
rect 9088 31464 9094 31476
rect 10965 31467 11023 31473
rect 9088 31436 10272 31464
rect 9088 31424 9094 31436
rect 7190 31396 7196 31408
rect 7024 31368 7196 31396
rect 2498 31288 2504 31340
rect 2556 31288 2562 31340
rect 4798 31288 4804 31340
rect 4856 31288 4862 31340
rect 5166 31288 5172 31340
rect 5224 31288 5230 31340
rect 5997 31331 6055 31337
rect 5997 31297 6009 31331
rect 6043 31328 6055 31331
rect 6086 31328 6092 31340
rect 6043 31300 6092 31328
rect 6043 31297 6055 31300
rect 5997 31291 6055 31297
rect 6086 31288 6092 31300
rect 6144 31288 6150 31340
rect 7024 31337 7052 31368
rect 7190 31356 7196 31368
rect 7248 31396 7254 31408
rect 10134 31396 10140 31408
rect 7248 31368 10140 31396
rect 7248 31356 7254 31368
rect 10134 31356 10140 31368
rect 10192 31356 10198 31408
rect 7009 31331 7067 31337
rect 7009 31297 7021 31331
rect 7055 31297 7067 31331
rect 9030 31328 9036 31340
rect 7009 31291 7067 31297
rect 7392 31300 9036 31328
rect 1673 31263 1731 31269
rect 1673 31229 1685 31263
rect 1719 31260 1731 31263
rect 3050 31260 3056 31272
rect 1719 31232 3056 31260
rect 1719 31229 1731 31232
rect 1673 31223 1731 31229
rect 3050 31220 3056 31232
rect 3108 31220 3114 31272
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31260 5687 31263
rect 5718 31260 5724 31272
rect 5675 31232 5724 31260
rect 5675 31229 5687 31232
rect 5629 31223 5687 31229
rect 5718 31220 5724 31232
rect 5776 31220 5782 31272
rect 6454 31220 6460 31272
rect 6512 31260 6518 31272
rect 6638 31260 6644 31272
rect 6512 31232 6644 31260
rect 6512 31220 6518 31232
rect 6638 31220 6644 31232
rect 6696 31260 6702 31272
rect 7392 31260 7420 31300
rect 9030 31288 9036 31300
rect 9088 31288 9094 31340
rect 9398 31337 9404 31340
rect 9392 31291 9404 31337
rect 9398 31288 9404 31291
rect 9456 31288 9462 31340
rect 6696 31232 7420 31260
rect 6696 31220 6702 31232
rect 7466 31220 7472 31272
rect 7524 31260 7530 31272
rect 8297 31263 8355 31269
rect 8297 31260 8309 31263
rect 7524 31232 8309 31260
rect 7524 31220 7530 31232
rect 8297 31229 8309 31232
rect 8343 31229 8355 31263
rect 8297 31223 8355 31229
rect 9122 31220 9128 31272
rect 9180 31220 9186 31272
rect 10244 31260 10272 31436
rect 10965 31433 10977 31467
rect 11011 31464 11023 31467
rect 11698 31464 11704 31476
rect 11011 31436 11704 31464
rect 11011 31433 11023 31436
rect 10965 31427 11023 31433
rect 11698 31424 11704 31436
rect 11756 31424 11762 31476
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 16482 31464 16488 31476
rect 13872 31436 16488 31464
rect 13872 31424 13878 31436
rect 16482 31424 16488 31436
rect 16540 31424 16546 31476
rect 16853 31467 16911 31473
rect 16853 31433 16865 31467
rect 16899 31464 16911 31467
rect 17402 31464 17408 31476
rect 16899 31436 17408 31464
rect 16899 31433 16911 31436
rect 16853 31427 16911 31433
rect 17402 31424 17408 31436
rect 17460 31424 17466 31476
rect 19058 31424 19064 31476
rect 19116 31464 19122 31476
rect 19116 31436 21404 31464
rect 19116 31424 19122 31436
rect 14734 31396 14740 31408
rect 11164 31368 14740 31396
rect 11164 31337 11192 31368
rect 14734 31356 14740 31368
rect 14792 31356 14798 31408
rect 15188 31399 15246 31405
rect 15188 31365 15200 31399
rect 15234 31396 15246 31399
rect 15234 31368 21312 31396
rect 15234 31365 15246 31368
rect 15188 31359 15246 31365
rect 11149 31331 11207 31337
rect 11149 31297 11161 31331
rect 11195 31297 11207 31331
rect 11149 31291 11207 31297
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 13354 31337 13360 31340
rect 12621 31331 12679 31337
rect 12621 31328 12633 31331
rect 12492 31300 12633 31328
rect 12492 31288 12498 31300
rect 12621 31297 12633 31300
rect 12667 31297 12679 31331
rect 12621 31291 12679 31297
rect 13348 31291 13360 31337
rect 13354 31288 13360 31291
rect 13412 31288 13418 31340
rect 15470 31288 15476 31340
rect 15528 31328 15534 31340
rect 15528 31300 15976 31328
rect 15528 31288 15534 31300
rect 12253 31263 12311 31269
rect 12253 31260 12265 31263
rect 10244 31232 12265 31260
rect 12253 31229 12265 31232
rect 12299 31229 12311 31263
rect 12253 31223 12311 31229
rect 13078 31220 13084 31272
rect 13136 31220 13142 31272
rect 14550 31220 14556 31272
rect 14608 31260 14614 31272
rect 14921 31263 14979 31269
rect 14921 31260 14933 31263
rect 14608 31232 14933 31260
rect 14608 31220 14614 31232
rect 14921 31229 14933 31232
rect 14967 31229 14979 31263
rect 15948 31260 15976 31300
rect 16574 31288 16580 31340
rect 16632 31328 16638 31340
rect 17037 31331 17095 31337
rect 17037 31328 17049 31331
rect 16632 31300 17049 31328
rect 16632 31288 16638 31300
rect 17037 31297 17049 31300
rect 17083 31297 17095 31331
rect 17753 31331 17811 31337
rect 17753 31328 17765 31331
rect 17037 31291 17095 31297
rect 17144 31300 17765 31328
rect 17144 31260 17172 31300
rect 17753 31297 17765 31300
rect 17799 31297 17811 31331
rect 19593 31331 19651 31337
rect 19593 31328 19605 31331
rect 17753 31291 17811 31297
rect 18524 31300 19605 31328
rect 15948 31232 17172 31260
rect 14921 31223 14979 31229
rect 17494 31220 17500 31272
rect 17552 31220 17558 31272
rect 2041 31195 2099 31201
rect 2041 31161 2053 31195
rect 2087 31192 2099 31195
rect 3234 31192 3240 31204
rect 2087 31164 3240 31192
rect 2087 31161 2099 31164
rect 2041 31155 2099 31161
rect 3234 31152 3240 31164
rect 3292 31152 3298 31204
rect 7834 31152 7840 31204
rect 7892 31192 7898 31204
rect 8665 31195 8723 31201
rect 8665 31192 8677 31195
rect 7892 31164 8677 31192
rect 7892 31152 7898 31164
rect 8665 31161 8677 31164
rect 8711 31161 8723 31195
rect 8665 31155 8723 31161
rect 16666 31152 16672 31204
rect 16724 31192 16730 31204
rect 17512 31192 17540 31220
rect 16724 31164 17540 31192
rect 16724 31152 16730 31164
rect 1578 31084 1584 31136
rect 1636 31124 1642 31136
rect 2498 31124 2504 31136
rect 1636 31096 2504 31124
rect 1636 31084 1642 31096
rect 2498 31084 2504 31096
rect 2556 31124 2562 31136
rect 3789 31127 3847 31133
rect 3789 31124 3801 31127
rect 2556 31096 3801 31124
rect 2556 31084 2562 31096
rect 3789 31093 3801 31096
rect 3835 31093 3847 31127
rect 3789 31087 3847 31093
rect 4338 31084 4344 31136
rect 4396 31124 4402 31136
rect 10226 31124 10232 31136
rect 4396 31096 10232 31124
rect 4396 31084 4402 31096
rect 10226 31084 10232 31096
rect 10284 31084 10290 31136
rect 10410 31084 10416 31136
rect 10468 31124 10474 31136
rect 10505 31127 10563 31133
rect 10505 31124 10517 31127
rect 10468 31096 10517 31124
rect 10468 31084 10474 31096
rect 10505 31093 10517 31096
rect 10551 31124 10563 31127
rect 10594 31124 10600 31136
rect 10551 31096 10600 31124
rect 10551 31093 10563 31096
rect 10505 31087 10563 31093
rect 10594 31084 10600 31096
rect 10652 31084 10658 31136
rect 12621 31127 12679 31133
rect 12621 31093 12633 31127
rect 12667 31124 12679 31127
rect 13722 31124 13728 31136
rect 12667 31096 13728 31124
rect 12667 31093 12679 31096
rect 12621 31087 12679 31093
rect 13722 31084 13728 31096
rect 13780 31084 13786 31136
rect 14458 31084 14464 31136
rect 14516 31084 14522 31136
rect 15194 31084 15200 31136
rect 15252 31124 15258 31136
rect 16301 31127 16359 31133
rect 16301 31124 16313 31127
rect 15252 31096 16313 31124
rect 15252 31084 15258 31096
rect 16301 31093 16313 31096
rect 16347 31093 16359 31127
rect 16301 31087 16359 31093
rect 17218 31084 17224 31136
rect 17276 31124 17282 31136
rect 18524 31124 18552 31300
rect 19593 31297 19605 31300
rect 19639 31297 19651 31331
rect 19593 31291 19651 31297
rect 19334 31220 19340 31272
rect 19392 31220 19398 31272
rect 21284 31260 21312 31368
rect 21376 31337 21404 31436
rect 21726 31424 21732 31476
rect 21784 31464 21790 31476
rect 24489 31467 24547 31473
rect 24489 31464 24501 31467
rect 21784 31436 24501 31464
rect 21784 31424 21790 31436
rect 24489 31433 24501 31436
rect 24535 31433 24547 31467
rect 24489 31427 24547 31433
rect 27157 31467 27215 31473
rect 27157 31433 27169 31467
rect 27203 31433 27215 31467
rect 27157 31427 27215 31433
rect 27172 31396 27200 31427
rect 21468 31368 27200 31396
rect 21361 31331 21419 31337
rect 21361 31297 21373 31331
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 21468 31260 21496 31368
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 22261 31331 22319 31337
rect 22261 31328 22273 31331
rect 21692 31300 22273 31328
rect 21692 31288 21698 31300
rect 22261 31297 22273 31300
rect 22307 31297 22319 31331
rect 22261 31291 22319 31297
rect 23658 31288 23664 31340
rect 23716 31328 23722 31340
rect 23845 31331 23903 31337
rect 23845 31328 23857 31331
rect 23716 31300 23857 31328
rect 23716 31288 23722 31300
rect 23845 31297 23857 31300
rect 23891 31297 23903 31331
rect 23845 31291 23903 31297
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 21284 31232 21496 31260
rect 21542 31220 21548 31272
rect 21600 31260 21606 31272
rect 22005 31263 22063 31269
rect 22005 31260 22017 31263
rect 21600 31232 22017 31260
rect 21600 31220 21606 31232
rect 22005 31229 22017 31232
rect 22051 31229 22063 31263
rect 24044 31260 24072 31291
rect 24670 31288 24676 31340
rect 24728 31288 24734 31340
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 25317 31331 25375 31337
rect 25317 31328 25329 31331
rect 25004 31300 25329 31328
rect 25004 31288 25010 31300
rect 25317 31297 25329 31300
rect 25363 31297 25375 31331
rect 25317 31291 25375 31297
rect 25958 31288 25964 31340
rect 26016 31328 26022 31340
rect 26421 31331 26479 31337
rect 26421 31328 26433 31331
rect 26016 31300 26433 31328
rect 26016 31288 26022 31300
rect 26421 31297 26433 31300
rect 26467 31297 26479 31331
rect 26421 31291 26479 31297
rect 26605 31331 26663 31337
rect 26605 31297 26617 31331
rect 26651 31297 26663 31331
rect 26605 31291 26663 31297
rect 26234 31260 26240 31272
rect 24044 31232 26240 31260
rect 22005 31223 22063 31229
rect 26234 31220 26240 31232
rect 26292 31220 26298 31272
rect 26620 31260 26648 31291
rect 26786 31288 26792 31340
rect 26844 31328 26850 31340
rect 27341 31331 27399 31337
rect 27341 31328 27353 31331
rect 26844 31300 27353 31328
rect 26844 31288 26850 31300
rect 27341 31297 27353 31300
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27985 31263 28043 31269
rect 27985 31260 27997 31263
rect 26620 31232 27997 31260
rect 27985 31229 27997 31232
rect 28031 31229 28043 31263
rect 27985 31223 28043 31229
rect 20714 31152 20720 31204
rect 20772 31152 20778 31204
rect 20990 31152 20996 31204
rect 21048 31192 21054 31204
rect 21048 31164 21588 31192
rect 21048 31152 21054 31164
rect 17276 31096 18552 31124
rect 17276 31084 17282 31096
rect 18690 31084 18696 31136
rect 18748 31124 18754 31136
rect 18877 31127 18935 31133
rect 18877 31124 18889 31127
rect 18748 31096 18889 31124
rect 18748 31084 18754 31096
rect 18877 31093 18889 31096
rect 18923 31093 18935 31127
rect 18877 31087 18935 31093
rect 21177 31127 21235 31133
rect 21177 31093 21189 31127
rect 21223 31124 21235 31127
rect 21450 31124 21456 31136
rect 21223 31096 21456 31124
rect 21223 31093 21235 31096
rect 21177 31087 21235 31093
rect 21450 31084 21456 31096
rect 21508 31084 21514 31136
rect 21560 31124 21588 31164
rect 25774 31152 25780 31204
rect 25832 31192 25838 31204
rect 25961 31195 26019 31201
rect 25961 31192 25973 31195
rect 25832 31164 25973 31192
rect 25832 31152 25838 31164
rect 25961 31161 25973 31164
rect 26007 31161 26019 31195
rect 25961 31155 26019 31161
rect 23385 31127 23443 31133
rect 23385 31124 23397 31127
rect 21560 31096 23397 31124
rect 23385 31093 23397 31096
rect 23431 31093 23443 31127
rect 23385 31087 23443 31093
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 26786 31124 26792 31136
rect 26568 31096 26792 31124
rect 26568 31084 26574 31096
rect 26786 31084 26792 31096
rect 26844 31084 26850 31136
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 9950 30880 9956 30932
rect 10008 30880 10014 30932
rect 13722 30880 13728 30932
rect 13780 30880 13786 30932
rect 13814 30880 13820 30932
rect 13872 30920 13878 30932
rect 15657 30923 15715 30929
rect 15657 30920 15669 30923
rect 13872 30892 15669 30920
rect 13872 30880 13878 30892
rect 15657 30889 15669 30892
rect 15703 30889 15715 30923
rect 18230 30920 18236 30932
rect 15657 30883 15715 30889
rect 17328 30892 18236 30920
rect 3878 30812 3884 30864
rect 3936 30852 3942 30864
rect 4065 30855 4123 30861
rect 4065 30852 4077 30855
rect 3936 30824 4077 30852
rect 3936 30812 3942 30824
rect 4065 30821 4077 30824
rect 4111 30821 4123 30855
rect 4065 30815 4123 30821
rect 6086 30812 6092 30864
rect 6144 30852 6150 30864
rect 6917 30855 6975 30861
rect 6917 30852 6929 30855
rect 6144 30824 6929 30852
rect 6144 30812 6150 30824
rect 6917 30821 6929 30824
rect 6963 30852 6975 30855
rect 6963 30824 7880 30852
rect 6963 30821 6975 30824
rect 6917 30815 6975 30821
rect 3326 30744 3332 30796
rect 3384 30744 3390 30796
rect 7852 30793 7880 30824
rect 13078 30812 13084 30864
rect 13136 30852 13142 30864
rect 13136 30824 14320 30852
rect 13136 30812 13142 30824
rect 7837 30787 7895 30793
rect 7837 30753 7849 30787
rect 7883 30753 7895 30787
rect 7837 30747 7895 30753
rect 9030 30744 9036 30796
rect 9088 30784 9094 30796
rect 9585 30787 9643 30793
rect 9585 30784 9597 30787
rect 9088 30756 9597 30784
rect 9088 30744 9094 30756
rect 9585 30753 9597 30756
rect 9631 30753 9643 30787
rect 9585 30747 9643 30753
rect 12161 30787 12219 30793
rect 12161 30753 12173 30787
rect 12207 30784 12219 30787
rect 13630 30784 13636 30796
rect 12207 30756 13636 30784
rect 12207 30753 12219 30756
rect 12161 30747 12219 30753
rect 13630 30744 13636 30756
rect 13688 30744 13694 30796
rect 13722 30744 13728 30796
rect 13780 30744 13786 30796
rect 14292 30793 14320 30824
rect 16482 30812 16488 30864
rect 16540 30852 16546 30864
rect 17328 30861 17356 30892
rect 18230 30880 18236 30892
rect 18288 30880 18294 30932
rect 18417 30923 18475 30929
rect 18417 30889 18429 30923
rect 18463 30920 18475 30923
rect 18782 30920 18788 30932
rect 18463 30892 18788 30920
rect 18463 30889 18475 30892
rect 18417 30883 18475 30889
rect 18782 30880 18788 30892
rect 18840 30880 18846 30932
rect 18874 30880 18880 30932
rect 18932 30920 18938 30932
rect 20901 30923 20959 30929
rect 20901 30920 20913 30923
rect 18932 30892 20913 30920
rect 18932 30880 18938 30892
rect 20901 30889 20913 30892
rect 20947 30889 20959 30923
rect 21542 30920 21548 30932
rect 20901 30883 20959 30889
rect 21376 30892 21548 30920
rect 17313 30855 17371 30861
rect 17313 30852 17325 30855
rect 16540 30824 17325 30852
rect 16540 30812 16546 30824
rect 17313 30821 17325 30824
rect 17359 30821 17371 30855
rect 17313 30815 17371 30821
rect 17773 30855 17831 30861
rect 17773 30821 17785 30855
rect 17819 30852 17831 30855
rect 19518 30852 19524 30864
rect 17819 30824 19524 30852
rect 17819 30821 17831 30824
rect 17773 30815 17831 30821
rect 19518 30812 19524 30824
rect 19576 30812 19582 30864
rect 14277 30787 14335 30793
rect 14277 30753 14289 30787
rect 14323 30753 14335 30787
rect 14277 30747 14335 30753
rect 15378 30744 15384 30796
rect 15436 30784 15442 30796
rect 16117 30787 16175 30793
rect 16117 30784 16129 30787
rect 15436 30756 16129 30784
rect 15436 30744 15442 30756
rect 16117 30753 16129 30756
rect 16163 30753 16175 30787
rect 17678 30784 17684 30796
rect 16117 30747 16175 30753
rect 17236 30756 17684 30784
rect 1578 30676 1584 30728
rect 1636 30676 1642 30728
rect 2406 30676 2412 30728
rect 2464 30716 2470 30728
rect 4617 30719 4675 30725
rect 4617 30716 4629 30719
rect 2464 30688 4629 30716
rect 2464 30676 2470 30688
rect 4617 30685 4629 30688
rect 4663 30685 4675 30719
rect 4617 30679 4675 30685
rect 4338 30608 4344 30660
rect 4396 30608 4402 30660
rect 4632 30648 4660 30679
rect 5718 30676 5724 30728
rect 5776 30716 5782 30728
rect 6546 30716 6552 30728
rect 5776 30688 6552 30716
rect 5776 30676 5782 30688
rect 6546 30676 6552 30688
rect 6604 30716 6610 30728
rect 6822 30716 6828 30728
rect 6604 30688 6828 30716
rect 6604 30676 6610 30688
rect 6822 30676 6828 30688
rect 6880 30676 6886 30728
rect 7561 30719 7619 30725
rect 7561 30685 7573 30719
rect 7607 30716 7619 30719
rect 8294 30716 8300 30728
rect 7607 30688 8300 30716
rect 7607 30685 7619 30688
rect 7561 30679 7619 30685
rect 8294 30676 8300 30688
rect 8352 30676 8358 30728
rect 9674 30676 9680 30728
rect 9732 30716 9738 30728
rect 9953 30719 10011 30725
rect 9953 30716 9965 30719
rect 9732 30688 9965 30716
rect 9732 30676 9738 30688
rect 9953 30685 9965 30688
rect 9999 30716 10011 30719
rect 10134 30716 10140 30728
rect 9999 30688 10140 30716
rect 9999 30685 10011 30688
rect 9953 30679 10011 30685
rect 10134 30676 10140 30688
rect 10192 30676 10198 30728
rect 10594 30676 10600 30728
rect 10652 30716 10658 30728
rect 12621 30719 12679 30725
rect 12621 30716 12633 30719
rect 10652 30688 12633 30716
rect 10652 30676 10658 30688
rect 12621 30685 12633 30688
rect 12667 30685 12679 30719
rect 13357 30719 13415 30725
rect 13357 30716 13369 30719
rect 12621 30679 12679 30685
rect 12820 30688 13369 30716
rect 6730 30648 6736 30660
rect 4632 30620 6736 30648
rect 6730 30608 6736 30620
rect 6788 30608 6794 30660
rect 10413 30651 10471 30657
rect 10413 30617 10425 30651
rect 10459 30648 10471 30651
rect 12710 30648 12716 30660
rect 10459 30620 12716 30648
rect 10459 30617 10471 30620
rect 10413 30611 10471 30617
rect 12710 30608 12716 30620
rect 12768 30608 12774 30660
rect 4246 30540 4252 30592
rect 4304 30580 4310 30592
rect 4525 30583 4583 30589
rect 4525 30580 4537 30583
rect 4304 30552 4537 30580
rect 4304 30540 4310 30552
rect 4525 30549 4537 30552
rect 4571 30549 4583 30583
rect 4525 30543 4583 30549
rect 5166 30540 5172 30592
rect 5224 30580 5230 30592
rect 6089 30583 6147 30589
rect 6089 30580 6101 30583
rect 5224 30552 6101 30580
rect 5224 30540 5230 30552
rect 6089 30549 6101 30552
rect 6135 30580 6147 30583
rect 6917 30583 6975 30589
rect 6917 30580 6929 30583
rect 6135 30552 6929 30580
rect 6135 30549 6147 30552
rect 6089 30543 6147 30549
rect 6917 30549 6929 30552
rect 6963 30549 6975 30583
rect 6917 30543 6975 30549
rect 7466 30540 7472 30592
rect 7524 30580 7530 30592
rect 11698 30580 11704 30592
rect 7524 30552 11704 30580
rect 7524 30540 7530 30552
rect 11698 30540 11704 30552
rect 11756 30580 11762 30592
rect 12820 30589 12848 30688
rect 13357 30685 13369 30688
rect 13403 30685 13415 30719
rect 15562 30716 15568 30728
rect 13357 30679 13415 30685
rect 14476 30688 15568 30716
rect 12894 30608 12900 30660
rect 12952 30648 12958 30660
rect 14476 30648 14504 30688
rect 15562 30676 15568 30688
rect 15620 30676 15626 30728
rect 16132 30716 16160 30747
rect 16945 30719 17003 30725
rect 16132 30712 16896 30716
rect 16945 30712 16957 30719
rect 16132 30688 16957 30712
rect 16868 30685 16957 30688
rect 16991 30712 17003 30719
rect 17236 30716 17264 30756
rect 17678 30744 17684 30756
rect 17736 30744 17742 30796
rect 18046 30744 18052 30796
rect 18104 30784 18110 30796
rect 21376 30793 21404 30892
rect 21542 30880 21548 30892
rect 21600 30880 21606 30932
rect 22278 30880 22284 30932
rect 22336 30920 22342 30932
rect 23934 30920 23940 30932
rect 22336 30892 23940 30920
rect 22336 30880 22342 30892
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 25130 30880 25136 30932
rect 25188 30920 25194 30932
rect 25409 30923 25467 30929
rect 25409 30920 25421 30923
rect 25188 30892 25421 30920
rect 25188 30880 25194 30892
rect 25409 30889 25421 30892
rect 25455 30889 25467 30923
rect 25409 30883 25467 30889
rect 26234 30880 26240 30932
rect 26292 30920 26298 30932
rect 26697 30923 26755 30929
rect 26697 30920 26709 30923
rect 26292 30892 26709 30920
rect 26292 30880 26298 30892
rect 26697 30889 26709 30892
rect 26743 30889 26755 30923
rect 26697 30883 26755 30889
rect 27798 30812 27804 30864
rect 27856 30812 27862 30864
rect 21361 30787 21419 30793
rect 18104 30756 19656 30784
rect 18104 30744 18110 30756
rect 17770 30716 17776 30728
rect 17052 30712 17264 30716
rect 16991 30688 17264 30712
rect 17328 30688 17776 30716
rect 16991 30685 17080 30688
rect 16868 30684 17080 30685
rect 17135 30684 17172 30688
rect 16945 30679 17003 30684
rect 12952 30620 14504 30648
rect 14544 30651 14602 30657
rect 12952 30608 12958 30620
rect 14544 30617 14556 30651
rect 14590 30648 14602 30651
rect 15930 30648 15936 30660
rect 14590 30620 15936 30648
rect 14590 30617 14602 30620
rect 14544 30611 14602 30617
rect 15930 30608 15936 30620
rect 15988 30608 15994 30660
rect 12805 30583 12863 30589
rect 12805 30580 12817 30583
rect 11756 30552 12817 30580
rect 11756 30540 11762 30552
rect 12805 30549 12817 30552
rect 12851 30549 12863 30583
rect 12805 30543 12863 30549
rect 14642 30540 14648 30592
rect 14700 30580 14706 30592
rect 15286 30580 15292 30592
rect 14700 30552 15292 30580
rect 14700 30540 14706 30552
rect 15286 30540 15292 30552
rect 15344 30540 15350 30592
rect 15470 30540 15476 30592
rect 15528 30580 15534 30592
rect 15654 30580 15660 30592
rect 15528 30552 15660 30580
rect 15528 30540 15534 30552
rect 15654 30540 15660 30552
rect 15712 30580 15718 30592
rect 17328 30589 17356 30688
rect 17770 30676 17776 30688
rect 17828 30676 17834 30728
rect 17954 30676 17960 30728
rect 18012 30676 18018 30728
rect 18601 30719 18659 30725
rect 18601 30685 18613 30719
rect 18647 30685 18659 30719
rect 18601 30679 18659 30685
rect 17862 30608 17868 30660
rect 17920 30648 17926 30660
rect 18616 30648 18644 30679
rect 19426 30676 19432 30728
rect 19484 30716 19490 30728
rect 19521 30719 19579 30725
rect 19521 30716 19533 30719
rect 19484 30688 19533 30716
rect 19484 30676 19490 30688
rect 19521 30685 19533 30688
rect 19567 30685 19579 30719
rect 19628 30716 19656 30756
rect 21361 30753 21373 30787
rect 21407 30753 21419 30787
rect 21361 30747 21419 30753
rect 24029 30787 24087 30793
rect 24029 30753 24041 30787
rect 24075 30784 24087 30787
rect 24075 30756 24808 30784
rect 24075 30753 24087 30756
rect 24029 30747 24087 30753
rect 19628 30688 21404 30716
rect 19521 30679 19579 30685
rect 17920 30620 18644 30648
rect 19788 30651 19846 30657
rect 17920 30608 17926 30620
rect 19788 30617 19800 30651
rect 19834 30648 19846 30651
rect 20714 30648 20720 30660
rect 19834 30620 20720 30648
rect 19834 30617 19846 30620
rect 19788 30611 19846 30617
rect 20714 30608 20720 30620
rect 20772 30608 20778 30660
rect 21376 30648 21404 30688
rect 21450 30676 21456 30728
rect 21508 30716 21514 30728
rect 21617 30719 21675 30725
rect 21617 30716 21629 30719
rect 21508 30688 21629 30716
rect 21508 30676 21514 30688
rect 21617 30685 21629 30688
rect 21663 30685 21675 30719
rect 21617 30679 21675 30685
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 23566 30716 23572 30728
rect 23431 30688 23572 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 24578 30676 24584 30728
rect 24636 30676 24642 30728
rect 24780 30725 24808 30756
rect 25958 30744 25964 30796
rect 26016 30784 26022 30796
rect 26016 30756 26188 30784
rect 26016 30744 26022 30756
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 26053 30719 26111 30725
rect 26053 30716 26065 30719
rect 25004 30688 26065 30716
rect 25004 30676 25010 30688
rect 26053 30685 26065 30688
rect 26099 30685 26111 30719
rect 26160 30716 26188 30756
rect 27062 30744 27068 30796
rect 27120 30784 27126 30796
rect 27295 30787 27353 30793
rect 27295 30784 27307 30787
rect 27120 30756 27307 30784
rect 27120 30744 27126 30756
rect 27295 30753 27307 30756
rect 27341 30753 27353 30787
rect 27295 30747 27353 30753
rect 27192 30719 27250 30725
rect 27192 30716 27204 30719
rect 26160 30688 27204 30716
rect 26053 30679 26111 30685
rect 27192 30685 27204 30688
rect 27238 30685 27250 30719
rect 27192 30679 27250 30685
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 21726 30648 21732 30660
rect 20824 30620 21036 30648
rect 21376 30620 21732 30648
rect 16485 30583 16543 30589
rect 16485 30580 16497 30583
rect 15712 30552 16497 30580
rect 15712 30540 15718 30552
rect 16485 30549 16497 30552
rect 16531 30580 16543 30583
rect 17313 30583 17371 30589
rect 17313 30580 17325 30583
rect 16531 30552 17325 30580
rect 16531 30549 16543 30552
rect 16485 30543 16543 30549
rect 17313 30549 17325 30552
rect 17359 30549 17371 30583
rect 17313 30543 17371 30549
rect 17402 30540 17408 30592
rect 17460 30580 17466 30592
rect 20824 30580 20852 30620
rect 17460 30552 20852 30580
rect 21008 30580 21036 30620
rect 21726 30608 21732 30620
rect 21784 30608 21790 30660
rect 28000 30648 28028 30679
rect 22066 30620 28028 30648
rect 22066 30580 22094 30620
rect 21008 30552 22094 30580
rect 17460 30540 17466 30552
rect 22370 30540 22376 30592
rect 22428 30580 22434 30592
rect 22741 30583 22799 30589
rect 22741 30580 22753 30583
rect 22428 30552 22753 30580
rect 22428 30540 22434 30552
rect 22741 30549 22753 30552
rect 22787 30549 22799 30583
rect 22741 30543 22799 30549
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 3970 30336 3976 30388
rect 4028 30376 4034 30388
rect 5261 30379 5319 30385
rect 5261 30376 5273 30379
rect 4028 30348 5273 30376
rect 4028 30336 4034 30348
rect 5261 30345 5273 30348
rect 5307 30376 5319 30379
rect 5534 30376 5540 30388
rect 5307 30348 5540 30376
rect 5307 30345 5319 30348
rect 5261 30339 5319 30345
rect 5534 30336 5540 30348
rect 5592 30336 5598 30388
rect 7558 30336 7564 30388
rect 7616 30336 7622 30388
rect 9950 30336 9956 30388
rect 10008 30376 10014 30388
rect 12066 30376 12072 30388
rect 10008 30348 12072 30376
rect 10008 30336 10014 30348
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 12158 30336 12164 30388
rect 12216 30376 12222 30388
rect 12216 30348 13400 30376
rect 12216 30336 12222 30348
rect 2130 30268 2136 30320
rect 2188 30268 2194 30320
rect 7006 30268 7012 30320
rect 7064 30308 7070 30320
rect 7193 30311 7251 30317
rect 7193 30308 7205 30311
rect 7064 30280 7205 30308
rect 7064 30268 7070 30280
rect 7193 30277 7205 30280
rect 7239 30308 7251 30311
rect 7576 30308 7604 30336
rect 7239 30280 7604 30308
rect 7239 30277 7251 30280
rect 7193 30271 7251 30277
rect 7650 30268 7656 30320
rect 7708 30308 7714 30320
rect 10036 30311 10094 30317
rect 7708 30280 8156 30308
rect 7708 30268 7714 30280
rect 1946 30200 1952 30252
rect 2004 30200 2010 30252
rect 2038 30200 2044 30252
rect 2096 30200 2102 30252
rect 2225 30243 2283 30249
rect 2225 30209 2237 30243
rect 2271 30209 2283 30243
rect 2225 30203 2283 30209
rect 1765 30039 1823 30045
rect 1765 30005 1777 30039
rect 1811 30036 1823 30039
rect 1854 30036 1860 30048
rect 1811 30008 1860 30036
rect 1811 30005 1823 30008
rect 1765 29999 1823 30005
rect 1854 29996 1860 30008
rect 1912 29996 1918 30048
rect 2240 30036 2268 30203
rect 2314 30200 2320 30252
rect 2372 30240 2378 30252
rect 2409 30243 2467 30249
rect 2409 30240 2421 30243
rect 2372 30212 2421 30240
rect 2372 30200 2378 30212
rect 2409 30209 2421 30212
rect 2455 30209 2467 30243
rect 2409 30203 2467 30209
rect 2866 30200 2872 30252
rect 2924 30200 2930 30252
rect 4890 30200 4896 30252
rect 4948 30240 4954 30252
rect 5261 30243 5319 30249
rect 5261 30240 5273 30243
rect 4948 30212 5273 30240
rect 4948 30200 4954 30212
rect 5261 30209 5273 30212
rect 5307 30209 5319 30243
rect 5261 30203 5319 30209
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30209 6791 30243
rect 6733 30203 6791 30209
rect 4617 30175 4675 30181
rect 4617 30141 4629 30175
rect 4663 30172 4675 30175
rect 4798 30172 4804 30184
rect 4663 30144 4804 30172
rect 4663 30141 4675 30144
rect 4617 30135 4675 30141
rect 4798 30132 4804 30144
rect 4856 30132 4862 30184
rect 5077 30175 5135 30181
rect 5077 30141 5089 30175
rect 5123 30141 5135 30175
rect 5077 30135 5135 30141
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30172 5687 30175
rect 5994 30172 6000 30184
rect 5675 30144 6000 30172
rect 5675 30141 5687 30144
rect 5629 30135 5687 30141
rect 5092 30104 5120 30135
rect 5994 30132 6000 30144
rect 6052 30132 6058 30184
rect 6748 30172 6776 30203
rect 6822 30200 6828 30252
rect 6880 30240 6886 30252
rect 8128 30249 8156 30280
rect 10036 30277 10048 30311
rect 10082 30308 10094 30311
rect 10134 30308 10140 30320
rect 10082 30280 10140 30308
rect 10082 30277 10094 30280
rect 10036 30271 10094 30277
rect 10134 30268 10140 30280
rect 10192 30268 10198 30320
rect 10686 30268 10692 30320
rect 10744 30268 10750 30320
rect 13078 30308 13084 30320
rect 10980 30280 12204 30308
rect 8113 30243 8171 30249
rect 6880 30212 7788 30240
rect 6880 30200 6886 30212
rect 7098 30172 7104 30184
rect 6748 30144 7104 30172
rect 7098 30132 7104 30144
rect 7156 30132 7162 30184
rect 7650 30132 7656 30184
rect 7708 30132 7714 30184
rect 7760 30172 7788 30212
rect 8113 30209 8125 30243
rect 8159 30209 8171 30243
rect 10704 30240 10732 30268
rect 10980 30240 11008 30280
rect 8113 30203 8171 30209
rect 9784 30212 11008 30240
rect 9784 30184 9812 30212
rect 12066 30200 12072 30252
rect 12124 30200 12130 30252
rect 12176 30240 12204 30280
rect 12728 30280 13084 30308
rect 12728 30249 12756 30280
rect 13078 30268 13084 30280
rect 13136 30268 13142 30320
rect 13372 30308 13400 30348
rect 13446 30336 13452 30388
rect 13504 30376 13510 30388
rect 14182 30376 14188 30388
rect 13504 30348 14188 30376
rect 13504 30336 13510 30348
rect 14182 30336 14188 30348
rect 14240 30336 14246 30388
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 14826 30376 14832 30388
rect 14516 30348 14832 30376
rect 14516 30336 14522 30348
rect 14826 30336 14832 30348
rect 14884 30336 14890 30388
rect 15746 30336 15752 30388
rect 15804 30376 15810 30388
rect 15841 30379 15899 30385
rect 15841 30376 15853 30379
rect 15804 30348 15853 30376
rect 15804 30336 15810 30348
rect 15841 30345 15853 30348
rect 15887 30345 15899 30379
rect 15841 30339 15899 30345
rect 17052 30348 17264 30376
rect 15378 30308 15384 30320
rect 13372 30280 15384 30308
rect 15378 30268 15384 30280
rect 15436 30268 15442 30320
rect 15930 30268 15936 30320
rect 15988 30308 15994 30320
rect 17052 30308 17080 30348
rect 17126 30317 17132 30320
rect 15988 30280 17080 30308
rect 15988 30268 15994 30280
rect 17120 30271 17132 30317
rect 17126 30268 17132 30271
rect 17184 30268 17190 30320
rect 17236 30308 17264 30348
rect 17678 30336 17684 30388
rect 17736 30376 17742 30388
rect 18690 30376 18696 30388
rect 17736 30348 18696 30376
rect 17736 30336 17742 30348
rect 18690 30336 18696 30348
rect 18748 30336 18754 30388
rect 20714 30336 20720 30388
rect 20772 30336 20778 30388
rect 22186 30376 22192 30388
rect 22020 30348 22192 30376
rect 18138 30308 18144 30320
rect 17236 30280 18144 30308
rect 18138 30268 18144 30280
rect 18196 30268 18202 30320
rect 12713 30243 12771 30249
rect 12713 30240 12725 30243
rect 12176 30212 12725 30240
rect 12713 30209 12725 30212
rect 12759 30209 12771 30243
rect 12713 30203 12771 30209
rect 12980 30243 13038 30249
rect 12980 30209 12992 30243
rect 13026 30240 13038 30243
rect 13722 30240 13728 30252
rect 13026 30212 13728 30240
rect 13026 30209 13038 30212
rect 12980 30203 13038 30209
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 15286 30200 15292 30252
rect 15344 30240 15350 30252
rect 20257 30243 20315 30249
rect 20257 30240 20269 30243
rect 15344 30212 20269 30240
rect 15344 30200 15350 30212
rect 20257 30209 20269 30212
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 20898 30200 20904 30252
rect 20956 30200 20962 30252
rect 22020 30249 22048 30348
rect 22186 30336 22192 30348
rect 22244 30376 22250 30388
rect 23198 30376 23204 30388
rect 22244 30348 23204 30376
rect 22244 30336 22250 30348
rect 23198 30336 23204 30348
rect 23256 30336 23262 30388
rect 23474 30308 23480 30320
rect 22204 30280 23480 30308
rect 22204 30249 22232 30280
rect 23474 30268 23480 30280
rect 23532 30268 23538 30320
rect 25332 30280 25636 30308
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 23089 30243 23147 30249
rect 23089 30240 23101 30243
rect 22189 30203 22247 30209
rect 22388 30212 23101 30240
rect 8389 30175 8447 30181
rect 8389 30172 8401 30175
rect 7760 30144 8401 30172
rect 8389 30141 8401 30144
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 9766 30132 9772 30184
rect 9824 30132 9830 30184
rect 11698 30132 11704 30184
rect 11756 30132 11762 30184
rect 14458 30132 14464 30184
rect 14516 30172 14522 30184
rect 14553 30175 14611 30181
rect 14553 30172 14565 30175
rect 14516 30144 14565 30172
rect 14516 30132 14522 30144
rect 14553 30141 14565 30144
rect 14599 30141 14611 30175
rect 14553 30135 14611 30141
rect 14734 30132 14740 30184
rect 14792 30172 14798 30184
rect 15013 30175 15071 30181
rect 15013 30172 15025 30175
rect 14792 30144 15025 30172
rect 14792 30132 14798 30144
rect 15013 30141 15025 30144
rect 15059 30141 15071 30175
rect 15013 30135 15071 30141
rect 15470 30132 15476 30184
rect 15528 30132 15534 30184
rect 16853 30175 16911 30181
rect 16853 30141 16865 30175
rect 16899 30141 16911 30175
rect 16853 30135 16911 30141
rect 5810 30104 5816 30116
rect 5092 30076 5816 30104
rect 5810 30064 5816 30076
rect 5868 30064 5874 30116
rect 7374 30104 7380 30116
rect 6472 30076 7380 30104
rect 6472 30036 6500 30076
rect 7374 30064 7380 30076
rect 7432 30064 7438 30116
rect 7561 30107 7619 30113
rect 7561 30073 7573 30107
rect 7607 30104 7619 30107
rect 11974 30104 11980 30116
rect 7607 30076 9812 30104
rect 7607 30073 7619 30076
rect 7561 30067 7619 30073
rect 2240 30008 6500 30036
rect 6549 30039 6607 30045
rect 6549 30005 6561 30039
rect 6595 30036 6607 30039
rect 9582 30036 9588 30048
rect 6595 30008 9588 30036
rect 6595 30005 6607 30008
rect 6549 29999 6607 30005
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 9784 30036 9812 30076
rect 10704 30076 11980 30104
rect 10704 30048 10732 30076
rect 11974 30064 11980 30076
rect 12032 30064 12038 30116
rect 14921 30107 14979 30113
rect 14921 30073 14933 30107
rect 14967 30073 14979 30107
rect 14921 30067 14979 30073
rect 10686 30036 10692 30048
rect 9784 30008 10692 30036
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 11146 29996 11152 30048
rect 11204 30036 11210 30048
rect 11790 30036 11796 30048
rect 11204 30008 11796 30036
rect 11204 29996 11210 30008
rect 11790 29996 11796 30008
rect 11848 29996 11854 30048
rect 12526 29996 12532 30048
rect 12584 30036 12590 30048
rect 14093 30039 14151 30045
rect 14093 30036 14105 30039
rect 12584 30008 14105 30036
rect 12584 29996 12590 30008
rect 14093 30005 14105 30008
rect 14139 30005 14151 30039
rect 14936 30036 14964 30067
rect 15838 30064 15844 30116
rect 15896 30064 15902 30116
rect 15562 30036 15568 30048
rect 14936 30008 15568 30036
rect 14093 29999 14151 30005
rect 15562 29996 15568 30008
rect 15620 30036 15626 30048
rect 15930 30036 15936 30048
rect 15620 30008 15936 30036
rect 15620 29996 15626 30008
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 16114 29996 16120 30048
rect 16172 30036 16178 30048
rect 16868 30036 16896 30135
rect 18230 30132 18236 30184
rect 18288 30172 18294 30184
rect 18785 30175 18843 30181
rect 18785 30172 18797 30175
rect 18288 30144 18797 30172
rect 18288 30132 18294 30144
rect 18785 30141 18797 30144
rect 18831 30141 18843 30175
rect 18785 30135 18843 30141
rect 19061 30175 19119 30181
rect 19061 30141 19073 30175
rect 19107 30172 19119 30175
rect 19426 30172 19432 30184
rect 19107 30144 19432 30172
rect 19107 30141 19119 30144
rect 19061 30135 19119 30141
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 20714 30132 20720 30184
rect 20772 30172 20778 30184
rect 22388 30172 22416 30212
rect 23089 30209 23101 30212
rect 23135 30209 23147 30243
rect 23089 30203 23147 30209
rect 23658 30200 23664 30252
rect 23716 30240 23722 30252
rect 24578 30240 24584 30252
rect 23716 30212 24584 30240
rect 23716 30200 23722 30212
rect 24578 30200 24584 30212
rect 24636 30240 24642 30252
rect 24673 30243 24731 30249
rect 24673 30240 24685 30243
rect 24636 30212 24685 30240
rect 24636 30200 24642 30212
rect 24673 30209 24685 30212
rect 24719 30209 24731 30243
rect 24673 30203 24731 30209
rect 20772 30144 22416 30172
rect 20772 30132 20778 30144
rect 22554 30132 22560 30184
rect 22612 30172 22618 30184
rect 22833 30175 22891 30181
rect 22833 30172 22845 30175
rect 22612 30144 22845 30172
rect 22612 30132 22618 30144
rect 22833 30141 22845 30144
rect 22879 30141 22891 30175
rect 24688 30172 24716 30203
rect 24854 30200 24860 30252
rect 24912 30200 24918 30252
rect 25332 30249 25360 30280
rect 25317 30243 25375 30249
rect 25317 30209 25329 30243
rect 25363 30209 25375 30243
rect 25317 30203 25375 30209
rect 25501 30243 25559 30249
rect 25501 30209 25513 30243
rect 25547 30209 25559 30243
rect 25608 30240 25636 30280
rect 26234 30268 26240 30320
rect 26292 30308 26298 30320
rect 27295 30311 27353 30317
rect 27295 30308 27307 30311
rect 26292 30280 27307 30308
rect 26292 30268 26298 30280
rect 27295 30277 27307 30280
rect 27341 30277 27353 30311
rect 27295 30271 27353 30277
rect 25958 30249 25964 30252
rect 25951 30243 25964 30249
rect 25951 30240 25963 30243
rect 25608 30212 25963 30240
rect 25501 30203 25559 30209
rect 25951 30209 25963 30212
rect 25951 30203 25964 30209
rect 25332 30172 25360 30203
rect 24688 30144 25360 30172
rect 25516 30172 25544 30203
rect 25958 30200 25964 30203
rect 26016 30200 26022 30252
rect 26050 30200 26056 30252
rect 26108 30240 26114 30252
rect 26145 30243 26203 30249
rect 26145 30240 26157 30243
rect 26108 30212 26157 30240
rect 26108 30200 26114 30212
rect 26145 30209 26157 30212
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27192 30243 27250 30249
rect 27192 30240 27204 30243
rect 27120 30212 27204 30240
rect 27120 30200 27126 30212
rect 27192 30209 27204 30212
rect 27238 30209 27250 30243
rect 27192 30203 27250 30209
rect 27982 30200 27988 30252
rect 28040 30200 28046 30252
rect 26786 30172 26792 30184
rect 25516 30144 26792 30172
rect 22833 30135 22891 30141
rect 26786 30132 26792 30144
rect 26844 30132 26850 30184
rect 22738 30104 22744 30116
rect 17788 30076 22744 30104
rect 17126 30036 17132 30048
rect 16172 30008 17132 30036
rect 16172 29996 16178 30008
rect 17126 29996 17132 30008
rect 17184 30036 17190 30048
rect 17494 30036 17500 30048
rect 17184 30008 17500 30036
rect 17184 29996 17190 30008
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 17586 29996 17592 30048
rect 17644 30036 17650 30048
rect 17788 30036 17816 30076
rect 22738 30064 22744 30076
rect 22796 30064 22802 30116
rect 17644 30008 17816 30036
rect 17644 29996 17650 30008
rect 18138 29996 18144 30048
rect 18196 30036 18202 30048
rect 18233 30039 18291 30045
rect 18233 30036 18245 30039
rect 18196 30008 18245 30036
rect 18196 29996 18202 30008
rect 18233 30005 18245 30008
rect 18279 30005 18291 30039
rect 18233 29999 18291 30005
rect 20073 30039 20131 30045
rect 20073 30005 20085 30039
rect 20119 30036 20131 30039
rect 21910 30036 21916 30048
rect 20119 30008 21916 30036
rect 20119 30005 20131 30008
rect 20073 29999 20131 30005
rect 21910 29996 21916 30008
rect 21968 29996 21974 30048
rect 23014 29996 23020 30048
rect 23072 30036 23078 30048
rect 24213 30039 24271 30045
rect 24213 30036 24225 30039
rect 23072 30008 24225 30036
rect 23072 29996 23078 30008
rect 24213 30005 24225 30008
rect 24259 30005 24271 30039
rect 24213 29999 24271 30005
rect 27798 29996 27804 30048
rect 27856 29996 27862 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 2774 29792 2780 29844
rect 2832 29792 2838 29844
rect 4062 29792 4068 29844
rect 4120 29832 4126 29844
rect 11054 29832 11060 29844
rect 4120 29804 11060 29832
rect 4120 29792 4126 29804
rect 11054 29792 11060 29804
rect 11112 29792 11118 29844
rect 11974 29792 11980 29844
rect 12032 29832 12038 29844
rect 13081 29835 13139 29841
rect 13081 29832 13093 29835
rect 12032 29804 13093 29832
rect 12032 29792 12038 29804
rect 13081 29801 13093 29804
rect 13127 29801 13139 29835
rect 13081 29795 13139 29801
rect 13541 29835 13599 29841
rect 13541 29801 13553 29835
rect 13587 29832 13599 29835
rect 13587 29804 16436 29832
rect 13587 29801 13599 29804
rect 13541 29795 13599 29801
rect 3234 29724 3240 29776
rect 3292 29764 3298 29776
rect 4433 29767 4491 29773
rect 4433 29764 4445 29767
rect 3292 29736 4445 29764
rect 3292 29724 3298 29736
rect 4433 29733 4445 29736
rect 4479 29764 4491 29767
rect 5258 29764 5264 29776
rect 4479 29736 5264 29764
rect 4479 29733 4491 29736
rect 4433 29727 4491 29733
rect 5258 29724 5264 29736
rect 5316 29724 5322 29776
rect 6086 29724 6092 29776
rect 6144 29724 6150 29776
rect 7745 29767 7803 29773
rect 7745 29733 7757 29767
rect 7791 29764 7803 29767
rect 8570 29764 8576 29776
rect 7791 29736 8576 29764
rect 7791 29733 7803 29736
rect 7745 29727 7803 29733
rect 8570 29724 8576 29736
rect 8628 29724 8634 29776
rect 14550 29724 14556 29776
rect 14608 29764 14614 29776
rect 14918 29764 14924 29776
rect 14608 29736 14924 29764
rect 14608 29724 14614 29736
rect 14918 29724 14924 29736
rect 14976 29724 14982 29776
rect 16408 29764 16436 29804
rect 16482 29792 16488 29844
rect 16540 29832 16546 29844
rect 17862 29832 17868 29844
rect 16540 29804 17868 29832
rect 16540 29792 16546 29804
rect 17862 29792 17868 29804
rect 17920 29792 17926 29844
rect 18046 29792 18052 29844
rect 18104 29832 18110 29844
rect 20809 29835 20867 29841
rect 20809 29832 20821 29835
rect 18104 29804 20821 29832
rect 18104 29792 18110 29804
rect 20809 29801 20821 29804
rect 20855 29801 20867 29835
rect 20809 29795 20867 29801
rect 21542 29792 21548 29844
rect 21600 29832 21606 29844
rect 22554 29832 22560 29844
rect 21600 29804 22560 29832
rect 21600 29792 21606 29804
rect 16758 29764 16764 29776
rect 16408 29736 16764 29764
rect 16758 29724 16764 29736
rect 16816 29724 16822 29776
rect 2133 29699 2191 29705
rect 2133 29665 2145 29699
rect 2179 29696 2191 29699
rect 3142 29696 3148 29708
rect 2179 29668 3148 29696
rect 2179 29665 2191 29668
rect 2133 29659 2191 29665
rect 3142 29656 3148 29668
rect 3200 29656 3206 29708
rect 5718 29656 5724 29708
rect 5776 29656 5782 29708
rect 7377 29699 7435 29705
rect 6564 29668 7328 29696
rect 2406 29588 2412 29640
rect 2464 29588 2470 29640
rect 4065 29631 4123 29637
rect 2608 29600 2774 29628
rect 1946 29520 1952 29572
rect 2004 29560 2010 29572
rect 2608 29569 2636 29600
rect 2593 29563 2651 29569
rect 2593 29560 2605 29563
rect 2004 29532 2605 29560
rect 2004 29520 2010 29532
rect 2593 29529 2605 29532
rect 2639 29529 2651 29563
rect 2746 29560 2774 29600
rect 4065 29597 4077 29631
rect 4111 29628 4123 29631
rect 4154 29628 4160 29640
rect 4111 29600 4160 29628
rect 4111 29597 4123 29600
rect 4065 29591 4123 29597
rect 4154 29588 4160 29600
rect 4212 29628 4218 29640
rect 4893 29631 4951 29637
rect 4893 29628 4905 29631
rect 4212 29600 4905 29628
rect 4212 29588 4218 29600
rect 4893 29597 4905 29600
rect 4939 29628 4951 29631
rect 4982 29628 4988 29640
rect 4939 29600 4988 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 5350 29588 5356 29640
rect 5408 29628 5414 29640
rect 6564 29637 6592 29668
rect 6549 29631 6607 29637
rect 6549 29628 6561 29631
rect 5408 29600 6561 29628
rect 5408 29588 5414 29600
rect 6549 29597 6561 29600
rect 6595 29597 6607 29631
rect 6549 29591 6607 29597
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29597 6975 29631
rect 7300 29628 7328 29668
rect 7377 29665 7389 29699
rect 7423 29696 7435 29699
rect 8294 29696 8300 29708
rect 7423 29668 8300 29696
rect 7423 29665 7435 29668
rect 7377 29659 7435 29665
rect 8294 29656 8300 29668
rect 8352 29656 8358 29708
rect 14090 29656 14096 29708
rect 14148 29696 14154 29708
rect 21836 29705 21864 29804
rect 22554 29792 22560 29804
rect 22612 29792 22618 29844
rect 22738 29792 22744 29844
rect 22796 29832 22802 29844
rect 23201 29835 23259 29841
rect 23201 29832 23213 29835
rect 22796 29804 23213 29832
rect 22796 29792 22802 29804
rect 23201 29801 23213 29804
rect 23247 29801 23259 29835
rect 23201 29795 23259 29801
rect 24228 29804 26096 29832
rect 24228 29764 24256 29804
rect 22940 29736 24256 29764
rect 26068 29764 26096 29804
rect 26142 29792 26148 29844
rect 26200 29832 26206 29844
rect 27617 29835 27675 29841
rect 27617 29832 27629 29835
rect 26200 29804 27629 29832
rect 26200 29792 26206 29804
rect 27617 29801 27629 29804
rect 27663 29801 27675 29835
rect 27617 29795 27675 29801
rect 26510 29764 26516 29776
rect 26068 29736 26516 29764
rect 21821 29699 21879 29705
rect 14148 29668 15148 29696
rect 14148 29656 14154 29668
rect 7466 29628 7472 29640
rect 7300 29600 7472 29628
rect 6917 29591 6975 29597
rect 5718 29560 5724 29572
rect 2746 29532 5724 29560
rect 2593 29523 2651 29529
rect 5718 29520 5724 29532
rect 5776 29520 5782 29572
rect 1486 29452 1492 29504
rect 1544 29492 1550 29504
rect 2038 29492 2044 29504
rect 1544 29464 2044 29492
rect 1544 29452 1550 29464
rect 2038 29452 2044 29464
rect 2096 29492 2102 29504
rect 2501 29495 2559 29501
rect 2501 29492 2513 29495
rect 2096 29464 2513 29492
rect 2096 29452 2102 29464
rect 2501 29461 2513 29464
rect 2547 29461 2559 29495
rect 2501 29455 2559 29461
rect 4433 29495 4491 29501
rect 4433 29461 4445 29495
rect 4479 29492 4491 29495
rect 5166 29492 5172 29504
rect 4479 29464 5172 29492
rect 4479 29461 4491 29464
rect 4433 29455 4491 29461
rect 5166 29452 5172 29464
rect 5224 29492 5230 29504
rect 6932 29501 6960 29591
rect 7466 29588 7472 29600
rect 7524 29628 7530 29640
rect 8205 29631 8263 29637
rect 8205 29628 8217 29631
rect 7524 29600 8217 29628
rect 7524 29588 7530 29600
rect 8205 29597 8217 29600
rect 8251 29597 8263 29631
rect 8205 29591 8263 29597
rect 8573 29631 8631 29637
rect 8573 29597 8585 29631
rect 8619 29597 8631 29631
rect 8573 29591 8631 29597
rect 5261 29495 5319 29501
rect 5261 29492 5273 29495
rect 5224 29464 5273 29492
rect 5224 29452 5230 29464
rect 5261 29461 5273 29464
rect 5307 29492 5319 29495
rect 6089 29495 6147 29501
rect 6089 29492 6101 29495
rect 5307 29464 6101 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 6089 29461 6101 29464
rect 6135 29492 6147 29495
rect 6917 29495 6975 29501
rect 6917 29492 6929 29495
rect 6135 29464 6929 29492
rect 6135 29461 6147 29464
rect 6089 29455 6147 29461
rect 6917 29461 6929 29464
rect 6963 29492 6975 29495
rect 7745 29495 7803 29501
rect 7745 29492 7757 29495
rect 6963 29464 7757 29492
rect 6963 29461 6975 29464
rect 6917 29455 6975 29461
rect 7745 29461 7757 29464
rect 7791 29492 7803 29495
rect 8478 29492 8484 29504
rect 7791 29464 8484 29492
rect 7791 29461 7803 29464
rect 7745 29455 7803 29461
rect 8478 29452 8484 29464
rect 8536 29492 8542 29504
rect 8588 29501 8616 29591
rect 9122 29588 9128 29640
rect 9180 29628 9186 29640
rect 9585 29631 9643 29637
rect 9585 29628 9597 29631
rect 9180 29600 9597 29628
rect 9180 29588 9186 29600
rect 9585 29597 9597 29600
rect 9631 29628 9643 29631
rect 11238 29628 11244 29640
rect 9631 29600 11244 29628
rect 9631 29597 9643 29600
rect 9585 29591 9643 29597
rect 11238 29588 11244 29600
rect 11296 29628 11302 29640
rect 11701 29631 11759 29637
rect 11701 29628 11713 29631
rect 11296 29600 11713 29628
rect 11296 29588 11302 29600
rect 11701 29597 11713 29600
rect 11747 29597 11759 29631
rect 11701 29591 11759 29597
rect 13722 29588 13728 29640
rect 13780 29588 13786 29640
rect 14274 29588 14280 29640
rect 14332 29628 14338 29640
rect 14550 29628 14556 29640
rect 14332 29600 14556 29628
rect 14332 29588 14338 29600
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 15010 29588 15016 29640
rect 15068 29588 15074 29640
rect 15120 29628 15148 29668
rect 21821 29665 21833 29699
rect 21867 29665 21879 29699
rect 21821 29659 21879 29665
rect 15269 29631 15327 29637
rect 15269 29628 15281 29631
rect 15120 29600 15281 29628
rect 15269 29597 15281 29600
rect 15315 29597 15327 29631
rect 15269 29591 15327 29597
rect 16390 29588 16396 29640
rect 16448 29588 16454 29640
rect 17126 29588 17132 29640
rect 17184 29588 17190 29640
rect 17218 29588 17224 29640
rect 17276 29628 17282 29640
rect 17276 29600 19334 29628
rect 17276 29588 17282 29600
rect 9852 29563 9910 29569
rect 9852 29529 9864 29563
rect 9898 29560 9910 29563
rect 11968 29563 12026 29569
rect 9898 29532 11928 29560
rect 9898 29529 9910 29532
rect 9852 29523 9910 29529
rect 11900 29504 11928 29532
rect 11968 29529 11980 29563
rect 12014 29560 12026 29563
rect 12250 29560 12256 29572
rect 12014 29532 12256 29560
rect 12014 29529 12026 29532
rect 11968 29523 12026 29529
rect 12250 29520 12256 29532
rect 12308 29520 12314 29572
rect 14369 29563 14427 29569
rect 14369 29529 14381 29563
rect 14415 29560 14427 29563
rect 15930 29560 15936 29572
rect 14415 29532 15936 29560
rect 14415 29529 14427 29532
rect 14369 29523 14427 29529
rect 15930 29520 15936 29532
rect 15988 29520 15994 29572
rect 16114 29520 16120 29572
rect 16172 29560 16178 29572
rect 16408 29560 16436 29588
rect 16172 29532 16712 29560
rect 16172 29520 16178 29532
rect 8573 29495 8631 29501
rect 8573 29492 8585 29495
rect 8536 29464 8585 29492
rect 8536 29452 8542 29464
rect 8573 29461 8585 29464
rect 8619 29461 8631 29495
rect 8573 29455 8631 29461
rect 10134 29452 10140 29504
rect 10192 29492 10198 29504
rect 10965 29495 11023 29501
rect 10965 29492 10977 29495
rect 10192 29464 10977 29492
rect 10192 29452 10198 29464
rect 10965 29461 10977 29464
rect 11011 29461 11023 29495
rect 10965 29455 11023 29461
rect 11882 29452 11888 29504
rect 11940 29452 11946 29504
rect 15470 29452 15476 29504
rect 15528 29492 15534 29504
rect 16393 29495 16451 29501
rect 16393 29492 16405 29495
rect 15528 29464 16405 29492
rect 15528 29452 15534 29464
rect 16393 29461 16405 29464
rect 16439 29461 16451 29495
rect 16684 29492 16712 29532
rect 16942 29520 16948 29572
rect 17000 29560 17006 29572
rect 17374 29563 17432 29569
rect 17374 29560 17386 29563
rect 17000 29532 17386 29560
rect 17000 29520 17006 29532
rect 17374 29529 17386 29532
rect 17420 29529 17432 29563
rect 19306 29560 19334 29600
rect 19426 29588 19432 29640
rect 19484 29588 19490 29640
rect 19518 29588 19524 29640
rect 19576 29628 19582 29640
rect 19685 29631 19743 29637
rect 19685 29628 19697 29631
rect 19576 29600 19697 29628
rect 19576 29588 19582 29600
rect 19685 29597 19697 29600
rect 19731 29597 19743 29631
rect 19685 29591 19743 29597
rect 21910 29588 21916 29640
rect 21968 29628 21974 29640
rect 22077 29631 22135 29637
rect 22077 29628 22089 29631
rect 21968 29600 22089 29628
rect 21968 29588 21974 29600
rect 22077 29597 22089 29600
rect 22123 29597 22135 29631
rect 22077 29591 22135 29597
rect 22940 29560 22968 29736
rect 26510 29724 26516 29736
rect 26568 29764 26574 29776
rect 26973 29767 27031 29773
rect 26973 29764 26985 29767
rect 26568 29736 26985 29764
rect 26568 29724 26574 29736
rect 26973 29733 26985 29736
rect 27019 29733 27031 29767
rect 26973 29727 27031 29733
rect 23658 29588 23664 29640
rect 23716 29588 23722 29640
rect 23842 29588 23848 29640
rect 23900 29588 23906 29640
rect 24578 29588 24584 29640
rect 24636 29628 24642 29640
rect 25133 29631 25191 29637
rect 25133 29628 25145 29631
rect 24636 29600 25145 29628
rect 24636 29588 24642 29600
rect 25133 29597 25145 29600
rect 25179 29597 25191 29631
rect 25133 29591 25191 29597
rect 26602 29588 26608 29640
rect 26660 29628 26666 29640
rect 27157 29631 27215 29637
rect 27157 29628 27169 29631
rect 26660 29600 27169 29628
rect 26660 29588 26666 29600
rect 27157 29597 27169 29600
rect 27203 29597 27215 29631
rect 27157 29591 27215 29597
rect 27614 29588 27620 29640
rect 27672 29628 27678 29640
rect 27801 29631 27859 29637
rect 27801 29628 27813 29631
rect 27672 29600 27813 29628
rect 27672 29588 27678 29600
rect 27801 29597 27813 29600
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 19306 29532 22968 29560
rect 23124 29532 23336 29560
rect 17374 29523 17432 29529
rect 18509 29495 18567 29501
rect 18509 29492 18521 29495
rect 16684 29464 18521 29492
rect 16393 29455 16451 29461
rect 18509 29461 18521 29464
rect 18555 29461 18567 29495
rect 18509 29455 18567 29461
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 20530 29492 20536 29504
rect 19392 29464 20536 29492
rect 19392 29452 19398 29464
rect 20530 29452 20536 29464
rect 20588 29452 20594 29504
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 23124 29492 23152 29532
rect 20680 29464 23152 29492
rect 23308 29492 23336 29532
rect 24486 29520 24492 29572
rect 24544 29560 24550 29572
rect 25378 29563 25436 29569
rect 25378 29560 25390 29563
rect 24544 29532 25390 29560
rect 24544 29520 24550 29532
rect 25378 29529 25390 29532
rect 25424 29529 25436 29563
rect 25378 29523 25436 29529
rect 26513 29495 26571 29501
rect 26513 29492 26525 29495
rect 23308 29464 26525 29492
rect 20680 29452 20686 29464
rect 26513 29461 26525 29464
rect 26559 29461 26571 29495
rect 26513 29455 26571 29461
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 2590 29248 2596 29300
rect 2648 29288 2654 29300
rect 2869 29291 2927 29297
rect 2869 29288 2881 29291
rect 2648 29260 2881 29288
rect 2648 29248 2654 29260
rect 2869 29257 2881 29260
rect 2915 29257 2927 29291
rect 2869 29251 2927 29257
rect 5077 29291 5135 29297
rect 5077 29257 5089 29291
rect 5123 29288 5135 29291
rect 5166 29288 5172 29300
rect 5123 29260 5172 29288
rect 5123 29257 5135 29260
rect 5077 29251 5135 29257
rect 3786 29180 3792 29232
rect 3844 29180 3850 29232
rect 3970 29180 3976 29232
rect 4028 29180 4034 29232
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 4798 29152 4804 29164
rect 1627 29124 4804 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 4798 29112 4804 29124
rect 4856 29112 4862 29164
rect 5092 29161 5120 29251
rect 5166 29248 5172 29260
rect 5224 29288 5230 29300
rect 5997 29291 6055 29297
rect 5997 29288 6009 29291
rect 5224 29260 6009 29288
rect 5224 29248 5230 29260
rect 5997 29257 6009 29260
rect 6043 29257 6055 29291
rect 5997 29251 6055 29257
rect 7653 29291 7711 29297
rect 7653 29257 7665 29291
rect 7699 29257 7711 29291
rect 7653 29251 7711 29257
rect 7668 29220 7696 29251
rect 8478 29248 8484 29300
rect 8536 29288 8542 29300
rect 8573 29291 8631 29297
rect 8573 29288 8585 29291
rect 8536 29260 8585 29288
rect 8536 29248 8542 29260
rect 8573 29257 8585 29260
rect 8619 29288 8631 29291
rect 9122 29288 9128 29300
rect 8619 29260 9128 29288
rect 8619 29257 8631 29260
rect 8573 29251 8631 29257
rect 9122 29248 9128 29260
rect 9180 29288 9186 29300
rect 9401 29291 9459 29297
rect 9401 29288 9413 29291
rect 9180 29260 9413 29288
rect 9180 29248 9186 29260
rect 9401 29257 9413 29260
rect 9447 29257 9459 29291
rect 9401 29251 9459 29257
rect 11701 29291 11759 29297
rect 11701 29257 11713 29291
rect 11747 29288 11759 29291
rect 12713 29291 12771 29297
rect 11747 29260 12434 29288
rect 11747 29257 11759 29260
rect 11701 29251 11759 29257
rect 12066 29220 12072 29232
rect 6104 29192 12072 29220
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 5258 29112 5264 29164
rect 5316 29152 5322 29164
rect 5997 29155 6055 29161
rect 5997 29152 6009 29155
rect 5316 29124 6009 29152
rect 5316 29112 5322 29124
rect 5997 29121 6009 29124
rect 6043 29121 6055 29155
rect 5997 29115 6055 29121
rect 4706 29044 4712 29096
rect 4764 29044 4770 29096
rect 4982 29044 4988 29096
rect 5040 29084 5046 29096
rect 5629 29087 5687 29093
rect 5629 29084 5641 29087
rect 5040 29056 5641 29084
rect 5040 29044 5046 29056
rect 5629 29053 5641 29056
rect 5675 29084 5687 29087
rect 6104 29084 6132 29192
rect 12066 29180 12072 29192
rect 12124 29180 12130 29232
rect 12406 29220 12434 29260
rect 12713 29257 12725 29291
rect 12759 29288 12771 29291
rect 13541 29291 13599 29297
rect 13541 29288 13553 29291
rect 12759 29260 13553 29288
rect 12759 29257 12771 29260
rect 12713 29251 12771 29257
rect 13541 29257 13553 29260
rect 13587 29288 13599 29291
rect 13630 29288 13636 29300
rect 13587 29260 13636 29288
rect 13587 29257 13599 29260
rect 13541 29251 13599 29257
rect 13630 29248 13636 29260
rect 13688 29248 13694 29300
rect 14366 29248 14372 29300
rect 14424 29288 14430 29300
rect 14737 29291 14795 29297
rect 14737 29288 14749 29291
rect 14424 29260 14749 29288
rect 14424 29248 14430 29260
rect 14737 29257 14749 29260
rect 14783 29257 14795 29291
rect 14737 29251 14795 29257
rect 15378 29248 15384 29300
rect 15436 29288 15442 29300
rect 16209 29291 16267 29297
rect 15436 29260 15608 29288
rect 15436 29248 15442 29260
rect 14090 29220 14096 29232
rect 12406 29192 14096 29220
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 14826 29180 14832 29232
rect 14884 29220 14890 29232
rect 15194 29220 15200 29232
rect 14884 29192 15200 29220
rect 14884 29180 14890 29192
rect 15194 29180 15200 29192
rect 15252 29180 15258 29232
rect 6730 29112 6736 29164
rect 6788 29112 6794 29164
rect 7009 29155 7067 29161
rect 7009 29121 7021 29155
rect 7055 29152 7067 29155
rect 7190 29152 7196 29164
rect 7055 29124 7196 29152
rect 7055 29121 7067 29124
rect 7009 29115 7067 29121
rect 7190 29112 7196 29124
rect 7248 29112 7254 29164
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29152 7527 29155
rect 7558 29152 7564 29164
rect 7515 29124 7564 29152
rect 7515 29121 7527 29124
rect 7469 29115 7527 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 8205 29155 8263 29161
rect 8205 29121 8217 29155
rect 8251 29152 8263 29155
rect 8294 29152 8300 29164
rect 8251 29124 8300 29152
rect 8251 29121 8263 29124
rect 8205 29115 8263 29121
rect 8294 29112 8300 29124
rect 8352 29152 8358 29164
rect 8754 29152 8760 29164
rect 8352 29124 8760 29152
rect 8352 29112 8358 29124
rect 8754 29112 8760 29124
rect 8812 29152 8818 29164
rect 9033 29155 9091 29161
rect 9033 29152 9045 29155
rect 8812 29124 9045 29152
rect 8812 29112 8818 29124
rect 9033 29121 9045 29124
rect 9079 29152 9091 29155
rect 9214 29152 9220 29164
rect 9079 29124 9220 29152
rect 9079 29121 9091 29124
rect 9033 29115 9091 29121
rect 9214 29112 9220 29124
rect 9272 29112 9278 29164
rect 11885 29155 11943 29161
rect 11885 29121 11897 29155
rect 11931 29152 11943 29155
rect 12158 29152 12164 29164
rect 11931 29124 12164 29152
rect 11931 29121 11943 29124
rect 11885 29115 11943 29121
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 12713 29155 12771 29161
rect 12713 29121 12725 29155
rect 12759 29152 12771 29155
rect 13541 29155 13599 29161
rect 13541 29152 13553 29155
rect 12759 29124 13553 29152
rect 12759 29121 12771 29124
rect 12713 29115 12771 29121
rect 13541 29121 13553 29124
rect 13587 29152 13599 29155
rect 13630 29152 13636 29164
rect 13587 29124 13636 29152
rect 13587 29121 13599 29124
rect 13541 29115 13599 29121
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 15378 29152 15384 29164
rect 13780 29124 15384 29152
rect 13780 29112 13786 29124
rect 15378 29112 15384 29124
rect 15436 29112 15442 29164
rect 5675 29056 6132 29084
rect 5675 29053 5687 29056
rect 5629 29047 5687 29053
rect 6546 29044 6552 29096
rect 6604 29044 6610 29096
rect 10229 29087 10287 29093
rect 10229 29084 10241 29087
rect 8496 29056 10241 29084
rect 4154 28976 4160 29028
rect 4212 28976 4218 29028
rect 5534 28976 5540 29028
rect 5592 29016 5598 29028
rect 6730 29016 6736 29028
rect 5592 28988 6736 29016
rect 5592 28976 5598 28988
rect 6730 28976 6736 28988
rect 6788 29016 6794 29028
rect 6917 29019 6975 29025
rect 6917 29016 6929 29019
rect 6788 28988 6929 29016
rect 6788 28976 6794 28988
rect 6917 28985 6929 28988
rect 6963 28985 6975 29019
rect 8496 29016 8524 29056
rect 10229 29053 10241 29056
rect 10275 29084 10287 29087
rect 10275 29056 10824 29084
rect 10275 29053 10287 29056
rect 10229 29047 10287 29053
rect 6917 28979 6975 28985
rect 7024 28988 8524 29016
rect 7024 28960 7052 28988
rect 8570 28976 8576 29028
rect 8628 29016 8634 29028
rect 9030 29016 9036 29028
rect 8628 28988 9036 29016
rect 8628 28976 8634 28988
rect 9030 28976 9036 28988
rect 9088 29016 9094 29028
rect 9401 29019 9459 29025
rect 9401 29016 9413 29019
rect 9088 28988 9413 29016
rect 9088 28976 9094 28988
rect 9401 28985 9413 28988
rect 9447 28985 9459 29019
rect 9401 28979 9459 28985
rect 10502 28976 10508 29028
rect 10560 28976 10566 29028
rect 10686 28976 10692 29028
rect 10744 28976 10750 29028
rect 10796 29016 10824 29056
rect 12342 29044 12348 29096
rect 12400 29084 12406 29096
rect 13173 29087 13231 29093
rect 13173 29084 13185 29087
rect 12400 29056 13185 29084
rect 12400 29044 12406 29056
rect 13173 29053 13185 29056
rect 13219 29053 13231 29087
rect 14277 29087 14335 29093
rect 14277 29084 14289 29087
rect 13173 29047 13231 29053
rect 13464 29056 14289 29084
rect 13464 29016 13492 29056
rect 14277 29053 14289 29056
rect 14323 29084 14335 29087
rect 14458 29084 14464 29096
rect 14323 29056 14464 29084
rect 14323 29053 14335 29056
rect 14277 29047 14335 29053
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 15470 29084 15476 29096
rect 14568 29056 15476 29084
rect 14568 29016 14596 29056
rect 15470 29044 15476 29056
rect 15528 29044 15534 29096
rect 10796 28988 12664 29016
rect 3973 28951 4031 28957
rect 3973 28917 3985 28951
rect 4019 28948 4031 28951
rect 5442 28948 5448 28960
rect 4019 28920 5448 28948
rect 4019 28917 4031 28920
rect 3973 28911 4031 28917
rect 5442 28908 5448 28920
rect 5500 28908 5506 28960
rect 7006 28908 7012 28960
rect 7064 28908 7070 28960
rect 12636 28948 12664 28988
rect 12820 28988 13492 29016
rect 14292 28988 14596 29016
rect 14645 29019 14703 29025
rect 12820 28948 12848 28988
rect 14292 28960 14320 28988
rect 14645 28985 14657 29019
rect 14691 29016 14703 29019
rect 14826 29016 14832 29028
rect 14691 28988 14832 29016
rect 14691 28985 14703 28988
rect 14645 28979 14703 28985
rect 14826 28976 14832 28988
rect 14884 28976 14890 29028
rect 15194 28976 15200 29028
rect 15252 29016 15258 29028
rect 15580 29016 15608 29260
rect 16209 29257 16221 29291
rect 16255 29288 16267 29291
rect 16482 29288 16488 29300
rect 16255 29260 16488 29288
rect 16255 29257 16267 29260
rect 16209 29251 16267 29257
rect 16482 29248 16488 29260
rect 16540 29248 16546 29300
rect 16666 29248 16672 29300
rect 16724 29288 16730 29300
rect 19334 29288 19340 29300
rect 16724 29260 19340 29288
rect 16724 29248 16730 29260
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19521 29291 19579 29297
rect 19521 29257 19533 29291
rect 19567 29288 19579 29291
rect 20898 29288 20904 29300
rect 19567 29260 20904 29288
rect 19567 29257 19579 29260
rect 19521 29251 19579 29257
rect 20898 29248 20904 29260
rect 20956 29248 20962 29300
rect 21453 29291 21511 29297
rect 21453 29257 21465 29291
rect 21499 29257 21511 29291
rect 21453 29251 21511 29257
rect 22005 29291 22063 29297
rect 22005 29257 22017 29291
rect 22051 29288 22063 29291
rect 22278 29288 22284 29300
rect 22051 29260 22284 29288
rect 22051 29257 22063 29260
rect 22005 29251 22063 29257
rect 16758 29180 16764 29232
rect 16816 29220 16822 29232
rect 17558 29223 17616 29229
rect 17558 29220 17570 29223
rect 16816 29192 17570 29220
rect 16816 29180 16822 29192
rect 17558 29189 17570 29192
rect 17604 29189 17616 29223
rect 17558 29183 17616 29189
rect 18138 29180 18144 29232
rect 18196 29220 18202 29232
rect 18598 29220 18604 29232
rect 18196 29192 18604 29220
rect 18196 29180 18202 29192
rect 18598 29180 18604 29192
rect 18656 29180 18662 29232
rect 18966 29180 18972 29232
rect 19024 29220 19030 29232
rect 19153 29223 19211 29229
rect 19153 29220 19165 29223
rect 19024 29192 19165 29220
rect 19024 29180 19030 29192
rect 19153 29189 19165 29192
rect 19199 29189 19211 29223
rect 21468 29220 21496 29251
rect 22278 29248 22284 29260
rect 22336 29248 22342 29300
rect 22830 29248 22836 29300
rect 22888 29288 22894 29300
rect 24946 29288 24952 29300
rect 22888 29260 24952 29288
rect 22888 29248 22894 29260
rect 24946 29248 24952 29260
rect 25004 29248 25010 29300
rect 25792 29260 26004 29288
rect 19153 29183 19211 29189
rect 19352 29192 21496 29220
rect 15749 29155 15807 29161
rect 15749 29121 15761 29155
rect 15795 29152 15807 29155
rect 16040 29152 16160 29156
rect 17034 29152 17040 29164
rect 15795 29128 17040 29152
rect 15795 29124 16068 29128
rect 16132 29124 17040 29128
rect 15795 29121 15807 29124
rect 15749 29115 15807 29121
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 17126 29112 17132 29164
rect 17184 29152 17190 29164
rect 19352 29161 19380 29192
rect 21542 29180 21548 29232
rect 21600 29220 21606 29232
rect 25792 29220 25820 29260
rect 21600 29192 25820 29220
rect 21600 29180 21606 29192
rect 25866 29180 25872 29232
rect 25924 29180 25930 29232
rect 25976 29220 26004 29260
rect 27154 29248 27160 29300
rect 27212 29288 27218 29300
rect 27295 29291 27353 29297
rect 27295 29288 27307 29291
rect 27212 29260 27307 29288
rect 27212 29248 27218 29260
rect 27295 29257 27307 29260
rect 27341 29257 27353 29291
rect 27295 29251 27353 29257
rect 26694 29220 26700 29232
rect 25976 29192 26700 29220
rect 17313 29155 17371 29161
rect 17313 29152 17325 29155
rect 17184 29124 17325 29152
rect 17184 29112 17190 29124
rect 17313 29121 17325 29124
rect 17359 29152 17371 29155
rect 19337 29155 19395 29161
rect 17359 29124 19104 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 17218 29084 17224 29096
rect 15948 29056 17224 29084
rect 15948 29016 15976 29056
rect 17218 29044 17224 29056
rect 17276 29044 17282 29096
rect 15252 28988 15608 29016
rect 15856 28988 15976 29016
rect 16117 29019 16175 29025
rect 15252 28976 15258 28988
rect 12636 28920 12848 28948
rect 14274 28908 14280 28960
rect 14332 28908 14338 28960
rect 14366 28908 14372 28960
rect 14424 28948 14430 28960
rect 15856 28948 15884 28988
rect 16117 28985 16129 29019
rect 16163 29016 16175 29019
rect 16206 29016 16212 29028
rect 16163 28988 16212 29016
rect 16163 28985 16175 28988
rect 16117 28979 16175 28985
rect 16206 28976 16212 28988
rect 16264 28976 16270 29028
rect 14424 28920 15884 28948
rect 14424 28908 14430 28920
rect 15930 28908 15936 28960
rect 15988 28948 15994 28960
rect 18230 28948 18236 28960
rect 15988 28920 18236 28948
rect 15988 28908 15994 28920
rect 18230 28908 18236 28920
rect 18288 28908 18294 28960
rect 18598 28908 18604 28960
rect 18656 28948 18662 28960
rect 18693 28951 18751 28957
rect 18693 28948 18705 28951
rect 18656 28920 18705 28948
rect 18656 28908 18662 28920
rect 18693 28917 18705 28920
rect 18739 28917 18751 28951
rect 19076 28948 19104 29124
rect 19337 29121 19349 29155
rect 19383 29121 19395 29155
rect 19337 29115 19395 29121
rect 19352 29084 19380 29115
rect 19426 29112 19432 29164
rect 19484 29152 19490 29164
rect 20073 29155 20131 29161
rect 20073 29152 20085 29155
rect 19484 29124 20085 29152
rect 19484 29112 19490 29124
rect 20073 29121 20085 29124
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 20340 29155 20398 29161
rect 20340 29121 20352 29155
rect 20386 29152 20398 29155
rect 21450 29152 21456 29164
rect 20386 29124 21456 29152
rect 20386 29121 20398 29124
rect 20340 29115 20398 29121
rect 21450 29112 21456 29124
rect 21508 29112 21514 29164
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22152 29124 22201 29152
rect 22152 29112 22158 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 22649 29115 22707 29121
rect 19168 29056 19380 29084
rect 19168 29028 19196 29056
rect 21082 29044 21088 29096
rect 21140 29084 21146 29096
rect 22664 29084 22692 29115
rect 22830 29112 22836 29164
rect 22888 29112 22894 29164
rect 24193 29155 24251 29161
rect 24193 29152 24205 29155
rect 23768 29124 24205 29152
rect 23658 29084 23664 29096
rect 21140 29056 23664 29084
rect 21140 29044 21146 29056
rect 23658 29044 23664 29056
rect 23716 29044 23722 29096
rect 19150 28976 19156 29028
rect 19208 28976 19214 29028
rect 23768 29016 23796 29124
rect 24193 29121 24205 29124
rect 24239 29121 24251 29155
rect 24193 29115 24251 29121
rect 25774 29112 25780 29164
rect 25832 29112 25838 29164
rect 25976 29161 26004 29192
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29121 26019 29155
rect 25961 29115 26019 29121
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29152 26479 29155
rect 26510 29152 26516 29164
rect 26467 29124 26516 29152
rect 26467 29121 26479 29124
rect 26421 29115 26479 29121
rect 26510 29112 26516 29124
rect 26568 29112 26574 29164
rect 26620 29161 26648 29192
rect 26694 29180 26700 29192
rect 26752 29180 26758 29232
rect 26605 29155 26663 29161
rect 26605 29121 26617 29155
rect 26651 29121 26663 29155
rect 27062 29152 27068 29164
rect 26605 29115 26663 29121
rect 26712 29124 27068 29152
rect 23937 29087 23995 29093
rect 23937 29084 23949 29087
rect 21008 28988 23796 29016
rect 23860 29056 23949 29084
rect 19702 28948 19708 28960
rect 19076 28920 19708 28948
rect 18693 28911 18751 28917
rect 19702 28908 19708 28920
rect 19760 28908 19766 28960
rect 20438 28908 20444 28960
rect 20496 28948 20502 28960
rect 21008 28948 21036 28988
rect 20496 28920 21036 28948
rect 20496 28908 20502 28920
rect 23474 28908 23480 28960
rect 23532 28908 23538 28960
rect 23658 28908 23664 28960
rect 23716 28948 23722 28960
rect 23860 28948 23888 29056
rect 23937 29053 23949 29056
rect 23983 29053 23995 29087
rect 23937 29047 23995 29053
rect 26234 29044 26240 29096
rect 26292 29084 26298 29096
rect 26712 29084 26740 29124
rect 27062 29112 27068 29124
rect 27120 29152 27126 29164
rect 27192 29155 27250 29161
rect 27192 29152 27204 29155
rect 27120 29124 27204 29152
rect 27120 29112 27126 29124
rect 27192 29121 27204 29124
rect 27238 29121 27250 29155
rect 27192 29115 27250 29121
rect 27890 29112 27896 29164
rect 27948 29152 27954 29164
rect 27985 29155 28043 29161
rect 27985 29152 27997 29155
rect 27948 29124 27997 29152
rect 27948 29112 27954 29124
rect 27985 29121 27997 29124
rect 28031 29121 28043 29155
rect 27985 29115 28043 29121
rect 26292 29056 26740 29084
rect 26292 29044 26298 29056
rect 24946 28976 24952 29028
rect 25004 29016 25010 29028
rect 25317 29019 25375 29025
rect 25317 29016 25329 29019
rect 25004 28988 25329 29016
rect 25004 28976 25010 28988
rect 25317 28985 25329 28988
rect 25363 28985 25375 29019
rect 25317 28979 25375 28985
rect 25590 28976 25596 29028
rect 25648 29016 25654 29028
rect 27801 29019 27859 29025
rect 27801 29016 27813 29019
rect 25648 28988 27813 29016
rect 25648 28976 25654 28988
rect 27801 28985 27813 28988
rect 27847 28985 27859 29019
rect 27801 28979 27859 28985
rect 23716 28920 23888 28948
rect 23716 28908 23722 28920
rect 25682 28908 25688 28960
rect 25740 28948 25746 28960
rect 26421 28951 26479 28957
rect 26421 28948 26433 28951
rect 25740 28920 26433 28948
rect 25740 28908 25746 28920
rect 26421 28917 26433 28920
rect 26467 28917 26479 28951
rect 26421 28911 26479 28917
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 7190 28704 7196 28756
rect 7248 28744 7254 28756
rect 15197 28747 15255 28753
rect 7248 28716 15148 28744
rect 7248 28704 7254 28716
rect 7742 28636 7748 28688
rect 7800 28676 7806 28688
rect 9309 28679 9367 28685
rect 7800 28648 8064 28676
rect 7800 28636 7806 28648
rect 3878 28568 3884 28620
rect 3936 28608 3942 28620
rect 8036 28617 8064 28648
rect 9309 28645 9321 28679
rect 9355 28676 9367 28679
rect 9674 28676 9680 28688
rect 9355 28648 9680 28676
rect 9355 28645 9367 28648
rect 9309 28639 9367 28645
rect 9674 28636 9680 28648
rect 9732 28636 9738 28688
rect 10962 28636 10968 28688
rect 11020 28676 11026 28688
rect 11057 28679 11115 28685
rect 11057 28676 11069 28679
rect 11020 28648 11069 28676
rect 11020 28636 11026 28648
rect 11057 28645 11069 28648
rect 11103 28676 11115 28679
rect 11885 28679 11943 28685
rect 11885 28676 11897 28679
rect 11103 28648 11897 28676
rect 11103 28645 11115 28648
rect 11057 28639 11115 28645
rect 11885 28645 11897 28648
rect 11931 28645 11943 28679
rect 11885 28639 11943 28645
rect 12544 28648 13952 28676
rect 8021 28611 8079 28617
rect 3936 28580 7972 28608
rect 3936 28568 3942 28580
rect 1765 28543 1823 28549
rect 1765 28509 1777 28543
rect 1811 28509 1823 28543
rect 1765 28503 1823 28509
rect 1780 28472 1808 28503
rect 1854 28500 1860 28552
rect 1912 28540 1918 28552
rect 2021 28543 2079 28549
rect 2021 28540 2033 28543
rect 1912 28512 2033 28540
rect 1912 28500 1918 28512
rect 2021 28509 2033 28512
rect 2067 28509 2079 28543
rect 2021 28503 2079 28509
rect 3234 28500 3240 28552
rect 3292 28540 3298 28552
rect 3973 28543 4031 28549
rect 3973 28540 3985 28543
rect 3292 28512 3985 28540
rect 3292 28500 3298 28512
rect 3973 28509 3985 28512
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 4249 28543 4307 28549
rect 4249 28509 4261 28543
rect 4295 28509 4307 28543
rect 4249 28503 4307 28509
rect 4264 28472 4292 28503
rect 4798 28500 4804 28552
rect 4856 28540 4862 28552
rect 5261 28543 5319 28549
rect 5261 28540 5273 28543
rect 4856 28512 5273 28540
rect 4856 28500 4862 28512
rect 5261 28509 5273 28512
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 6822 28500 6828 28552
rect 6880 28500 6886 28552
rect 7466 28500 7472 28552
rect 7524 28500 7530 28552
rect 7653 28543 7711 28549
rect 7653 28509 7665 28543
rect 7699 28509 7711 28543
rect 7944 28540 7972 28580
rect 8021 28577 8033 28611
rect 8067 28577 8079 28611
rect 11146 28608 11152 28620
rect 8021 28571 8079 28577
rect 9048 28580 11152 28608
rect 9048 28540 9076 28580
rect 11146 28568 11152 28580
rect 11204 28568 11210 28620
rect 12158 28568 12164 28620
rect 12216 28608 12222 28620
rect 12544 28608 12572 28648
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12216 28580 12572 28608
rect 12636 28580 13185 28608
rect 12216 28568 12222 28580
rect 7944 28512 9076 28540
rect 9125 28543 9183 28549
rect 7653 28503 7711 28509
rect 9125 28509 9137 28543
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 4982 28472 4988 28484
rect 1780 28444 1992 28472
rect 4264 28444 4988 28472
rect 1964 28416 1992 28444
rect 4982 28432 4988 28444
rect 5040 28432 5046 28484
rect 5074 28432 5080 28484
rect 5132 28472 5138 28484
rect 7668 28472 7696 28503
rect 9140 28472 9168 28503
rect 9858 28500 9864 28552
rect 9916 28500 9922 28552
rect 10229 28543 10287 28549
rect 10229 28509 10241 28543
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28540 10747 28543
rect 11517 28543 11575 28549
rect 11517 28540 11529 28543
rect 10735 28512 11529 28540
rect 10735 28509 10747 28512
rect 10689 28503 10747 28509
rect 11517 28509 11529 28512
rect 11563 28540 11575 28543
rect 11882 28540 11888 28552
rect 11563 28512 11888 28540
rect 11563 28509 11575 28512
rect 11517 28503 11575 28509
rect 9674 28472 9680 28484
rect 5132 28444 7696 28472
rect 9054 28444 9680 28472
rect 5132 28432 5138 28444
rect 1946 28364 1952 28416
rect 2004 28364 2010 28416
rect 3142 28364 3148 28416
rect 3200 28364 3206 28416
rect 4246 28364 4252 28416
rect 4304 28364 4310 28416
rect 4338 28364 4344 28416
rect 4396 28404 4402 28416
rect 7653 28407 7711 28413
rect 7653 28404 7665 28407
rect 4396 28376 7665 28404
rect 4396 28364 4402 28376
rect 7653 28373 7665 28376
rect 7699 28404 7711 28407
rect 9054 28404 9082 28444
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 7699 28376 9082 28404
rect 7699 28373 7711 28376
rect 7653 28367 7711 28373
rect 9122 28364 9128 28416
rect 9180 28404 9186 28416
rect 10244 28413 10272 28503
rect 11882 28500 11888 28512
rect 11940 28540 11946 28552
rect 12342 28540 12348 28552
rect 11940 28512 12348 28540
rect 11940 28500 11946 28512
rect 12342 28500 12348 28512
rect 12400 28540 12406 28552
rect 12636 28540 12664 28580
rect 13173 28577 13185 28580
rect 13219 28577 13231 28611
rect 13173 28571 13231 28577
rect 12400 28512 12664 28540
rect 12713 28543 12771 28549
rect 12400 28500 12406 28512
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13630 28540 13636 28552
rect 13587 28512 13636 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 10229 28407 10287 28413
rect 10229 28404 10241 28407
rect 9180 28376 10241 28404
rect 9180 28364 9186 28376
rect 10229 28373 10241 28376
rect 10275 28404 10287 28407
rect 10962 28404 10968 28416
rect 10275 28376 10968 28404
rect 10275 28373 10287 28376
rect 10229 28367 10287 28373
rect 10962 28364 10968 28376
rect 11020 28404 11026 28416
rect 11057 28407 11115 28413
rect 11057 28404 11069 28407
rect 11020 28376 11069 28404
rect 11020 28364 11026 28376
rect 11057 28373 11069 28376
rect 11103 28404 11115 28407
rect 11885 28407 11943 28413
rect 11885 28404 11897 28407
rect 11103 28376 11897 28404
rect 11103 28373 11115 28376
rect 11057 28367 11115 28373
rect 11885 28373 11897 28376
rect 11931 28404 11943 28407
rect 12618 28404 12624 28416
rect 11931 28376 12624 28404
rect 11931 28373 11943 28376
rect 11885 28367 11943 28373
rect 12618 28364 12624 28376
rect 12676 28404 12682 28416
rect 12728 28413 12756 28503
rect 13556 28413 13584 28503
rect 13630 28500 13636 28512
rect 13688 28500 13694 28552
rect 13924 28540 13952 28648
rect 13998 28636 14004 28688
rect 14056 28676 14062 28688
rect 14642 28676 14648 28688
rect 14056 28648 14648 28676
rect 14056 28636 14062 28648
rect 14642 28636 14648 28648
rect 14700 28676 14706 28688
rect 15013 28679 15071 28685
rect 15013 28676 15025 28679
rect 14700 28648 15025 28676
rect 14700 28636 14706 28648
rect 15013 28645 15025 28648
rect 15059 28645 15071 28679
rect 15120 28676 15148 28716
rect 15197 28713 15209 28747
rect 15243 28744 15255 28747
rect 16022 28744 16028 28756
rect 15243 28716 16028 28744
rect 15243 28713 15255 28716
rect 15197 28707 15255 28713
rect 16022 28704 16028 28716
rect 16080 28704 16086 28756
rect 17129 28747 17187 28753
rect 17129 28713 17141 28747
rect 17175 28744 17187 28747
rect 21082 28744 21088 28756
rect 17175 28716 21088 28744
rect 17175 28713 17187 28716
rect 17129 28707 17187 28713
rect 21082 28704 21088 28716
rect 21140 28704 21146 28756
rect 21450 28704 21456 28756
rect 21508 28704 21514 28756
rect 22281 28747 22339 28753
rect 22281 28713 22293 28747
rect 22327 28744 22339 28747
rect 23842 28744 23848 28756
rect 22327 28716 23848 28744
rect 22327 28713 22339 28716
rect 22281 28707 22339 28713
rect 23842 28704 23848 28716
rect 23900 28704 23906 28756
rect 26050 28744 26056 28756
rect 24596 28716 26056 28744
rect 17402 28676 17408 28688
rect 15120 28648 17408 28676
rect 15013 28639 15071 28645
rect 17402 28636 17408 28648
rect 17460 28636 17466 28688
rect 17954 28636 17960 28688
rect 18012 28676 18018 28688
rect 18690 28676 18696 28688
rect 18012 28648 18696 28676
rect 18012 28636 18018 28648
rect 18690 28636 18696 28648
rect 18748 28636 18754 28688
rect 18785 28679 18843 28685
rect 18785 28645 18797 28679
rect 18831 28676 18843 28679
rect 18966 28676 18972 28688
rect 18831 28648 18972 28676
rect 18831 28645 18843 28648
rect 18785 28639 18843 28645
rect 18966 28636 18972 28648
rect 19024 28636 19030 28688
rect 23569 28679 23627 28685
rect 23569 28645 23581 28679
rect 23615 28676 23627 28679
rect 24596 28676 24624 28716
rect 26050 28704 26056 28716
rect 26108 28704 26114 28756
rect 23615 28648 24624 28676
rect 25961 28679 26019 28685
rect 23615 28645 23627 28648
rect 23569 28639 23627 28645
rect 25961 28645 25973 28679
rect 26007 28676 26019 28679
rect 26234 28676 26240 28688
rect 26007 28648 26240 28676
rect 26007 28645 26019 28648
rect 25961 28639 26019 28645
rect 26234 28636 26240 28648
rect 26292 28636 26298 28688
rect 14090 28568 14096 28620
rect 14148 28608 14154 28620
rect 14148 28580 19748 28608
rect 14148 28568 14154 28580
rect 13924 28512 15608 28540
rect 14737 28475 14795 28481
rect 14737 28441 14749 28475
rect 14783 28472 14795 28475
rect 15580 28472 15608 28512
rect 15654 28500 15660 28552
rect 15712 28500 15718 28552
rect 17034 28500 17040 28552
rect 17092 28540 17098 28552
rect 17862 28540 17868 28552
rect 17092 28512 17868 28540
rect 17092 28500 17098 28512
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 19518 28540 19524 28552
rect 18340 28512 19524 28540
rect 18340 28484 18368 28512
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28509 19671 28543
rect 19720 28540 19748 28580
rect 20640 28580 24716 28608
rect 19869 28543 19927 28549
rect 19869 28540 19881 28543
rect 19720 28512 19881 28540
rect 19613 28503 19671 28509
rect 19869 28509 19881 28512
rect 19915 28509 19927 28543
rect 19869 28503 19927 28509
rect 18230 28472 18236 28484
rect 14783 28444 15516 28472
rect 15580 28444 18236 28472
rect 14783 28441 14795 28444
rect 14737 28435 14795 28441
rect 12713 28407 12771 28413
rect 12713 28404 12725 28407
rect 12676 28376 12725 28404
rect 12676 28364 12682 28376
rect 12713 28373 12725 28376
rect 12759 28404 12771 28407
rect 13541 28407 13599 28413
rect 13541 28404 13553 28407
rect 12759 28376 13553 28404
rect 12759 28373 12771 28376
rect 12713 28367 12771 28373
rect 13541 28373 13553 28376
rect 13587 28373 13599 28407
rect 13541 28367 13599 28373
rect 13722 28364 13728 28416
rect 13780 28404 13786 28416
rect 14826 28404 14832 28416
rect 13780 28376 14832 28404
rect 13780 28364 13786 28376
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 15488 28404 15516 28444
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 18322 28432 18328 28484
rect 18380 28432 18386 28484
rect 18417 28475 18475 28481
rect 18417 28441 18429 28475
rect 18463 28441 18475 28475
rect 19628 28472 19656 28503
rect 20346 28500 20352 28552
rect 20404 28540 20410 28552
rect 20640 28540 20668 28580
rect 20404 28512 20668 28540
rect 20404 28500 20410 28512
rect 21266 28500 21272 28552
rect 21324 28540 21330 28552
rect 21637 28543 21695 28549
rect 21637 28540 21649 28543
rect 21324 28512 21649 28540
rect 21324 28500 21330 28512
rect 21637 28509 21649 28512
rect 21683 28509 21695 28543
rect 21637 28503 21695 28509
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 19702 28472 19708 28484
rect 19628 28444 19708 28472
rect 18417 28435 18475 28441
rect 18432 28404 18460 28435
rect 19702 28432 19708 28444
rect 19760 28432 19766 28484
rect 22094 28472 22100 28484
rect 20456 28444 22100 28472
rect 18690 28404 18696 28416
rect 15488 28376 18696 28404
rect 18690 28364 18696 28376
rect 18748 28364 18754 28416
rect 18877 28407 18935 28413
rect 18877 28373 18889 28407
rect 18923 28404 18935 28407
rect 20456 28404 20484 28444
rect 22094 28432 22100 28444
rect 22152 28432 22158 28484
rect 22940 28472 22968 28503
rect 23658 28500 23664 28552
rect 23716 28540 23722 28552
rect 24578 28540 24584 28552
rect 23716 28512 24584 28540
rect 23716 28500 23722 28512
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 24688 28540 24716 28580
rect 25590 28568 25596 28620
rect 25648 28608 25654 28620
rect 26881 28611 26939 28617
rect 26881 28608 26893 28611
rect 25648 28580 26893 28608
rect 25648 28568 25654 28580
rect 26881 28577 26893 28580
rect 26927 28577 26939 28611
rect 26881 28571 26939 28577
rect 24837 28543 24895 28549
rect 24837 28540 24849 28543
rect 24688 28512 24849 28540
rect 24837 28509 24849 28512
rect 24883 28509 24895 28543
rect 24837 28503 24895 28509
rect 25774 28500 25780 28552
rect 25832 28540 25838 28552
rect 25832 28512 26004 28540
rect 25832 28500 25838 28512
rect 25866 28472 25872 28484
rect 22940 28444 25872 28472
rect 25866 28432 25872 28444
rect 25924 28432 25930 28484
rect 25976 28472 26004 28512
rect 27126 28475 27184 28481
rect 27126 28472 27138 28475
rect 25976 28444 27138 28472
rect 27126 28441 27138 28444
rect 27172 28441 27184 28475
rect 27126 28435 27184 28441
rect 18923 28376 20484 28404
rect 18923 28373 18935 28376
rect 18877 28367 18935 28373
rect 20622 28364 20628 28416
rect 20680 28404 20686 28416
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20680 28376 21005 28404
rect 20680 28364 20686 28376
rect 20993 28373 21005 28376
rect 21039 28373 21051 28407
rect 20993 28367 21051 28373
rect 25038 28364 25044 28416
rect 25096 28404 25102 28416
rect 28261 28407 28319 28413
rect 28261 28404 28273 28407
rect 25096 28376 28273 28404
rect 25096 28364 25102 28376
rect 28261 28373 28273 28376
rect 28307 28373 28319 28407
rect 28261 28367 28319 28373
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 2314 28200 2320 28212
rect 1780 28172 2320 28200
rect 1780 28076 1808 28172
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 3142 28160 3148 28212
rect 3200 28200 3206 28212
rect 4985 28203 5043 28209
rect 3200 28172 4016 28200
rect 3200 28160 3206 28172
rect 3878 28132 3884 28144
rect 1872 28104 3884 28132
rect 1762 28024 1768 28076
rect 1820 28024 1826 28076
rect 1872 28073 1900 28104
rect 3878 28092 3884 28104
rect 3936 28092 3942 28144
rect 3988 28132 4016 28172
rect 4985 28169 4997 28203
rect 5031 28200 5043 28203
rect 5166 28200 5172 28212
rect 5031 28172 5172 28200
rect 5031 28169 5043 28172
rect 4985 28163 5043 28169
rect 5166 28160 5172 28172
rect 5224 28160 5230 28212
rect 7190 28160 7196 28212
rect 7248 28160 7254 28212
rect 7374 28160 7380 28212
rect 7432 28200 7438 28212
rect 8113 28203 8171 28209
rect 8113 28200 8125 28203
rect 7432 28172 8125 28200
rect 7432 28160 7438 28172
rect 8113 28169 8125 28172
rect 8159 28169 8171 28203
rect 8113 28163 8171 28169
rect 9122 28160 9128 28212
rect 9180 28160 9186 28212
rect 11882 28160 11888 28212
rect 11940 28160 11946 28212
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 14461 28203 14519 28209
rect 14461 28200 14473 28203
rect 14240 28172 14473 28200
rect 14240 28160 14246 28172
rect 14461 28169 14473 28172
rect 14507 28169 14519 28203
rect 14461 28163 14519 28169
rect 15746 28160 15752 28212
rect 15804 28200 15810 28212
rect 16206 28200 16212 28212
rect 15804 28172 16212 28200
rect 15804 28160 15810 28172
rect 16206 28160 16212 28172
rect 16264 28200 16270 28212
rect 16301 28203 16359 28209
rect 16301 28200 16313 28203
rect 16264 28172 16313 28200
rect 16264 28160 16270 28172
rect 16301 28169 16313 28172
rect 16347 28169 16359 28203
rect 18966 28200 18972 28212
rect 16301 28163 16359 28169
rect 18708 28172 18972 28200
rect 8205 28135 8263 28141
rect 3988 28104 7880 28132
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28033 1915 28067
rect 1857 28027 1915 28033
rect 1946 28024 1952 28076
rect 2004 28064 2010 28076
rect 2593 28067 2651 28073
rect 2593 28064 2605 28067
rect 2004 28036 2605 28064
rect 2004 28024 2010 28036
rect 2593 28033 2605 28036
rect 2639 28033 2651 28067
rect 2593 28027 2651 28033
rect 2860 28067 2918 28073
rect 2860 28033 2872 28067
rect 2906 28064 2918 28067
rect 4062 28064 4068 28076
rect 2906 28036 4068 28064
rect 2906 28033 2918 28036
rect 2860 28027 2918 28033
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28064 5043 28067
rect 5166 28064 5172 28076
rect 5031 28036 5172 28064
rect 5031 28033 5043 28036
rect 4985 28027 5043 28033
rect 5166 28024 5172 28036
rect 5224 28024 5230 28076
rect 5629 28067 5687 28073
rect 5629 28064 5641 28067
rect 5368 28036 5641 28064
rect 2038 27956 2044 28008
rect 2096 27956 2102 28008
rect 4617 27999 4675 28005
rect 4617 27965 4629 27999
rect 4663 27996 4675 27999
rect 5258 27996 5264 28008
rect 4663 27968 5264 27996
rect 4663 27965 4675 27968
rect 4617 27959 4675 27965
rect 5258 27956 5264 27968
rect 5316 27956 5322 28008
rect 3694 27888 3700 27940
rect 3752 27928 3758 27940
rect 5368 27928 5396 28036
rect 5629 28033 5641 28036
rect 5675 28033 5687 28067
rect 5629 28027 5687 28033
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 6822 28064 6828 28076
rect 5776 28036 6828 28064
rect 5776 28024 5782 28036
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 7006 28024 7012 28076
rect 7064 28064 7070 28076
rect 7374 28064 7380 28076
rect 7064 28036 7380 28064
rect 7064 28024 7070 28036
rect 7374 28024 7380 28036
rect 7432 28024 7438 28076
rect 7852 28073 7880 28104
rect 8205 28101 8217 28135
rect 8251 28132 8263 28135
rect 8478 28132 8484 28144
rect 8251 28104 8484 28132
rect 8251 28101 8263 28104
rect 8205 28095 8263 28101
rect 8478 28092 8484 28104
rect 8536 28092 8542 28144
rect 11698 28132 11704 28144
rect 9048 28104 11704 28132
rect 7837 28067 7895 28073
rect 7837 28033 7849 28067
rect 7883 28033 7895 28067
rect 7837 28027 7895 28033
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28033 8355 28067
rect 8297 28027 8355 28033
rect 5445 27999 5503 28005
rect 5445 27965 5457 27999
rect 5491 27996 5503 27999
rect 5736 27996 5764 28024
rect 5491 27968 5764 27996
rect 5491 27965 5503 27968
rect 5445 27959 5503 27965
rect 5994 27956 6000 28008
rect 6052 27956 6058 28008
rect 6733 27999 6791 28005
rect 6733 27965 6745 27999
rect 6779 27965 6791 27999
rect 6840 27996 6868 28024
rect 7466 27996 7472 28008
rect 6840 27968 7472 27996
rect 6733 27959 6791 27965
rect 3752 27900 5396 27928
rect 3752 27888 3758 27900
rect 5902 27888 5908 27940
rect 5960 27888 5966 27940
rect 6748 27928 6776 27959
rect 7466 27956 7472 27968
rect 7524 27996 7530 28008
rect 8312 27996 8340 28027
rect 7524 27968 8340 27996
rect 7524 27956 7530 27968
rect 8754 27956 8760 28008
rect 8812 27956 8818 28008
rect 7006 27928 7012 27940
rect 6748 27900 7012 27928
rect 7006 27888 7012 27900
rect 7064 27888 7070 27940
rect 7101 27931 7159 27937
rect 7101 27897 7113 27931
rect 7147 27928 7159 27931
rect 9048 27928 9076 28104
rect 11698 28092 11704 28104
rect 11756 28092 11762 28144
rect 11793 28135 11851 28141
rect 11793 28101 11805 28135
rect 11839 28132 11851 28135
rect 14366 28132 14372 28144
rect 11839 28104 14372 28132
rect 11839 28101 11851 28104
rect 11793 28095 11851 28101
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 12452 28073 12480 28104
rect 14366 28092 14372 28104
rect 14424 28092 14430 28144
rect 17402 28132 17408 28144
rect 16684 28104 17408 28132
rect 9841 28067 9899 28073
rect 9841 28064 9853 28067
rect 9272 28036 9853 28064
rect 9272 28024 9278 28036
rect 9841 28033 9853 28036
rect 9887 28033 9899 28067
rect 9841 28027 9899 28033
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28064 12495 28067
rect 12483 28036 12517 28064
rect 12483 28033 12495 28036
rect 12437 28027 12495 28033
rect 14090 28024 14096 28076
rect 14148 28024 14154 28076
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28064 14335 28067
rect 14323 28036 14412 28064
rect 14323 28033 14335 28036
rect 14277 28027 14335 28033
rect 14384 28008 14412 28036
rect 14458 28024 14464 28076
rect 14516 28064 14522 28076
rect 14921 28067 14979 28073
rect 14921 28064 14933 28067
rect 14516 28036 14933 28064
rect 14516 28024 14522 28036
rect 14921 28033 14933 28036
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 15102 28024 15108 28076
rect 15160 28024 15166 28076
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28064 15347 28067
rect 16684 28064 16712 28104
rect 17402 28092 17408 28104
rect 17460 28132 17466 28144
rect 18506 28132 18512 28144
rect 17460 28104 18512 28132
rect 17460 28092 17466 28104
rect 18506 28092 18512 28104
rect 18564 28092 18570 28144
rect 15335 28036 16712 28064
rect 15335 28033 15347 28036
rect 15289 28027 15347 28033
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 18708 28073 18736 28172
rect 18966 28160 18972 28172
rect 19024 28200 19030 28212
rect 19024 28172 19334 28200
rect 19024 28160 19030 28172
rect 19306 28132 19334 28172
rect 19978 28160 19984 28212
rect 20036 28200 20042 28212
rect 20622 28200 20628 28212
rect 20036 28172 20628 28200
rect 20036 28160 20042 28172
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 21450 28160 21456 28212
rect 21508 28200 21514 28212
rect 24670 28200 24676 28212
rect 21508 28172 24676 28200
rect 21508 28160 21514 28172
rect 24670 28160 24676 28172
rect 24728 28160 24734 28212
rect 24762 28160 24768 28212
rect 24820 28160 24826 28212
rect 25130 28160 25136 28212
rect 25188 28200 25194 28212
rect 25409 28203 25467 28209
rect 25409 28200 25421 28203
rect 25188 28172 25421 28200
rect 25188 28160 25194 28172
rect 25409 28169 25421 28172
rect 25455 28169 25467 28203
rect 25409 28163 25467 28169
rect 26050 28160 26056 28212
rect 26108 28200 26114 28212
rect 26145 28203 26203 28209
rect 26145 28200 26157 28203
rect 26108 28172 26157 28200
rect 26108 28160 26114 28172
rect 26145 28169 26157 28172
rect 26191 28169 26203 28203
rect 26145 28163 26203 28169
rect 26326 28160 26332 28212
rect 26384 28200 26390 28212
rect 27939 28203 27997 28209
rect 27939 28200 27951 28203
rect 26384 28172 27951 28200
rect 26384 28160 26390 28172
rect 27939 28169 27951 28172
rect 27985 28169 27997 28203
rect 27939 28163 27997 28169
rect 22370 28132 22376 28144
rect 19306 28104 22376 28132
rect 22370 28092 22376 28104
rect 22428 28092 22434 28144
rect 17109 28067 17167 28073
rect 17109 28064 17121 28067
rect 16816 28036 17121 28064
rect 16816 28024 16822 28036
rect 17109 28033 17121 28036
rect 17155 28033 17167 28067
rect 17109 28027 17167 28033
rect 18693 28067 18751 28073
rect 18693 28033 18705 28067
rect 18739 28033 18751 28067
rect 18693 28027 18751 28033
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 18969 28067 19027 28073
rect 18969 28033 18981 28067
rect 19015 28033 19027 28067
rect 18969 28027 19027 28033
rect 9585 27999 9643 28005
rect 9585 27965 9597 27999
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 7147 27900 9076 27928
rect 9125 27931 9183 27937
rect 7147 27897 7159 27900
rect 7101 27891 7159 27897
rect 9125 27897 9137 27931
rect 9171 27897 9183 27931
rect 9125 27891 9183 27897
rect 3973 27863 4031 27869
rect 3973 27829 3985 27863
rect 4019 27860 4031 27863
rect 7190 27860 7196 27872
rect 4019 27832 7196 27860
rect 4019 27829 4031 27832
rect 3973 27823 4031 27829
rect 7190 27820 7196 27832
rect 7248 27820 7254 27872
rect 9030 27820 9036 27872
rect 9088 27860 9094 27872
rect 9140 27860 9168 27891
rect 9088 27832 9168 27860
rect 9600 27860 9628 27959
rect 10962 27956 10968 28008
rect 11020 27996 11026 28008
rect 11238 27996 11244 28008
rect 11020 27968 11244 27996
rect 11020 27956 11026 27968
rect 11238 27956 11244 27968
rect 11296 27956 11302 28008
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27965 12771 27999
rect 12713 27959 12771 27965
rect 12728 27928 12756 27959
rect 14366 27956 14372 28008
rect 14424 27956 14430 28008
rect 15470 27996 15476 28008
rect 14476 27968 15476 27996
rect 13262 27928 13268 27940
rect 12728 27900 13268 27928
rect 13262 27888 13268 27900
rect 13320 27928 13326 27940
rect 14476 27928 14504 27968
rect 15470 27956 15476 27968
rect 15528 27996 15534 28008
rect 15933 27999 15991 28005
rect 15933 27996 15945 27999
rect 15528 27968 15945 27996
rect 15528 27956 15534 27968
rect 15933 27965 15945 27968
rect 15979 27965 15991 27999
rect 15933 27959 15991 27965
rect 16206 27956 16212 28008
rect 16264 27996 16270 28008
rect 16301 27999 16359 28005
rect 16301 27996 16313 27999
rect 16264 27968 16313 27996
rect 16264 27956 16270 27968
rect 16301 27965 16313 27968
rect 16347 27965 16359 27999
rect 16301 27959 16359 27965
rect 16853 27999 16911 28005
rect 16853 27965 16865 27999
rect 16899 27965 16911 27999
rect 16853 27959 16911 27965
rect 13320 27900 14504 27928
rect 13320 27888 13326 27900
rect 15102 27888 15108 27940
rect 15160 27928 15166 27940
rect 15160 27900 15792 27928
rect 15160 27888 15166 27900
rect 9766 27860 9772 27872
rect 9600 27832 9772 27860
rect 9088 27820 9094 27832
rect 9766 27820 9772 27832
rect 9824 27820 9830 27872
rect 9950 27820 9956 27872
rect 10008 27860 10014 27872
rect 10965 27863 11023 27869
rect 10965 27860 10977 27863
rect 10008 27832 10977 27860
rect 10008 27820 10014 27832
rect 10965 27829 10977 27832
rect 11011 27829 11023 27863
rect 10965 27823 11023 27829
rect 15473 27863 15531 27869
rect 15473 27829 15485 27863
rect 15519 27860 15531 27863
rect 15654 27860 15660 27872
rect 15519 27832 15660 27860
rect 15519 27829 15531 27832
rect 15473 27823 15531 27829
rect 15654 27820 15660 27832
rect 15712 27820 15718 27872
rect 15764 27860 15792 27900
rect 16022 27888 16028 27940
rect 16080 27928 16086 27940
rect 16482 27928 16488 27940
rect 16080 27900 16488 27928
rect 16080 27888 16086 27900
rect 16482 27888 16488 27900
rect 16540 27928 16546 27940
rect 16868 27928 16896 27959
rect 16540 27900 16896 27928
rect 18233 27931 18291 27937
rect 16540 27888 16546 27900
rect 18233 27897 18245 27931
rect 18279 27928 18291 27931
rect 18322 27928 18328 27940
rect 18279 27900 18328 27928
rect 18279 27897 18291 27900
rect 18233 27891 18291 27897
rect 18322 27888 18328 27900
rect 18380 27888 18386 27940
rect 17586 27860 17592 27872
rect 15764 27832 17592 27860
rect 17586 27820 17592 27832
rect 17644 27860 17650 27872
rect 18892 27860 18920 28027
rect 18984 27928 19012 28027
rect 19058 28024 19064 28076
rect 19116 28024 19122 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 20329 28067 20387 28073
rect 20329 28064 20341 28067
rect 19484 28036 20341 28064
rect 19484 28024 19490 28036
rect 20329 28033 20341 28036
rect 20375 28033 20387 28067
rect 20329 28027 20387 28033
rect 20622 28024 20628 28076
rect 20680 28064 20686 28076
rect 22537 28067 22595 28073
rect 22537 28064 22549 28067
rect 20680 28036 22549 28064
rect 20680 28024 20686 28036
rect 22537 28033 22549 28036
rect 22583 28033 22595 28067
rect 22537 28027 22595 28033
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28064 24363 28067
rect 24854 28064 24860 28076
rect 24351 28036 24860 28064
rect 24351 28033 24363 28036
rect 24305 28027 24363 28033
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 24949 28067 25007 28073
rect 24949 28033 24961 28067
rect 24995 28064 25007 28067
rect 25130 28064 25136 28076
rect 24995 28036 25136 28064
rect 24995 28033 25007 28036
rect 24949 28027 25007 28033
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 25590 28024 25596 28076
rect 25648 28024 25654 28076
rect 26050 28024 26056 28076
rect 26108 28024 26114 28076
rect 26418 28024 26424 28076
rect 26476 28064 26482 28076
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 26476 28036 27169 28064
rect 26476 28024 26482 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 27836 28067 27894 28073
rect 27836 28064 27848 28067
rect 27672 28036 27848 28064
rect 27672 28024 27678 28036
rect 27836 28033 27848 28036
rect 27882 28033 27894 28067
rect 27836 28027 27894 28033
rect 19242 27956 19248 28008
rect 19300 27956 19306 28008
rect 19518 27956 19524 28008
rect 19576 27996 19582 28008
rect 19794 27996 19800 28008
rect 19576 27968 19800 27996
rect 19576 27956 19582 27968
rect 19794 27956 19800 27968
rect 19852 27996 19858 28008
rect 20073 27999 20131 28005
rect 20073 27996 20085 27999
rect 19852 27968 20085 27996
rect 19852 27956 19858 27968
rect 20073 27965 20085 27968
rect 20119 27965 20131 27999
rect 20073 27959 20131 27965
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27965 22339 27999
rect 22281 27959 22339 27965
rect 19260 27928 19288 27956
rect 18984 27900 19288 27928
rect 17644 27832 18920 27860
rect 17644 27820 17650 27832
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 19245 27863 19303 27869
rect 19245 27860 19257 27863
rect 19116 27832 19257 27860
rect 19116 27820 19122 27832
rect 19245 27829 19257 27832
rect 19291 27829 19303 27863
rect 19245 27823 19303 27829
rect 19886 27820 19892 27872
rect 19944 27860 19950 27872
rect 21453 27863 21511 27869
rect 21453 27860 21465 27863
rect 19944 27832 21465 27860
rect 19944 27820 19950 27832
rect 21453 27829 21465 27832
rect 21499 27829 21511 27863
rect 22296 27860 22324 27959
rect 22646 27860 22652 27872
rect 22296 27832 22652 27860
rect 21453 27823 21511 27829
rect 22646 27820 22652 27832
rect 22704 27820 22710 27872
rect 23661 27863 23719 27869
rect 23661 27829 23673 27863
rect 23707 27860 23719 27863
rect 24026 27860 24032 27872
rect 23707 27832 24032 27860
rect 23707 27829 23719 27832
rect 23661 27823 23719 27829
rect 24026 27820 24032 27832
rect 24084 27820 24090 27872
rect 24118 27820 24124 27872
rect 24176 27860 24182 27872
rect 27341 27863 27399 27869
rect 27341 27860 27353 27863
rect 24176 27832 27353 27860
rect 24176 27820 24182 27832
rect 27341 27829 27353 27832
rect 27387 27829 27399 27863
rect 27341 27823 27399 27829
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 474 27616 480 27668
rect 532 27656 538 27668
rect 3602 27656 3608 27668
rect 532 27628 3608 27656
rect 532 27616 538 27628
rect 3602 27616 3608 27628
rect 3660 27616 3666 27668
rect 9766 27616 9772 27668
rect 9824 27656 9830 27668
rect 10042 27656 10048 27668
rect 9824 27628 10048 27656
rect 9824 27616 9830 27628
rect 10042 27616 10048 27628
rect 10100 27616 10106 27668
rect 11698 27616 11704 27668
rect 11756 27656 11762 27668
rect 12066 27656 12072 27668
rect 11756 27628 12072 27656
rect 11756 27616 11762 27628
rect 12066 27616 12072 27628
rect 12124 27656 12130 27668
rect 13814 27656 13820 27668
rect 12124 27628 13820 27656
rect 12124 27616 12130 27628
rect 13814 27616 13820 27628
rect 13872 27616 13878 27668
rect 14366 27616 14372 27668
rect 14424 27656 14430 27668
rect 18046 27656 18052 27668
rect 14424 27628 18052 27656
rect 14424 27616 14430 27628
rect 18046 27616 18052 27628
rect 18104 27616 18110 27668
rect 18340 27628 19380 27656
rect 3970 27548 3976 27600
rect 4028 27548 4034 27600
rect 4062 27548 4068 27600
rect 4120 27548 4126 27600
rect 5166 27548 5172 27600
rect 5224 27588 5230 27600
rect 5629 27591 5687 27597
rect 5629 27588 5641 27591
rect 5224 27560 5641 27588
rect 5224 27548 5230 27560
rect 5629 27557 5641 27560
rect 5675 27588 5687 27591
rect 5718 27588 5724 27600
rect 5675 27560 5724 27588
rect 5675 27557 5687 27560
rect 5629 27551 5687 27557
rect 5718 27548 5724 27560
rect 5776 27588 5782 27600
rect 7285 27591 7343 27597
rect 7285 27588 7297 27591
rect 5776 27560 7297 27588
rect 5776 27548 5782 27560
rect 7285 27557 7297 27560
rect 7331 27588 7343 27591
rect 7466 27588 7472 27600
rect 7331 27560 7472 27588
rect 7331 27557 7343 27560
rect 7285 27551 7343 27557
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 7760 27560 10456 27588
rect 3988 27520 4016 27548
rect 6457 27523 6515 27529
rect 6457 27520 6469 27523
rect 3988 27492 6469 27520
rect 6457 27489 6469 27492
rect 6503 27489 6515 27523
rect 6457 27483 6515 27489
rect 6914 27480 6920 27532
rect 6972 27520 6978 27532
rect 7760 27529 7788 27560
rect 7745 27523 7803 27529
rect 6972 27492 7328 27520
rect 6972 27480 6978 27492
rect 1946 27412 1952 27464
rect 2004 27452 2010 27464
rect 2041 27455 2099 27461
rect 2041 27452 2053 27455
rect 2004 27424 2053 27452
rect 2004 27412 2010 27424
rect 2041 27421 2053 27424
rect 2087 27421 2099 27455
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 2041 27415 2099 27421
rect 2240 27424 3985 27452
rect 1762 27344 1768 27396
rect 1820 27384 1826 27396
rect 2240 27384 2268 27424
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 4246 27412 4252 27464
rect 4304 27412 4310 27464
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27421 4583 27455
rect 4525 27415 4583 27421
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 4982 27452 4988 27464
rect 4847 27424 4988 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 1820 27356 2268 27384
rect 2308 27387 2366 27393
rect 1820 27344 1826 27356
rect 2308 27353 2320 27387
rect 2354 27384 2366 27387
rect 2406 27384 2412 27396
rect 2354 27356 2412 27384
rect 2354 27353 2366 27356
rect 2308 27347 2366 27353
rect 2406 27344 2412 27356
rect 2464 27344 2470 27396
rect 4540 27384 4568 27415
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5258 27412 5264 27464
rect 5316 27452 5322 27464
rect 5534 27452 5540 27464
rect 5316 27424 5540 27452
rect 5316 27412 5322 27424
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 5626 27412 5632 27464
rect 5684 27452 5690 27464
rect 5994 27452 6000 27464
rect 5684 27424 6000 27452
rect 5684 27412 5690 27424
rect 5994 27412 6000 27424
rect 6052 27452 6058 27464
rect 6089 27455 6147 27461
rect 6089 27452 6101 27455
rect 6052 27424 6101 27452
rect 6052 27412 6058 27424
rect 6089 27421 6101 27424
rect 6135 27421 6147 27455
rect 6089 27415 6147 27421
rect 4890 27384 4896 27396
rect 4540 27356 4896 27384
rect 4890 27344 4896 27356
rect 4948 27344 4954 27396
rect 6104 27384 6132 27415
rect 6270 27412 6276 27464
rect 6328 27412 6334 27464
rect 7300 27452 7328 27492
rect 7745 27489 7757 27523
rect 7791 27489 7803 27523
rect 7745 27483 7803 27489
rect 9585 27523 9643 27529
rect 9585 27489 9597 27523
rect 9631 27520 9643 27523
rect 9858 27520 9864 27532
rect 9631 27492 9864 27520
rect 9631 27489 9643 27492
rect 9585 27483 9643 27489
rect 9858 27480 9864 27492
rect 9916 27480 9922 27532
rect 10428 27520 10456 27560
rect 12618 27548 12624 27600
rect 12676 27588 12682 27600
rect 12713 27591 12771 27597
rect 12713 27588 12725 27591
rect 12676 27560 12725 27588
rect 12676 27548 12682 27560
rect 12713 27557 12725 27560
rect 12759 27557 12771 27591
rect 12713 27551 12771 27557
rect 14921 27591 14979 27597
rect 14921 27557 14933 27591
rect 14967 27588 14979 27591
rect 15286 27588 15292 27600
rect 14967 27560 15292 27588
rect 14967 27557 14979 27560
rect 14921 27551 14979 27557
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 18340 27588 18368 27628
rect 15396 27560 18368 27588
rect 18417 27591 18475 27597
rect 15396 27520 15424 27560
rect 18417 27557 18429 27591
rect 18463 27588 18475 27591
rect 19242 27588 19248 27600
rect 18463 27560 19248 27588
rect 18463 27557 18475 27560
rect 18417 27551 18475 27557
rect 19242 27548 19248 27560
rect 19300 27548 19306 27600
rect 19352 27588 19380 27628
rect 19996 27628 20852 27656
rect 19996 27588 20024 27628
rect 19352 27560 20024 27588
rect 20073 27591 20131 27597
rect 20073 27557 20085 27591
rect 20119 27588 20131 27591
rect 20714 27588 20720 27600
rect 20119 27560 20720 27588
rect 20119 27557 20131 27560
rect 20073 27551 20131 27557
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 20824 27588 20852 27628
rect 20898 27616 20904 27668
rect 20956 27656 20962 27668
rect 26234 27656 26240 27668
rect 20956 27628 26240 27656
rect 20956 27616 20962 27628
rect 26234 27616 26240 27628
rect 26292 27616 26298 27668
rect 21542 27588 21548 27600
rect 20824 27560 21548 27588
rect 21542 27548 21548 27560
rect 21600 27588 21606 27600
rect 22002 27588 22008 27600
rect 21600 27560 22008 27588
rect 21600 27548 21606 27560
rect 22002 27548 22008 27560
rect 22060 27548 22066 27600
rect 10428 27492 10548 27520
rect 8021 27455 8079 27461
rect 8021 27452 8033 27455
rect 7300 27424 8033 27452
rect 8021 27421 8033 27424
rect 8067 27421 8079 27455
rect 8021 27415 8079 27421
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9953 27455 10011 27461
rect 9953 27452 9965 27455
rect 9180 27424 9965 27452
rect 9180 27412 9186 27424
rect 7006 27384 7012 27396
rect 6104 27356 7012 27384
rect 7006 27344 7012 27356
rect 7064 27344 7070 27396
rect 3326 27276 3332 27328
rect 3384 27316 3390 27328
rect 3421 27319 3479 27325
rect 3421 27316 3433 27319
rect 3384 27288 3433 27316
rect 3384 27276 3390 27288
rect 3421 27285 3433 27288
rect 3467 27285 3479 27319
rect 3421 27279 3479 27285
rect 5629 27319 5687 27325
rect 5629 27285 5641 27319
rect 5675 27316 5687 27319
rect 5718 27316 5724 27328
rect 5675 27288 5724 27316
rect 5675 27285 5687 27288
rect 5629 27279 5687 27285
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 6362 27276 6368 27328
rect 6420 27316 6426 27328
rect 6638 27316 6644 27328
rect 6420 27288 6644 27316
rect 6420 27276 6426 27288
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 7285 27319 7343 27325
rect 7285 27285 7297 27319
rect 7331 27316 7343 27319
rect 7466 27316 7472 27328
rect 7331 27288 7472 27316
rect 7331 27285 7343 27288
rect 7285 27279 7343 27285
rect 7466 27276 7472 27288
rect 7524 27276 7530 27328
rect 8386 27276 8392 27328
rect 8444 27316 8450 27328
rect 9214 27316 9220 27328
rect 8444 27288 9220 27316
rect 8444 27276 8450 27288
rect 9214 27276 9220 27288
rect 9272 27276 9278 27328
rect 9508 27316 9536 27424
rect 9953 27421 9965 27424
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10042 27412 10048 27464
rect 10100 27452 10106 27464
rect 10413 27455 10471 27461
rect 10413 27452 10425 27455
rect 10100 27424 10425 27452
rect 10100 27412 10106 27424
rect 10413 27421 10425 27424
rect 10459 27421 10471 27455
rect 10520 27452 10548 27492
rect 11440 27492 15424 27520
rect 11238 27452 11244 27464
rect 10520 27424 11244 27452
rect 10413 27415 10471 27421
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 10658 27387 10716 27393
rect 10658 27384 10670 27387
rect 9640 27356 10670 27384
rect 9640 27344 9646 27356
rect 10658 27353 10670 27356
rect 10704 27353 10716 27387
rect 10658 27347 10716 27353
rect 10778 27344 10784 27396
rect 10836 27384 10842 27396
rect 11440 27384 11468 27492
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 17129 27523 17187 27529
rect 15804 27492 16528 27520
rect 15804 27480 15810 27492
rect 12342 27412 12348 27464
rect 12400 27412 12406 27464
rect 12618 27412 12624 27464
rect 12676 27412 12682 27464
rect 13170 27412 13176 27464
rect 13228 27412 13234 27464
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27421 13599 27455
rect 13541 27415 13599 27421
rect 10836 27356 11468 27384
rect 10836 27344 10842 27356
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 9508 27288 9965 27316
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 11698 27276 11704 27328
rect 11756 27316 11762 27328
rect 11793 27319 11851 27325
rect 11793 27316 11805 27319
rect 11756 27288 11805 27316
rect 11756 27276 11762 27288
rect 11793 27285 11805 27288
rect 11839 27285 11851 27319
rect 12636 27316 12664 27412
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 12636 27288 12725 27316
rect 11793 27279 11851 27285
rect 12713 27285 12725 27288
rect 12759 27316 12771 27319
rect 12802 27316 12808 27328
rect 12759 27288 12808 27316
rect 12759 27285 12771 27288
rect 12713 27279 12771 27285
rect 12802 27276 12808 27288
rect 12860 27316 12866 27328
rect 13556 27325 13584 27415
rect 13906 27412 13912 27464
rect 13964 27452 13970 27464
rect 14366 27452 14372 27464
rect 13964 27424 14372 27452
rect 13964 27412 13970 27424
rect 14366 27412 14372 27424
rect 14424 27452 14430 27464
rect 14737 27455 14795 27461
rect 14737 27452 14749 27455
rect 14424 27424 14749 27452
rect 14424 27412 14430 27424
rect 14737 27421 14749 27424
rect 14783 27421 14795 27455
rect 14737 27415 14795 27421
rect 15381 27455 15439 27461
rect 15381 27421 15393 27455
rect 15427 27452 15439 27455
rect 15470 27452 15476 27464
rect 15427 27424 15476 27452
rect 15427 27421 15439 27424
rect 15381 27415 15439 27421
rect 15470 27412 15476 27424
rect 15528 27412 15534 27464
rect 16393 27455 16451 27461
rect 16393 27421 16405 27455
rect 16439 27421 16451 27455
rect 16500 27452 16528 27492
rect 17129 27489 17141 27523
rect 17175 27520 17187 27523
rect 19613 27523 19671 27529
rect 19613 27520 19625 27523
rect 17175 27492 19625 27520
rect 17175 27489 17187 27492
rect 17129 27483 17187 27489
rect 19613 27489 19625 27492
rect 19659 27489 19671 27523
rect 19613 27483 19671 27489
rect 20162 27480 20168 27532
rect 20220 27520 20226 27532
rect 20220 27492 22784 27520
rect 20220 27480 20226 27492
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 16500 27424 17509 27452
rect 16393 27415 16451 27421
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 14550 27344 14556 27396
rect 14608 27344 14614 27396
rect 15194 27344 15200 27396
rect 15252 27384 15258 27396
rect 16408 27384 16436 27415
rect 15252 27356 16436 27384
rect 15252 27344 15258 27356
rect 13541 27319 13599 27325
rect 13541 27316 13553 27319
rect 12860 27288 13553 27316
rect 12860 27276 12866 27288
rect 13541 27285 13553 27288
rect 13587 27285 13599 27319
rect 13541 27279 13599 27285
rect 15746 27276 15752 27328
rect 15804 27276 15810 27328
rect 16209 27319 16267 27325
rect 16209 27285 16221 27319
rect 16255 27316 16267 27319
rect 17310 27316 17316 27328
rect 16255 27288 17316 27316
rect 16255 27285 16267 27288
rect 16209 27279 16267 27285
rect 17310 27276 17316 27288
rect 17368 27276 17374 27328
rect 17512 27325 17540 27415
rect 17862 27412 17868 27464
rect 17920 27452 17926 27464
rect 18049 27455 18107 27461
rect 18049 27452 18061 27455
rect 17920 27424 18061 27452
rect 17920 27412 17926 27424
rect 18049 27421 18061 27424
rect 18095 27421 18107 27455
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 18049 27415 18107 27421
rect 18340 27424 20269 27452
rect 17497 27319 17555 27325
rect 17497 27285 17509 27319
rect 17543 27285 17555 27319
rect 18340 27316 18368 27424
rect 20257 27421 20269 27424
rect 20303 27421 20315 27455
rect 20806 27452 20812 27464
rect 20257 27415 20315 27421
rect 20640 27424 20812 27452
rect 18414 27344 18420 27396
rect 18472 27384 18478 27396
rect 20640 27384 20668 27424
rect 20806 27412 20812 27424
rect 20864 27412 20870 27464
rect 20898 27412 20904 27464
rect 20956 27412 20962 27464
rect 21358 27412 21364 27464
rect 21416 27412 21422 27464
rect 22002 27412 22008 27464
rect 22060 27412 22066 27464
rect 22646 27412 22652 27464
rect 22704 27412 22710 27464
rect 22756 27452 22784 27492
rect 24581 27455 24639 27461
rect 22756 27424 23060 27452
rect 21634 27384 21640 27396
rect 18472 27356 20668 27384
rect 20732 27356 21640 27384
rect 18472 27344 18478 27356
rect 18509 27319 18567 27325
rect 18509 27316 18521 27319
rect 18340 27288 18521 27316
rect 17497 27279 17555 27285
rect 18509 27285 18521 27288
rect 18555 27285 18567 27319
rect 18509 27279 18567 27285
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 19610 27316 19616 27328
rect 19392 27288 19616 27316
rect 19392 27276 19398 27288
rect 19610 27276 19616 27288
rect 19668 27276 19674 27328
rect 20070 27276 20076 27328
rect 20128 27316 20134 27328
rect 20622 27316 20628 27328
rect 20128 27288 20628 27316
rect 20128 27276 20134 27288
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 20732 27325 20760 27356
rect 21634 27344 21640 27356
rect 21692 27344 21698 27396
rect 22370 27344 22376 27396
rect 22428 27384 22434 27396
rect 22894 27387 22952 27393
rect 22894 27384 22906 27387
rect 22428 27356 22906 27384
rect 22428 27344 22434 27356
rect 22894 27353 22906 27356
rect 22940 27353 22952 27387
rect 23032 27384 23060 27424
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 24670 27452 24676 27464
rect 24627 27424 24676 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 24670 27412 24676 27424
rect 24728 27452 24734 27464
rect 26973 27455 27031 27461
rect 26973 27452 26985 27455
rect 24728 27424 26985 27452
rect 24728 27412 24734 27424
rect 26973 27421 26985 27424
rect 27019 27421 27031 27455
rect 26973 27415 27031 27421
rect 24826 27387 24884 27393
rect 24826 27384 24838 27387
rect 23032 27356 24838 27384
rect 22894 27347 22952 27353
rect 24826 27353 24838 27356
rect 24872 27353 24884 27387
rect 27218 27387 27276 27393
rect 27218 27384 27230 27387
rect 24826 27347 24884 27353
rect 24964 27356 27230 27384
rect 20717 27319 20775 27325
rect 20717 27285 20729 27319
rect 20763 27285 20775 27319
rect 20717 27279 20775 27285
rect 21542 27276 21548 27328
rect 21600 27276 21606 27328
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22186 27316 22192 27328
rect 22143 27288 22192 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22186 27276 22192 27288
rect 22244 27276 22250 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 24029 27319 24087 27325
rect 24029 27316 24041 27319
rect 22336 27288 24041 27316
rect 22336 27276 22342 27288
rect 24029 27285 24041 27288
rect 24075 27285 24087 27319
rect 24029 27279 24087 27285
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 24964 27316 24992 27356
rect 27218 27353 27230 27356
rect 27264 27353 27276 27387
rect 27218 27347 27276 27353
rect 24176 27288 24992 27316
rect 24176 27276 24182 27288
rect 25130 27276 25136 27328
rect 25188 27316 25194 27328
rect 25961 27319 26019 27325
rect 25961 27316 25973 27319
rect 25188 27288 25973 27316
rect 25188 27276 25194 27288
rect 25961 27285 25973 27288
rect 26007 27285 26019 27319
rect 25961 27279 26019 27285
rect 27614 27276 27620 27328
rect 27672 27316 27678 27328
rect 28353 27319 28411 27325
rect 28353 27316 28365 27319
rect 27672 27288 28365 27316
rect 27672 27276 27678 27288
rect 28353 27285 28365 27288
rect 28399 27285 28411 27319
rect 28353 27279 28411 27285
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 2866 27072 2872 27124
rect 2924 27112 2930 27124
rect 2924 27084 8892 27112
rect 2924 27072 2930 27084
rect 2498 27004 2504 27056
rect 2556 27044 2562 27056
rect 2593 27047 2651 27053
rect 2593 27044 2605 27047
rect 2556 27016 2605 27044
rect 2556 27004 2562 27016
rect 2593 27013 2605 27016
rect 2639 27013 2651 27047
rect 2593 27007 2651 27013
rect 5000 27016 5856 27044
rect 5000 26988 5028 27016
rect 1762 26936 1768 26988
rect 1820 26936 1826 26988
rect 2041 26979 2099 26985
rect 2041 26945 2053 26979
rect 2087 26976 2099 26979
rect 2087 26948 2360 26976
rect 2087 26945 2099 26948
rect 2041 26939 2099 26945
rect 2130 26868 2136 26920
rect 2188 26868 2194 26920
rect 2332 26908 2360 26948
rect 4798 26936 4804 26988
rect 4856 26936 4862 26988
rect 4982 26936 4988 26988
rect 5040 26936 5046 26988
rect 5828 26985 5856 27016
rect 6086 27004 6092 27056
rect 6144 27044 6150 27056
rect 7929 27047 7987 27053
rect 7929 27044 7941 27047
rect 6144 27016 7941 27044
rect 6144 27004 6150 27016
rect 7929 27013 7941 27016
rect 7975 27013 7987 27047
rect 8864 27044 8892 27084
rect 9122 27072 9128 27124
rect 9180 27112 9186 27124
rect 9306 27112 9312 27124
rect 9180 27084 9312 27112
rect 9180 27072 9186 27084
rect 9306 27072 9312 27084
rect 9364 27072 9370 27124
rect 9769 27115 9827 27121
rect 9769 27081 9781 27115
rect 9815 27112 9827 27115
rect 10226 27112 10232 27124
rect 9815 27084 10232 27112
rect 9815 27081 9827 27084
rect 9769 27075 9827 27081
rect 10226 27072 10232 27084
rect 10284 27072 10290 27124
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27112 11023 27115
rect 12618 27112 12624 27124
rect 11011 27084 12624 27112
rect 11011 27081 11023 27084
rect 10965 27075 11023 27081
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 12713 27115 12771 27121
rect 12713 27081 12725 27115
rect 12759 27112 12771 27115
rect 12802 27112 12808 27124
rect 12759 27084 12808 27112
rect 12759 27081 12771 27084
rect 12713 27075 12771 27081
rect 12802 27072 12808 27084
rect 12860 27112 12866 27124
rect 13541 27115 13599 27121
rect 13541 27112 13553 27115
rect 12860 27084 13553 27112
rect 12860 27072 12866 27084
rect 13541 27081 13553 27084
rect 13587 27081 13599 27115
rect 13541 27075 13599 27081
rect 14090 27072 14096 27124
rect 14148 27112 14154 27124
rect 14550 27112 14556 27124
rect 14148 27084 14556 27112
rect 14148 27072 14154 27084
rect 14550 27072 14556 27084
rect 14608 27112 14614 27124
rect 15289 27115 15347 27121
rect 14608 27084 14964 27112
rect 14608 27072 14614 27084
rect 14734 27044 14740 27056
rect 8864 27016 14740 27044
rect 7929 27007 7987 27013
rect 14734 27004 14740 27016
rect 14792 27004 14798 27056
rect 14936 27053 14964 27084
rect 15289 27081 15301 27115
rect 15335 27112 15347 27115
rect 15378 27112 15384 27124
rect 15335 27084 15384 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 15378 27072 15384 27084
rect 15436 27072 15442 27124
rect 16117 27115 16175 27121
rect 16117 27081 16129 27115
rect 16163 27112 16175 27115
rect 16574 27112 16580 27124
rect 16163 27084 16580 27112
rect 16163 27081 16175 27084
rect 16117 27075 16175 27081
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17865 27115 17923 27121
rect 17865 27112 17877 27115
rect 16908 27084 17877 27112
rect 16908 27072 16914 27084
rect 17865 27081 17877 27084
rect 17911 27081 17923 27115
rect 17865 27075 17923 27081
rect 17954 27072 17960 27124
rect 18012 27112 18018 27124
rect 19058 27112 19064 27124
rect 18012 27084 19064 27112
rect 18012 27072 18018 27084
rect 19058 27072 19064 27084
rect 19116 27072 19122 27124
rect 19334 27112 19340 27124
rect 19306 27072 19340 27112
rect 19392 27072 19398 27124
rect 19426 27072 19432 27124
rect 19484 27072 19490 27124
rect 19518 27072 19524 27124
rect 19576 27112 19582 27124
rect 20990 27112 20996 27124
rect 19576 27084 20996 27112
rect 19576 27072 19582 27084
rect 20990 27072 20996 27084
rect 21048 27072 21054 27124
rect 14921 27047 14979 27053
rect 14921 27013 14933 27047
rect 14967 27044 14979 27047
rect 15470 27044 15476 27056
rect 14967 27016 15476 27044
rect 14967 27013 14979 27016
rect 14921 27007 14979 27013
rect 15470 27004 15476 27016
rect 15528 27004 15534 27056
rect 15838 27004 15844 27056
rect 15896 27044 15902 27056
rect 15933 27047 15991 27053
rect 15933 27044 15945 27047
rect 15896 27016 15945 27044
rect 15896 27004 15902 27016
rect 15933 27013 15945 27016
rect 15979 27044 15991 27047
rect 17405 27047 17463 27053
rect 15979 27016 17356 27044
rect 15979 27013 15991 27016
rect 15933 27007 15991 27013
rect 5721 26979 5779 26985
rect 5721 26945 5733 26979
rect 5767 26945 5779 26979
rect 5721 26939 5779 26945
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 3510 26908 3516 26920
rect 2332 26880 3516 26908
rect 3510 26868 3516 26880
rect 3568 26868 3574 26920
rect 5736 26908 5764 26939
rect 6638 26936 6644 26988
rect 6696 26976 6702 26988
rect 6733 26979 6791 26985
rect 6733 26976 6745 26979
rect 6696 26948 6745 26976
rect 6696 26936 6702 26948
rect 6733 26945 6745 26948
rect 6779 26945 6791 26979
rect 6733 26939 6791 26945
rect 7006 26936 7012 26988
rect 7064 26976 7070 26988
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 7064 26948 7113 26976
rect 7064 26936 7070 26948
rect 7101 26945 7113 26948
rect 7147 26976 7159 26979
rect 7742 26976 7748 26988
rect 7147 26948 7748 26976
rect 7147 26945 7159 26948
rect 7101 26939 7159 26945
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 6178 26908 6184 26920
rect 5736 26880 6184 26908
rect 6178 26868 6184 26880
rect 6236 26868 6242 26920
rect 6549 26911 6607 26917
rect 6549 26877 6561 26911
rect 6595 26908 6607 26911
rect 6822 26908 6828 26920
rect 6595 26880 6828 26908
rect 6595 26877 6607 26880
rect 6549 26871 6607 26877
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7650 26868 7656 26920
rect 7708 26908 7714 26920
rect 8036 26908 8064 26939
rect 8478 26936 8484 26988
rect 8536 26976 8542 26988
rect 10137 26979 10195 26985
rect 10137 26976 10149 26979
rect 8536 26948 10149 26976
rect 8536 26936 8542 26948
rect 10137 26945 10149 26948
rect 10183 26976 10195 26979
rect 10183 26948 11100 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 7708 26880 8064 26908
rect 7708 26868 7714 26880
rect 8938 26868 8944 26920
rect 8996 26868 9002 26920
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 10229 26911 10287 26917
rect 10229 26908 10241 26911
rect 9456 26880 10241 26908
rect 9456 26868 9462 26880
rect 10229 26877 10241 26880
rect 10275 26877 10287 26911
rect 10229 26871 10287 26877
rect 10318 26868 10324 26920
rect 10376 26868 10382 26920
rect 11072 26908 11100 26948
rect 11146 26936 11152 26988
rect 11204 26936 11210 26988
rect 11256 26948 12297 26976
rect 11256 26908 11284 26948
rect 11072 26880 11284 26908
rect 11701 26911 11759 26917
rect 11701 26877 11713 26911
rect 11747 26877 11759 26911
rect 12269 26908 12297 26948
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 13170 26976 13176 26988
rect 12400 26948 13176 26976
rect 12400 26936 12406 26948
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 14090 26936 14096 26988
rect 14148 26936 14154 26988
rect 14182 26936 14188 26988
rect 14240 26976 14246 26988
rect 14277 26979 14335 26985
rect 14277 26976 14289 26979
rect 14240 26948 14289 26976
rect 14240 26936 14246 26948
rect 14277 26945 14289 26948
rect 14323 26945 14335 26979
rect 14277 26939 14335 26945
rect 15102 26936 15108 26988
rect 15160 26936 15166 26988
rect 15378 26936 15384 26988
rect 15436 26976 15442 26988
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15436 26948 15761 26976
rect 15436 26936 15442 26948
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 17034 26936 17040 26988
rect 17092 26936 17098 26988
rect 17218 26936 17224 26988
rect 17276 26936 17282 26988
rect 17328 26976 17356 27016
rect 17405 27013 17417 27047
rect 17451 27044 17463 27047
rect 19306 27044 19334 27072
rect 17451 27016 19334 27044
rect 17451 27013 17463 27016
rect 17405 27007 17463 27013
rect 21634 27004 21640 27056
rect 21692 27044 21698 27056
rect 22250 27047 22308 27053
rect 22250 27044 22262 27047
rect 21692 27016 22262 27044
rect 21692 27004 21698 27016
rect 22250 27013 22262 27016
rect 22296 27013 22308 27047
rect 22250 27007 22308 27013
rect 22370 27004 22376 27056
rect 22428 27004 22434 27056
rect 23198 27004 23204 27056
rect 23256 27044 23262 27056
rect 23256 27016 27844 27044
rect 23256 27004 23262 27016
rect 17954 26976 17960 26988
rect 17328 26948 17960 26976
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18046 26936 18052 26988
rect 18104 26936 18110 26988
rect 19426 26982 19432 26988
rect 19352 26976 19432 26982
rect 18156 26954 19432 26976
rect 18156 26948 19380 26954
rect 17862 26908 17868 26920
rect 12269 26880 17868 26908
rect 11701 26871 11759 26877
rect 4062 26800 4068 26852
rect 4120 26800 4126 26852
rect 4154 26800 4160 26852
rect 4212 26840 4218 26852
rect 5077 26843 5135 26849
rect 5077 26840 5089 26843
rect 4212 26812 5089 26840
rect 4212 26800 4218 26812
rect 5077 26809 5089 26812
rect 5123 26809 5135 26843
rect 5077 26803 5135 26809
rect 5902 26800 5908 26852
rect 5960 26800 5966 26852
rect 7006 26800 7012 26852
rect 7064 26800 7070 26852
rect 9309 26843 9367 26849
rect 9309 26809 9321 26843
rect 9355 26840 9367 26843
rect 11716 26840 11744 26871
rect 17862 26868 17868 26880
rect 17920 26868 17926 26920
rect 9355 26812 11744 26840
rect 9355 26809 9367 26812
rect 9309 26803 9367 26809
rect 11974 26800 11980 26852
rect 12032 26840 12038 26852
rect 12713 26843 12771 26849
rect 12713 26840 12725 26843
rect 12032 26812 12725 26840
rect 12032 26800 12038 26812
rect 12713 26809 12725 26812
rect 12759 26840 12771 26843
rect 12802 26840 12808 26852
rect 12759 26812 12808 26840
rect 12759 26809 12771 26812
rect 12713 26803 12771 26809
rect 12802 26800 12808 26812
rect 12860 26840 12866 26852
rect 13541 26843 13599 26849
rect 13541 26840 13553 26843
rect 12860 26812 13553 26840
rect 12860 26800 12866 26812
rect 13541 26809 13553 26812
rect 13587 26840 13599 26843
rect 13630 26840 13636 26852
rect 13587 26812 13636 26840
rect 13587 26809 13599 26812
rect 13541 26803 13599 26809
rect 13630 26800 13636 26812
rect 13688 26800 13694 26852
rect 14461 26843 14519 26849
rect 14461 26809 14473 26843
rect 14507 26840 14519 26843
rect 16298 26840 16304 26852
rect 14507 26812 16304 26840
rect 14507 26809 14519 26812
rect 14461 26803 14519 26809
rect 16298 26800 16304 26812
rect 16356 26800 16362 26852
rect 16574 26800 16580 26852
rect 16632 26840 16638 26852
rect 17218 26840 17224 26852
rect 16632 26812 17224 26840
rect 16632 26800 16638 26812
rect 17218 26800 17224 26812
rect 17276 26840 17282 26852
rect 18156 26840 18184 26948
rect 19426 26936 19432 26954
rect 19484 26936 19490 26988
rect 19610 26985 19616 26988
rect 19605 26939 19616 26985
rect 19610 26936 19616 26939
rect 19668 26936 19674 26988
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26945 20499 26979
rect 20441 26939 20499 26945
rect 18414 26868 18420 26920
rect 18472 26868 18478 26920
rect 18509 26911 18567 26917
rect 18509 26877 18521 26911
rect 18555 26908 18567 26911
rect 18690 26908 18696 26920
rect 18555 26880 18696 26908
rect 18555 26877 18567 26880
rect 18509 26871 18567 26877
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 18969 26911 19027 26917
rect 18969 26877 18981 26911
rect 19015 26908 19027 26911
rect 20456 26908 20484 26939
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20772 26948 21097 26976
rect 20772 26936 20778 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 21174 26936 21180 26988
rect 21232 26976 21238 26988
rect 22388 26976 22416 27004
rect 21232 26948 22416 26976
rect 24029 26979 24087 26985
rect 21232 26936 21238 26948
rect 24029 26945 24041 26979
rect 24075 26976 24087 26979
rect 24302 26976 24308 26988
rect 24075 26948 24308 26976
rect 24075 26945 24087 26948
rect 24029 26939 24087 26945
rect 24302 26936 24308 26948
rect 24360 26936 24366 26988
rect 24489 26979 24547 26985
rect 24489 26945 24501 26979
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 19015 26880 19334 26908
rect 19015 26877 19027 26880
rect 18969 26871 19027 26877
rect 17276 26812 18184 26840
rect 18432 26840 18460 26868
rect 18785 26843 18843 26849
rect 18785 26840 18797 26843
rect 18432 26812 18797 26840
rect 17276 26800 17282 26812
rect 18785 26809 18797 26812
rect 18831 26809 18843 26843
rect 19306 26840 19334 26880
rect 19689 26880 20484 26908
rect 19689 26840 19717 26880
rect 21542 26868 21548 26920
rect 21600 26908 21606 26920
rect 22005 26911 22063 26917
rect 22005 26908 22017 26911
rect 21600 26880 22017 26908
rect 21600 26868 21606 26880
rect 22005 26877 22017 26880
rect 22051 26877 22063 26911
rect 22005 26871 22063 26877
rect 24504 26840 24532 26939
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 25481 26979 25539 26985
rect 25481 26976 25493 26979
rect 24820 26948 25493 26976
rect 24820 26936 24826 26948
rect 25481 26945 25493 26948
rect 25527 26945 25539 26979
rect 25481 26939 25539 26945
rect 25866 26936 25872 26988
rect 25924 26976 25930 26988
rect 27157 26979 27215 26985
rect 25924 26948 27108 26976
rect 25924 26936 25930 26948
rect 24946 26868 24952 26920
rect 25004 26908 25010 26920
rect 25225 26911 25283 26917
rect 25225 26908 25237 26911
rect 25004 26880 25237 26908
rect 25004 26868 25010 26880
rect 25225 26877 25237 26880
rect 25271 26877 25283 26911
rect 27080 26908 27108 26948
rect 27157 26945 27169 26979
rect 27203 26974 27215 26979
rect 27264 26974 27292 27016
rect 27816 26985 27844 27016
rect 27203 26946 27292 26974
rect 27341 26979 27399 26985
rect 27203 26945 27215 26946
rect 27157 26939 27215 26945
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 27801 26979 27859 26985
rect 27801 26945 27813 26979
rect 27847 26945 27859 26979
rect 27801 26939 27859 26945
rect 27985 26979 28043 26985
rect 27985 26945 27997 26979
rect 28031 26976 28043 26979
rect 28074 26976 28080 26988
rect 28031 26948 28080 26976
rect 28031 26945 28043 26948
rect 27985 26939 28043 26945
rect 27356 26908 27384 26939
rect 28074 26936 28080 26948
rect 28132 26936 28138 26988
rect 27080 26880 27384 26908
rect 25225 26871 25283 26877
rect 19306 26812 19717 26840
rect 20180 26812 21036 26840
rect 18785 26803 18843 26809
rect 7561 26775 7619 26781
rect 7561 26741 7573 26775
rect 7607 26772 7619 26775
rect 9214 26772 9220 26784
rect 7607 26744 9220 26772
rect 7607 26741 7619 26744
rect 7561 26735 7619 26741
rect 9214 26732 9220 26744
rect 9272 26732 9278 26784
rect 15102 26732 15108 26784
rect 15160 26772 15166 26784
rect 17678 26772 17684 26784
rect 15160 26744 17684 26772
rect 15160 26732 15166 26744
rect 17678 26732 17684 26744
rect 17736 26732 17742 26784
rect 17862 26732 17868 26784
rect 17920 26772 17926 26784
rect 19334 26772 19340 26784
rect 17920 26744 19340 26772
rect 17920 26732 17926 26744
rect 19334 26732 19340 26744
rect 19392 26732 19398 26784
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 20180 26772 20208 26812
rect 19668 26744 20208 26772
rect 20257 26775 20315 26781
rect 19668 26732 19674 26744
rect 20257 26741 20269 26775
rect 20303 26772 20315 26775
rect 20438 26772 20444 26784
rect 20303 26744 20444 26772
rect 20303 26741 20315 26744
rect 20257 26735 20315 26741
rect 20438 26732 20444 26744
rect 20496 26732 20502 26784
rect 20530 26732 20536 26784
rect 20588 26772 20594 26784
rect 20901 26775 20959 26781
rect 20901 26772 20913 26775
rect 20588 26744 20913 26772
rect 20588 26732 20594 26744
rect 20901 26741 20913 26744
rect 20947 26741 20959 26775
rect 21008 26772 21036 26812
rect 22940 26812 24532 26840
rect 22940 26772 22968 26812
rect 21008 26744 22968 26772
rect 20901 26735 20959 26741
rect 23382 26732 23388 26784
rect 23440 26732 23446 26784
rect 23750 26732 23756 26784
rect 23808 26772 23814 26784
rect 23845 26775 23903 26781
rect 23845 26772 23857 26775
rect 23808 26744 23857 26772
rect 23808 26732 23814 26744
rect 23845 26741 23857 26744
rect 23891 26741 23903 26775
rect 23845 26735 23903 26741
rect 23934 26732 23940 26784
rect 23992 26772 23998 26784
rect 24581 26775 24639 26781
rect 24581 26772 24593 26775
rect 23992 26744 24593 26772
rect 23992 26732 23998 26744
rect 24581 26741 24593 26744
rect 24627 26741 24639 26775
rect 24581 26735 24639 26741
rect 25958 26732 25964 26784
rect 26016 26772 26022 26784
rect 26605 26775 26663 26781
rect 26605 26772 26617 26775
rect 26016 26744 26617 26772
rect 26016 26732 26022 26744
rect 26605 26741 26617 26744
rect 26651 26741 26663 26775
rect 26605 26735 26663 26741
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 3786 26528 3792 26580
rect 3844 26568 3850 26580
rect 5994 26568 6000 26580
rect 3844 26540 6000 26568
rect 3844 26528 3850 26540
rect 5994 26528 6000 26540
rect 6052 26528 6058 26580
rect 7561 26571 7619 26577
rect 7561 26537 7573 26571
rect 7607 26568 7619 26571
rect 8386 26568 8392 26580
rect 7607 26540 8392 26568
rect 7607 26537 7619 26540
rect 7561 26531 7619 26537
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 8496 26540 9536 26568
rect 4982 26500 4988 26512
rect 3436 26472 4988 26500
rect 3436 26441 3464 26472
rect 3421 26435 3479 26441
rect 3421 26401 3433 26435
rect 3467 26401 3479 26435
rect 3421 26395 3479 26401
rect 4154 26392 4160 26444
rect 4212 26392 4218 26444
rect 4816 26441 4844 26472
rect 4982 26460 4988 26472
rect 5040 26460 5046 26512
rect 5810 26460 5816 26512
rect 5868 26500 5874 26512
rect 7282 26500 7288 26512
rect 5868 26472 7288 26500
rect 5868 26460 5874 26472
rect 4801 26435 4859 26441
rect 4801 26401 4813 26435
rect 4847 26401 4859 26435
rect 4801 26395 4859 26401
rect 5629 26435 5687 26441
rect 5629 26401 5641 26435
rect 5675 26432 5687 26435
rect 6454 26432 6460 26444
rect 5675 26404 6460 26432
rect 5675 26401 5687 26404
rect 5629 26395 5687 26401
rect 6454 26392 6460 26404
rect 6512 26392 6518 26444
rect 7116 26441 7144 26472
rect 7282 26460 7288 26472
rect 7340 26460 7346 26512
rect 8496 26500 8524 26540
rect 7392 26472 8524 26500
rect 8573 26503 8631 26509
rect 7101 26435 7159 26441
rect 7101 26401 7113 26435
rect 7147 26401 7159 26435
rect 7101 26395 7159 26401
rect 1762 26324 1768 26376
rect 1820 26364 1826 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 1820 26336 3985 26364
rect 1820 26324 1826 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4525 26367 4583 26373
rect 4525 26333 4537 26367
rect 4571 26364 4583 26367
rect 5074 26364 5080 26376
rect 4571 26336 5080 26364
rect 4571 26333 4583 26336
rect 4525 26327 4583 26333
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 5258 26324 5264 26376
rect 5316 26324 5322 26376
rect 5350 26324 5356 26376
rect 5408 26364 5414 26376
rect 5445 26367 5503 26373
rect 5445 26364 5457 26367
rect 5408 26336 5457 26364
rect 5408 26324 5414 26336
rect 5445 26333 5457 26336
rect 5491 26333 5503 26367
rect 5445 26327 5503 26333
rect 6362 26324 6368 26376
rect 6420 26364 6426 26376
rect 6825 26367 6883 26373
rect 6825 26364 6837 26367
rect 6420 26336 6837 26364
rect 6420 26324 6426 26336
rect 6825 26333 6837 26336
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 6914 26324 6920 26376
rect 6972 26364 6978 26376
rect 7009 26367 7067 26373
rect 7009 26364 7021 26367
rect 6972 26336 7021 26364
rect 6972 26324 6978 26336
rect 7009 26333 7021 26336
rect 7055 26333 7067 26367
rect 7009 26327 7067 26333
rect 1670 26256 1676 26308
rect 1728 26256 1734 26308
rect 4062 26256 4068 26308
rect 4120 26256 4126 26308
rect 4982 26256 4988 26308
rect 5040 26296 5046 26308
rect 6380 26296 6408 26324
rect 5040 26268 6408 26296
rect 5040 26256 5046 26268
rect 6638 26256 6644 26308
rect 6696 26256 6702 26308
rect 5718 26188 5724 26240
rect 5776 26228 5782 26240
rect 7392 26228 7420 26472
rect 8573 26469 8585 26503
rect 8619 26500 8631 26503
rect 8662 26500 8668 26512
rect 8619 26472 8668 26500
rect 8619 26469 8631 26472
rect 8573 26463 8631 26469
rect 8662 26460 8668 26472
rect 8720 26500 8726 26512
rect 8720 26472 9260 26500
rect 8720 26460 8726 26472
rect 8205 26435 8263 26441
rect 8205 26401 8217 26435
rect 8251 26432 8263 26435
rect 9122 26432 9128 26444
rect 8251 26404 9128 26432
rect 8251 26401 8263 26404
rect 8205 26395 8263 26401
rect 9122 26392 9128 26404
rect 9180 26392 9186 26444
rect 7742 26324 7748 26376
rect 7800 26324 7806 26376
rect 9232 26364 9260 26472
rect 9508 26432 9536 26540
rect 9582 26528 9588 26580
rect 9640 26568 9646 26580
rect 10778 26568 10784 26580
rect 9640 26540 10784 26568
rect 9640 26528 9646 26540
rect 10778 26528 10784 26540
rect 10836 26528 10842 26580
rect 11974 26528 11980 26580
rect 12032 26528 12038 26580
rect 13998 26568 14004 26580
rect 13556 26540 14004 26568
rect 10689 26503 10747 26509
rect 10689 26469 10701 26503
rect 10735 26500 10747 26503
rect 11882 26500 11888 26512
rect 10735 26472 11888 26500
rect 10735 26469 10747 26472
rect 10689 26463 10747 26469
rect 11882 26460 11888 26472
rect 11940 26460 11946 26512
rect 9508 26404 9674 26432
rect 9493 26367 9551 26373
rect 9232 26360 9444 26364
rect 9493 26360 9505 26367
rect 9232 26336 9505 26360
rect 9416 26333 9505 26336
rect 9539 26333 9551 26367
rect 9416 26332 9551 26333
rect 9493 26327 9551 26332
rect 5776 26200 7420 26228
rect 5776 26188 5782 26200
rect 8570 26188 8576 26240
rect 8628 26188 8634 26240
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9493 26231 9551 26237
rect 9493 26228 9505 26231
rect 9364 26200 9505 26228
rect 9364 26188 9370 26200
rect 9493 26197 9505 26200
rect 9539 26197 9551 26231
rect 9646 26228 9674 26404
rect 9858 26392 9864 26444
rect 9916 26432 9922 26444
rect 11992 26441 12020 26528
rect 12269 26472 13308 26500
rect 11977 26435 12035 26441
rect 9916 26404 11652 26432
rect 9916 26392 9922 26404
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10137 26367 10195 26373
rect 10137 26364 10149 26367
rect 10008 26336 10149 26364
rect 10008 26324 10014 26336
rect 10137 26333 10149 26336
rect 10183 26333 10195 26367
rect 10137 26327 10195 26333
rect 10410 26324 10416 26376
rect 10468 26324 10474 26376
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26364 10563 26367
rect 10686 26364 10692 26376
rect 10551 26336 10692 26364
rect 10551 26333 10563 26336
rect 10505 26327 10563 26333
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 11624 26373 11652 26404
rect 11977 26401 11989 26435
rect 12023 26401 12035 26435
rect 11977 26395 12035 26401
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26364 11667 26367
rect 12269 26364 12297 26472
rect 13280 26444 13308 26472
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12400 26404 12817 26432
rect 12400 26392 12406 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 13262 26392 13268 26444
rect 13320 26392 13326 26444
rect 11655 26336 12297 26364
rect 12621 26367 12679 26373
rect 11655 26333 11667 26336
rect 11609 26327 11667 26333
rect 12621 26333 12633 26367
rect 12667 26364 12679 26367
rect 13556 26364 13584 26540
rect 13998 26528 14004 26540
rect 14056 26568 14062 26580
rect 17865 26571 17923 26577
rect 17865 26568 17877 26571
rect 14056 26540 17877 26568
rect 14056 26528 14062 26540
rect 17865 26537 17877 26540
rect 17911 26537 17923 26571
rect 17865 26531 17923 26537
rect 18877 26571 18935 26577
rect 18877 26537 18889 26571
rect 18923 26568 18935 26571
rect 20898 26568 20904 26580
rect 18923 26540 20904 26568
rect 18923 26537 18935 26540
rect 18877 26531 18935 26537
rect 20898 26528 20904 26540
rect 20956 26528 20962 26580
rect 21082 26528 21088 26580
rect 21140 26568 21146 26580
rect 21140 26540 26188 26568
rect 21140 26528 21146 26540
rect 13630 26460 13636 26512
rect 13688 26460 13694 26512
rect 14458 26460 14464 26512
rect 14516 26500 14522 26512
rect 15102 26500 15108 26512
rect 14516 26472 15108 26500
rect 14516 26460 14522 26472
rect 15102 26460 15108 26472
rect 15160 26460 15166 26512
rect 16114 26500 16120 26512
rect 15212 26472 16120 26500
rect 14642 26392 14648 26444
rect 14700 26432 14706 26444
rect 14700 26404 14964 26432
rect 14700 26392 14706 26404
rect 12667 26336 13584 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 14826 26324 14832 26376
rect 14884 26324 14890 26376
rect 14936 26373 14964 26404
rect 15212 26373 15240 26472
rect 16114 26460 16120 26472
rect 16172 26460 16178 26512
rect 17954 26460 17960 26512
rect 18012 26500 18018 26512
rect 18785 26503 18843 26509
rect 18785 26500 18797 26503
rect 18012 26472 18797 26500
rect 18012 26460 18018 26472
rect 18785 26469 18797 26472
rect 18831 26500 18843 26503
rect 19242 26500 19248 26512
rect 18831 26472 19248 26500
rect 18831 26469 18843 26472
rect 18785 26463 18843 26469
rect 19242 26460 19248 26472
rect 19300 26460 19306 26512
rect 22922 26460 22928 26512
rect 22980 26500 22986 26512
rect 23382 26500 23388 26512
rect 22980 26472 23388 26500
rect 22980 26460 22986 26472
rect 23382 26460 23388 26472
rect 23440 26460 23446 26512
rect 17678 26392 17684 26444
rect 17736 26432 17742 26444
rect 17736 26404 19564 26432
rect 17736 26392 17742 26404
rect 14922 26367 14980 26373
rect 14922 26333 14934 26367
rect 14968 26333 14980 26367
rect 14922 26327 14980 26333
rect 15197 26367 15255 26373
rect 15197 26333 15209 26367
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 15335 26367 15393 26373
rect 15335 26333 15347 26367
rect 15381 26364 15393 26367
rect 16114 26364 16120 26376
rect 15381 26336 16120 26364
rect 15381 26333 15393 26336
rect 15335 26327 15393 26333
rect 16114 26324 16120 26336
rect 16172 26324 16178 26376
rect 16482 26324 16488 26376
rect 16540 26324 16546 26376
rect 17310 26324 17316 26376
rect 17368 26364 17374 26376
rect 17368 26336 18552 26364
rect 17368 26324 17374 26336
rect 10318 26256 10324 26308
rect 10376 26256 10382 26308
rect 11054 26256 11060 26308
rect 11112 26296 11118 26308
rect 12437 26299 12495 26305
rect 12437 26296 12449 26299
rect 11112 26268 12449 26296
rect 11112 26256 11118 26268
rect 12437 26265 12449 26268
rect 12483 26296 12495 26299
rect 12986 26296 12992 26308
rect 12483 26268 12992 26296
rect 12483 26265 12495 26268
rect 12437 26259 12495 26265
rect 12986 26256 12992 26268
rect 13044 26256 13050 26308
rect 15105 26299 15163 26305
rect 15105 26265 15117 26299
rect 15151 26296 15163 26299
rect 15930 26296 15936 26308
rect 15151 26268 15936 26296
rect 15151 26265 15163 26268
rect 15105 26259 15163 26265
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 16022 26256 16028 26308
rect 16080 26296 16086 26308
rect 16730 26299 16788 26305
rect 16730 26296 16742 26299
rect 16080 26268 16742 26296
rect 16080 26256 16086 26268
rect 16730 26265 16742 26268
rect 16776 26265 16788 26299
rect 16730 26259 16788 26265
rect 18417 26299 18475 26305
rect 18417 26265 18429 26299
rect 18463 26265 18475 26299
rect 18524 26296 18552 26336
rect 19426 26324 19432 26376
rect 19484 26324 19490 26376
rect 19536 26364 19564 26404
rect 20456 26404 21404 26432
rect 20456 26364 20484 26404
rect 21269 26367 21327 26373
rect 21269 26364 21281 26367
rect 19536 26336 20484 26364
rect 20548 26336 21281 26364
rect 19674 26299 19732 26305
rect 19674 26296 19686 26299
rect 18524 26268 19686 26296
rect 18417 26259 18475 26265
rect 19674 26265 19686 26268
rect 19720 26265 19732 26299
rect 19674 26259 19732 26265
rect 10778 26228 10784 26240
rect 9646 26200 10784 26228
rect 9493 26191 9551 26197
rect 10778 26188 10784 26200
rect 10836 26228 10842 26240
rect 11422 26228 11428 26240
rect 10836 26200 11428 26228
rect 10836 26188 10842 26200
rect 11422 26188 11428 26200
rect 11480 26188 11486 26240
rect 13630 26188 13636 26240
rect 13688 26188 13694 26240
rect 14642 26188 14648 26240
rect 14700 26228 14706 26240
rect 15286 26228 15292 26240
rect 14700 26200 15292 26228
rect 14700 26188 14706 26200
rect 15286 26188 15292 26200
rect 15344 26188 15350 26240
rect 15470 26188 15476 26240
rect 15528 26188 15534 26240
rect 18432 26228 18460 26259
rect 19794 26256 19800 26308
rect 19852 26296 19858 26308
rect 20548 26296 20576 26336
rect 21269 26333 21281 26336
rect 21315 26333 21327 26367
rect 21376 26364 21404 26404
rect 22388 26404 23980 26432
rect 22278 26364 22284 26376
rect 21376 26336 22284 26364
rect 21269 26327 21327 26333
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 19852 26268 20576 26296
rect 19852 26256 19858 26268
rect 20898 26256 20904 26308
rect 20956 26296 20962 26308
rect 21514 26299 21572 26305
rect 21514 26296 21526 26299
rect 20956 26268 21526 26296
rect 20956 26256 20962 26268
rect 21514 26265 21526 26268
rect 21560 26265 21572 26299
rect 21514 26259 21572 26265
rect 21634 26256 21640 26308
rect 21692 26296 21698 26308
rect 22388 26296 22416 26404
rect 22462 26324 22468 26376
rect 22520 26364 22526 26376
rect 22738 26364 22744 26376
rect 22520 26336 22744 26364
rect 22520 26324 22526 26336
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23106 26324 23112 26376
rect 23164 26324 23170 26376
rect 23290 26324 23296 26376
rect 23348 26324 23354 26376
rect 23952 26373 23980 26404
rect 24670 26392 24676 26444
rect 24728 26432 24734 26444
rect 25133 26435 25191 26441
rect 25133 26432 25145 26435
rect 24728 26404 25145 26432
rect 24728 26392 24734 26404
rect 25133 26401 25145 26404
rect 25179 26401 25191 26435
rect 26160 26432 26188 26540
rect 26160 26404 27088 26432
rect 25133 26395 25191 26401
rect 23753 26367 23811 26373
rect 23753 26333 23765 26367
rect 23799 26333 23811 26367
rect 23753 26327 23811 26333
rect 23937 26367 23995 26373
rect 23937 26333 23949 26367
rect 23983 26333 23995 26367
rect 23937 26327 23995 26333
rect 21692 26268 22416 26296
rect 22460 26268 22784 26296
rect 21692 26256 21698 26268
rect 18782 26228 18788 26240
rect 18432 26200 18788 26228
rect 18782 26188 18788 26200
rect 18840 26188 18846 26240
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 20346 26228 20352 26240
rect 19484 26200 20352 26228
rect 19484 26188 19490 26200
rect 20346 26188 20352 26200
rect 20404 26188 20410 26240
rect 20806 26188 20812 26240
rect 20864 26188 20870 26240
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 22460 26228 22488 26268
rect 21048 26200 22488 26228
rect 21048 26188 21054 26200
rect 22646 26188 22652 26240
rect 22704 26188 22710 26240
rect 22756 26228 22784 26268
rect 23198 26256 23204 26308
rect 23256 26256 23262 26308
rect 23768 26228 23796 26327
rect 26142 26324 26148 26376
rect 26200 26364 26206 26376
rect 26973 26367 27031 26373
rect 26973 26364 26985 26367
rect 26200 26336 26985 26364
rect 26200 26324 26206 26336
rect 26973 26333 26985 26336
rect 27019 26333 27031 26367
rect 27060 26364 27088 26404
rect 27229 26367 27287 26373
rect 27229 26364 27241 26367
rect 27060 26336 27241 26364
rect 26973 26327 27031 26333
rect 27229 26333 27241 26336
rect 27275 26333 27287 26367
rect 27229 26327 27287 26333
rect 23842 26256 23848 26308
rect 23900 26256 23906 26308
rect 24854 26256 24860 26308
rect 24912 26296 24918 26308
rect 25378 26299 25436 26305
rect 25378 26296 25390 26299
rect 24912 26268 25390 26296
rect 24912 26256 24918 26268
rect 25378 26265 25390 26268
rect 25424 26265 25436 26299
rect 25378 26259 25436 26265
rect 22756 26200 23796 26228
rect 26510 26188 26516 26240
rect 26568 26188 26574 26240
rect 28350 26188 28356 26240
rect 28408 26188 28414 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 2406 25984 2412 26036
rect 2464 25984 2470 26036
rect 5902 26024 5908 26036
rect 2746 25996 5908 26024
rect 2746 25956 2774 25996
rect 5902 25984 5908 25996
rect 5960 25984 5966 26036
rect 7466 25984 7472 26036
rect 7524 26024 7530 26036
rect 8113 26027 8171 26033
rect 8113 26024 8125 26027
rect 7524 25996 8125 26024
rect 7524 25984 7530 25996
rect 8113 25993 8125 25996
rect 8159 26024 8171 26027
rect 8570 26024 8576 26036
rect 8159 25996 8576 26024
rect 8159 25993 8171 25996
rect 8113 25987 8171 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 9401 26027 9459 26033
rect 9401 25993 9413 26027
rect 9447 26024 9459 26027
rect 9490 26024 9496 26036
rect 9447 25996 9496 26024
rect 9447 25993 9459 25996
rect 9401 25987 9459 25993
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 9766 25984 9772 26036
rect 9824 25984 9830 26036
rect 9858 25984 9864 26036
rect 9916 25984 9922 26036
rect 11057 26027 11115 26033
rect 11057 25993 11069 26027
rect 11103 26024 11115 26027
rect 11146 26024 11152 26036
rect 11103 25996 11152 26024
rect 11103 25993 11115 25996
rect 11057 25987 11115 25993
rect 11146 25984 11152 25996
rect 11204 25984 11210 26036
rect 11422 25984 11428 26036
rect 11480 26024 11486 26036
rect 19613 26027 19671 26033
rect 11480 25996 19334 26024
rect 11480 25984 11486 25996
rect 2424 25928 2774 25956
rect 2424 25897 2452 25928
rect 3418 25916 3424 25968
rect 3476 25916 3482 25968
rect 6917 25959 6975 25965
rect 6917 25925 6929 25959
rect 6963 25956 6975 25959
rect 9122 25956 9128 25968
rect 6963 25928 9128 25956
rect 6963 25925 6975 25928
rect 6917 25919 6975 25925
rect 9122 25916 9128 25928
rect 9180 25956 9186 25968
rect 9180 25928 9260 25956
rect 9180 25916 9186 25928
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 3694 25888 3700 25900
rect 2639 25860 3700 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 1394 25780 1400 25832
rect 1452 25820 1458 25832
rect 1854 25820 1860 25832
rect 1452 25792 1860 25820
rect 1452 25780 1458 25792
rect 1854 25780 1860 25792
rect 1912 25820 1918 25832
rect 2133 25823 2191 25829
rect 2133 25820 2145 25823
rect 1912 25792 2145 25820
rect 1912 25780 1918 25792
rect 2133 25789 2145 25792
rect 2179 25789 2191 25823
rect 2133 25783 2191 25789
rect 2314 25780 2320 25832
rect 2372 25820 2378 25832
rect 2608 25820 2636 25851
rect 3694 25848 3700 25860
rect 3752 25848 3758 25900
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 5626 25888 5632 25900
rect 4856 25860 5632 25888
rect 4856 25848 4862 25860
rect 5626 25848 5632 25860
rect 5684 25848 5690 25900
rect 5905 25891 5963 25897
rect 5905 25857 5917 25891
rect 5951 25888 5963 25891
rect 6454 25888 6460 25900
rect 5951 25860 6460 25888
rect 5951 25857 5963 25860
rect 5905 25851 5963 25857
rect 6454 25848 6460 25860
rect 6512 25848 6518 25900
rect 7101 25891 7159 25897
rect 7101 25857 7113 25891
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7745 25891 7803 25897
rect 7745 25857 7757 25891
rect 7791 25888 7803 25891
rect 8202 25888 8208 25900
rect 7791 25860 8208 25888
rect 7791 25857 7803 25860
rect 7745 25851 7803 25857
rect 2372 25792 2636 25820
rect 2372 25780 2378 25792
rect 2958 25780 2964 25832
rect 3016 25780 3022 25832
rect 7116 25820 7144 25851
rect 8202 25848 8208 25860
rect 8260 25848 8266 25900
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 9232 25888 9260 25928
rect 9306 25916 9312 25968
rect 9364 25956 9370 25968
rect 15166 25959 15224 25965
rect 15166 25956 15178 25959
rect 9364 25928 15178 25956
rect 9364 25916 9370 25928
rect 15166 25925 15178 25928
rect 15212 25925 15224 25959
rect 15166 25919 15224 25925
rect 16853 25959 16911 25965
rect 16853 25925 16865 25959
rect 16899 25956 16911 25959
rect 16942 25956 16948 25968
rect 16899 25928 16948 25956
rect 16899 25925 16911 25928
rect 16853 25919 16911 25925
rect 16942 25916 16948 25928
rect 17000 25916 17006 25968
rect 17221 25959 17279 25965
rect 17221 25925 17233 25959
rect 17267 25956 17279 25959
rect 18598 25956 18604 25968
rect 17267 25928 18604 25956
rect 17267 25925 17279 25928
rect 17221 25919 17279 25925
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 19306 25956 19334 25996
rect 19613 25993 19625 26027
rect 19659 26024 19671 26027
rect 20070 26024 20076 26036
rect 19659 25996 20076 26024
rect 19659 25993 19671 25996
rect 19613 25987 19671 25993
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 21177 26027 21235 26033
rect 21177 25993 21189 26027
rect 21223 26024 21235 26027
rect 25038 26024 25044 26036
rect 21223 25996 25044 26024
rect 21223 25993 21235 25996
rect 21177 25987 21235 25993
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 20990 25956 20996 25968
rect 19306 25928 20996 25956
rect 20990 25916 20996 25928
rect 21048 25916 21054 25968
rect 22278 25965 22284 25968
rect 22261 25959 22284 25965
rect 22261 25925 22273 25959
rect 22261 25919 22284 25925
rect 22278 25916 22284 25919
rect 22336 25916 22342 25968
rect 23014 25956 23020 25968
rect 22388 25928 23020 25956
rect 10502 25888 10508 25900
rect 9232 25860 10508 25888
rect 10502 25848 10508 25860
rect 10560 25888 10566 25900
rect 10689 25891 10747 25897
rect 10689 25888 10701 25891
rect 10560 25860 10701 25888
rect 10560 25848 10566 25860
rect 10689 25857 10701 25860
rect 10735 25857 10747 25891
rect 10873 25891 10931 25897
rect 10873 25888 10885 25891
rect 10689 25851 10747 25857
rect 10796 25860 10885 25888
rect 7116 25792 8524 25820
rect 1670 25712 1676 25764
rect 1728 25752 1734 25764
rect 2590 25752 2596 25764
rect 1728 25724 2596 25752
rect 1728 25712 1734 25724
rect 2590 25712 2596 25724
rect 2648 25752 2654 25764
rect 4709 25755 4767 25761
rect 4709 25752 4721 25755
rect 2648 25724 4721 25752
rect 2648 25712 2654 25724
rect 4709 25721 4721 25724
rect 4755 25721 4767 25755
rect 4709 25715 4767 25721
rect 5902 25712 5908 25764
rect 5960 25752 5966 25764
rect 6914 25752 6920 25764
rect 5960 25724 6920 25752
rect 5960 25712 5966 25724
rect 6914 25712 6920 25724
rect 6972 25752 6978 25764
rect 7834 25752 7840 25764
rect 6972 25724 7840 25752
rect 6972 25712 6978 25724
rect 7834 25712 7840 25724
rect 7892 25712 7898 25764
rect 8110 25712 8116 25764
rect 8168 25712 8174 25764
rect 8496 25752 8524 25792
rect 8570 25780 8576 25832
rect 8628 25780 8634 25832
rect 9030 25780 9036 25832
rect 9088 25820 9094 25832
rect 9490 25820 9496 25832
rect 9088 25792 9496 25820
rect 9088 25780 9094 25792
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9640 25792 9965 25820
rect 9640 25780 9646 25792
rect 9953 25789 9965 25792
rect 9999 25789 10011 25823
rect 10796 25820 10824 25860
rect 10873 25857 10885 25860
rect 10919 25857 10931 25891
rect 10873 25851 10931 25857
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 11793 25891 11851 25897
rect 11793 25888 11805 25891
rect 11020 25860 11805 25888
rect 11020 25848 11026 25860
rect 11793 25857 11805 25860
rect 11839 25857 11851 25891
rect 12526 25888 12532 25900
rect 11793 25851 11851 25857
rect 11900 25860 12532 25888
rect 11900 25820 11928 25860
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 12710 25897 12716 25900
rect 12704 25851 12716 25897
rect 12710 25848 12716 25851
rect 12768 25848 12774 25900
rect 13446 25848 13452 25900
rect 13504 25888 13510 25900
rect 14461 25891 14519 25897
rect 14461 25888 14473 25891
rect 13504 25860 14473 25888
rect 13504 25848 13510 25860
rect 14461 25857 14473 25860
rect 14507 25857 14519 25891
rect 14461 25851 14519 25857
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25888 14979 25891
rect 16206 25888 16212 25900
rect 14967 25860 16212 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 16206 25848 16212 25860
rect 16264 25888 16270 25900
rect 16482 25888 16488 25900
rect 16264 25860 16488 25888
rect 16264 25848 16270 25860
rect 16482 25848 16488 25860
rect 16540 25848 16546 25900
rect 16666 25848 16672 25900
rect 16724 25888 16730 25900
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16724 25860 17049 25888
rect 16724 25848 16730 25860
rect 17037 25857 17049 25860
rect 17083 25888 17095 25891
rect 17494 25888 17500 25900
rect 17083 25860 17500 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 17862 25848 17868 25900
rect 17920 25888 17926 25900
rect 19153 25891 19211 25897
rect 19153 25888 19165 25891
rect 17920 25860 19165 25888
rect 17920 25848 17926 25860
rect 19153 25857 19165 25860
rect 19199 25857 19211 25891
rect 19153 25851 19211 25857
rect 19794 25848 19800 25900
rect 19852 25848 19858 25900
rect 20070 25848 20076 25900
rect 20128 25888 20134 25900
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20128 25860 20453 25888
rect 20128 25848 20134 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20530 25848 20536 25900
rect 20588 25888 20594 25900
rect 21361 25891 21419 25897
rect 21361 25888 21373 25891
rect 20588 25860 21373 25888
rect 20588 25848 20594 25860
rect 21361 25857 21373 25860
rect 21407 25857 21419 25891
rect 22388 25888 22416 25928
rect 23014 25916 23020 25928
rect 23072 25916 23078 25968
rect 23198 25916 23204 25968
rect 23256 25956 23262 25968
rect 24946 25956 24952 25968
rect 23256 25928 24952 25956
rect 23256 25916 23262 25928
rect 24946 25916 24952 25928
rect 25004 25956 25010 25968
rect 25590 25956 25596 25968
rect 25004 25928 25596 25956
rect 25004 25916 25010 25928
rect 25590 25916 25596 25928
rect 25648 25916 25654 25968
rect 21361 25851 21419 25857
rect 21468 25860 22416 25888
rect 10796 25792 11928 25820
rect 11977 25823 12035 25829
rect 9953 25783 10011 25789
rect 11977 25789 11989 25823
rect 12023 25820 12035 25823
rect 12434 25820 12440 25832
rect 12023 25792 12440 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 12434 25780 12440 25792
rect 12492 25820 12498 25832
rect 12492 25792 12537 25820
rect 12492 25780 12498 25792
rect 17770 25780 17776 25832
rect 17828 25820 17834 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 17828 25792 18061 25820
rect 17828 25780 17834 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 18230 25780 18236 25832
rect 18288 25820 18294 25832
rect 18509 25823 18567 25829
rect 18509 25820 18521 25823
rect 18288 25792 18521 25820
rect 18288 25780 18294 25792
rect 18509 25789 18521 25792
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 18598 25780 18604 25832
rect 18656 25820 18662 25832
rect 19242 25820 19248 25832
rect 18656 25792 19248 25820
rect 18656 25780 18662 25792
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 21174 25820 21180 25832
rect 20272 25792 21180 25820
rect 11146 25752 11152 25764
rect 8496 25724 11152 25752
rect 11146 25712 11152 25724
rect 11204 25752 11210 25764
rect 12250 25752 12256 25764
rect 11204 25724 12256 25752
rect 11204 25712 11210 25724
rect 12250 25712 12256 25724
rect 12308 25712 12314 25764
rect 18138 25712 18144 25764
rect 18196 25752 18202 25764
rect 20272 25761 20300 25792
rect 21174 25780 21180 25792
rect 21232 25780 21238 25832
rect 18417 25755 18475 25761
rect 18417 25752 18429 25755
rect 18196 25724 18429 25752
rect 18196 25712 18202 25724
rect 18417 25721 18429 25724
rect 18463 25752 18475 25755
rect 20257 25755 20315 25761
rect 18463 25724 19472 25752
rect 18463 25721 18475 25724
rect 18417 25715 18475 25721
rect 7282 25644 7288 25696
rect 7340 25644 7346 25696
rect 7650 25644 7656 25696
rect 7708 25684 7714 25696
rect 7926 25684 7932 25696
rect 7708 25656 7932 25684
rect 7708 25644 7714 25656
rect 7926 25644 7932 25656
rect 7984 25684 7990 25696
rect 8941 25687 8999 25693
rect 8941 25684 8953 25687
rect 7984 25656 8953 25684
rect 7984 25644 7990 25656
rect 8941 25653 8953 25656
rect 8987 25653 8999 25687
rect 8941 25647 8999 25653
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10962 25684 10968 25696
rect 9732 25656 10968 25684
rect 9732 25644 9738 25656
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 13817 25687 13875 25693
rect 13817 25684 13829 25687
rect 12860 25656 13829 25684
rect 12860 25644 12866 25656
rect 13817 25653 13829 25656
rect 13863 25653 13875 25687
rect 13817 25647 13875 25653
rect 14277 25687 14335 25693
rect 14277 25653 14289 25687
rect 14323 25684 14335 25687
rect 14458 25684 14464 25696
rect 14323 25656 14464 25684
rect 14323 25653 14335 25656
rect 14277 25647 14335 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 16298 25644 16304 25696
rect 16356 25644 16362 25696
rect 18969 25687 19027 25693
rect 18969 25653 18981 25687
rect 19015 25684 19027 25687
rect 19334 25684 19340 25696
rect 19015 25656 19340 25684
rect 19015 25653 19027 25656
rect 18969 25647 19027 25653
rect 19334 25644 19340 25656
rect 19392 25644 19398 25696
rect 19444 25684 19472 25724
rect 20257 25721 20269 25755
rect 20303 25721 20315 25755
rect 20257 25715 20315 25721
rect 21468 25684 21496 25860
rect 22738 25848 22744 25900
rect 22796 25888 22802 25900
rect 22796 25860 23060 25888
rect 22796 25848 22802 25860
rect 21542 25780 21548 25832
rect 21600 25820 21606 25832
rect 22005 25823 22063 25829
rect 22005 25820 22017 25823
rect 21600 25792 22017 25820
rect 21600 25780 21606 25792
rect 22005 25789 22017 25792
rect 22051 25789 22063 25823
rect 23032 25820 23060 25860
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 24101 25891 24159 25897
rect 24101 25888 24113 25891
rect 23532 25860 24113 25888
rect 23532 25848 23538 25860
rect 24101 25857 24113 25860
rect 24147 25857 24159 25891
rect 24101 25851 24159 25857
rect 25682 25848 25688 25900
rect 25740 25848 25746 25900
rect 23845 25823 23903 25829
rect 23845 25820 23857 25823
rect 23032 25792 23857 25820
rect 22005 25783 22063 25789
rect 23845 25789 23857 25792
rect 23891 25789 23903 25823
rect 23845 25783 23903 25789
rect 22020 25696 22048 25783
rect 19444 25656 21496 25684
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 22370 25684 22376 25696
rect 22060 25656 22376 25684
rect 22060 25644 22066 25656
rect 22370 25644 22376 25656
rect 22428 25644 22434 25696
rect 22738 25644 22744 25696
rect 22796 25684 22802 25696
rect 23385 25687 23443 25693
rect 23385 25684 23397 25687
rect 22796 25656 23397 25684
rect 22796 25644 22802 25656
rect 23385 25653 23397 25656
rect 23431 25653 23443 25687
rect 23860 25684 23888 25783
rect 25866 25712 25872 25764
rect 25924 25712 25930 25764
rect 24578 25684 24584 25696
rect 23860 25656 24584 25684
rect 23385 25647 23443 25653
rect 24578 25644 24584 25656
rect 24636 25644 24642 25696
rect 24946 25644 24952 25696
rect 25004 25684 25010 25696
rect 25225 25687 25283 25693
rect 25225 25684 25237 25687
rect 25004 25656 25237 25684
rect 25004 25644 25010 25656
rect 25225 25653 25237 25656
rect 25271 25653 25283 25687
rect 25225 25647 25283 25653
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 3329 25483 3387 25489
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 7466 25480 7472 25492
rect 3375 25452 7472 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 7466 25440 7472 25452
rect 7524 25440 7530 25492
rect 8202 25440 8208 25492
rect 8260 25480 8266 25492
rect 8389 25483 8447 25489
rect 8389 25480 8401 25483
rect 8260 25452 8401 25480
rect 8260 25440 8266 25452
rect 8389 25449 8401 25452
rect 8435 25480 8447 25483
rect 8754 25480 8760 25492
rect 8435 25452 8760 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 9861 25483 9919 25489
rect 9861 25449 9873 25483
rect 9907 25480 9919 25483
rect 10594 25480 10600 25492
rect 9907 25452 10600 25480
rect 9907 25449 9919 25452
rect 9861 25443 9919 25449
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 13078 25480 13084 25492
rect 12584 25452 13084 25480
rect 12584 25440 12590 25452
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 15010 25440 15016 25492
rect 15068 25440 15074 25492
rect 17862 25440 17868 25492
rect 17920 25440 17926 25492
rect 19242 25440 19248 25492
rect 19300 25480 19306 25492
rect 19300 25440 19334 25480
rect 19794 25440 19800 25492
rect 19852 25440 19858 25492
rect 20257 25483 20315 25489
rect 20257 25449 20269 25483
rect 20303 25480 20315 25483
rect 20898 25480 20904 25492
rect 20303 25452 20904 25480
rect 20303 25449 20315 25452
rect 20257 25443 20315 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 21177 25483 21235 25489
rect 21177 25449 21189 25483
rect 21223 25480 21235 25483
rect 21223 25452 21956 25480
rect 21223 25449 21235 25452
rect 21177 25443 21235 25449
rect 5534 25372 5540 25424
rect 5592 25412 5598 25424
rect 5997 25415 6055 25421
rect 5997 25412 6009 25415
rect 5592 25384 6009 25412
rect 5592 25372 5598 25384
rect 5997 25381 6009 25384
rect 6043 25381 6055 25415
rect 6822 25412 6828 25424
rect 5997 25375 6055 25381
rect 6288 25384 6828 25412
rect 5902 25304 5908 25356
rect 5960 25344 5966 25356
rect 5960 25316 6224 25344
rect 5960 25304 5966 25316
rect 1946 25236 1952 25288
rect 2004 25236 2010 25288
rect 2038 25236 2044 25288
rect 2096 25276 2102 25288
rect 2205 25279 2263 25285
rect 2205 25276 2217 25279
rect 2096 25248 2217 25276
rect 2096 25236 2102 25248
rect 2205 25245 2217 25248
rect 2251 25245 2263 25279
rect 2205 25239 2263 25245
rect 2498 25236 2504 25288
rect 2556 25276 2562 25288
rect 6196 25285 6224 25316
rect 6288 25285 6316 25384
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 10410 25412 10416 25424
rect 10336 25384 10416 25412
rect 6362 25304 6368 25356
rect 6420 25344 6426 25356
rect 8021 25347 8079 25353
rect 8021 25344 8033 25347
rect 6420 25316 8033 25344
rect 6420 25304 6426 25316
rect 8021 25313 8033 25316
rect 8067 25344 8079 25347
rect 8570 25344 8576 25356
rect 8067 25316 8576 25344
rect 8067 25313 8079 25316
rect 8021 25307 8079 25313
rect 8570 25304 8576 25316
rect 8628 25344 8634 25356
rect 9766 25344 9772 25356
rect 8628 25316 9772 25344
rect 8628 25304 8634 25316
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 10336 25344 10364 25384
rect 10410 25372 10416 25384
rect 10468 25372 10474 25424
rect 10962 25412 10968 25424
rect 10520 25384 10968 25412
rect 10520 25353 10548 25384
rect 10962 25372 10968 25384
rect 11020 25372 11026 25424
rect 13814 25372 13820 25424
rect 13872 25412 13878 25424
rect 16022 25412 16028 25424
rect 13872 25384 16028 25412
rect 13872 25372 13878 25384
rect 16022 25372 16028 25384
rect 16080 25372 16086 25424
rect 16114 25372 16120 25424
rect 16172 25412 16178 25424
rect 18693 25415 18751 25421
rect 18693 25412 18705 25415
rect 16172 25384 18705 25412
rect 16172 25372 16178 25384
rect 18693 25381 18705 25384
rect 18739 25381 18751 25415
rect 19306 25412 19334 25440
rect 21266 25412 21272 25424
rect 19306 25384 21272 25412
rect 18693 25375 18751 25381
rect 21266 25372 21272 25384
rect 21324 25372 21330 25424
rect 21928 25412 21956 25452
rect 22002 25440 22008 25492
rect 22060 25440 22066 25492
rect 22554 25440 22560 25492
rect 22612 25480 22618 25492
rect 22741 25483 22799 25489
rect 22741 25480 22753 25483
rect 22612 25452 22753 25480
rect 22612 25440 22618 25452
rect 22741 25449 22753 25452
rect 22787 25480 22799 25483
rect 23198 25480 23204 25492
rect 22787 25452 23204 25480
rect 22787 25449 22799 25452
rect 22741 25443 22799 25449
rect 23198 25440 23204 25452
rect 23256 25440 23262 25492
rect 23293 25483 23351 25489
rect 23293 25449 23305 25483
rect 23339 25480 23351 25483
rect 24118 25480 24124 25492
rect 23339 25452 24124 25480
rect 23339 25449 23351 25452
rect 23293 25443 23351 25449
rect 24118 25440 24124 25452
rect 24176 25440 24182 25492
rect 25682 25440 25688 25492
rect 25740 25480 25746 25492
rect 27614 25480 27620 25492
rect 25740 25452 27620 25480
rect 25740 25440 25746 25452
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 24762 25412 24768 25424
rect 21928 25384 24768 25412
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 9968 25316 10364 25344
rect 10505 25347 10563 25353
rect 3973 25279 4031 25285
rect 3973 25276 3985 25279
rect 2556 25248 3985 25276
rect 2556 25236 2562 25248
rect 3973 25245 3985 25248
rect 4019 25245 4031 25279
rect 3973 25239 4031 25245
rect 6181 25279 6239 25285
rect 6181 25245 6193 25279
rect 6227 25245 6239 25279
rect 6181 25239 6239 25245
rect 6273 25279 6331 25285
rect 6273 25245 6285 25279
rect 6319 25245 6331 25279
rect 6273 25239 6331 25245
rect 6454 25236 6460 25288
rect 6512 25286 6518 25288
rect 6512 25285 6526 25286
rect 6512 25279 6541 25285
rect 6529 25245 6541 25279
rect 6512 25239 6541 25245
rect 6641 25279 6699 25285
rect 6641 25245 6653 25279
rect 6687 25276 6699 25279
rect 6730 25276 6736 25288
rect 6687 25248 6736 25276
rect 6687 25245 6699 25248
rect 6641 25239 6699 25245
rect 6512 25236 6518 25239
rect 6730 25236 6736 25248
rect 6788 25236 6794 25288
rect 7193 25279 7251 25285
rect 7193 25245 7205 25279
rect 7239 25276 7251 25279
rect 7926 25276 7932 25288
rect 7239 25248 7932 25276
rect 7239 25245 7251 25248
rect 7193 25239 7251 25245
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 9214 25236 9220 25288
rect 9272 25236 9278 25288
rect 9401 25279 9459 25285
rect 9401 25245 9413 25279
rect 9447 25276 9459 25279
rect 9490 25276 9496 25288
rect 9447 25248 9496 25276
rect 9447 25245 9459 25248
rect 9401 25239 9459 25245
rect 9490 25236 9496 25248
rect 9548 25276 9554 25288
rect 9968 25276 9996 25316
rect 10505 25313 10517 25347
rect 10551 25313 10563 25347
rect 10505 25307 10563 25313
rect 13633 25347 13691 25353
rect 13633 25313 13645 25347
rect 13679 25344 13691 25347
rect 18046 25344 18052 25356
rect 13679 25316 18052 25344
rect 13679 25313 13691 25316
rect 13633 25307 13691 25313
rect 18046 25304 18052 25316
rect 18104 25304 18110 25356
rect 19242 25344 19248 25356
rect 18156 25316 18552 25344
rect 9548 25248 9996 25276
rect 9548 25236 9554 25248
rect 10042 25236 10048 25288
rect 10100 25276 10106 25288
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 10100 25248 11437 25276
rect 10100 25236 10106 25248
rect 11425 25245 11437 25248
rect 11471 25276 11483 25279
rect 12434 25276 12440 25288
rect 11471 25248 12440 25276
rect 11471 25245 11483 25248
rect 11425 25239 11483 25245
rect 12434 25236 12440 25248
rect 12492 25276 12498 25288
rect 12618 25276 12624 25288
rect 12492 25248 12624 25276
rect 12492 25236 12498 25248
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25276 13507 25279
rect 13998 25276 14004 25288
rect 13495 25248 14004 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 13998 25236 14004 25248
rect 14056 25276 14062 25288
rect 14182 25276 14188 25288
rect 14056 25248 14188 25276
rect 14056 25236 14062 25248
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 15378 25276 15384 25288
rect 14292 25248 15384 25276
rect 1854 25168 1860 25220
rect 1912 25208 1918 25220
rect 4218 25211 4276 25217
rect 4218 25208 4230 25211
rect 1912 25180 4230 25208
rect 1912 25168 1918 25180
rect 4218 25177 4230 25180
rect 4264 25177 4276 25211
rect 4218 25171 4276 25177
rect 6365 25211 6423 25217
rect 6365 25177 6377 25211
rect 6411 25177 6423 25211
rect 6365 25171 6423 25177
rect 5350 25100 5356 25152
rect 5408 25100 5414 25152
rect 6380 25140 6408 25171
rect 7282 25168 7288 25220
rect 7340 25208 7346 25220
rect 7561 25211 7619 25217
rect 7561 25208 7573 25211
rect 7340 25180 7573 25208
rect 7340 25168 7346 25180
rect 7561 25177 7573 25180
rect 7607 25177 7619 25211
rect 7561 25171 7619 25177
rect 7834 25168 7840 25220
rect 7892 25208 7898 25220
rect 7892 25180 8708 25208
rect 7892 25168 7898 25180
rect 6546 25140 6552 25152
rect 6380 25112 6552 25140
rect 6546 25100 6552 25112
rect 6604 25140 6610 25152
rect 6822 25140 6828 25152
rect 6604 25112 6828 25140
rect 6604 25100 6610 25112
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 6914 25100 6920 25152
rect 6972 25140 6978 25152
rect 8202 25140 8208 25152
rect 6972 25112 8208 25140
rect 6972 25100 6978 25112
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 8386 25100 8392 25152
rect 8444 25100 8450 25152
rect 8478 25100 8484 25152
rect 8536 25140 8542 25152
rect 8573 25143 8631 25149
rect 8573 25140 8585 25143
rect 8536 25112 8585 25140
rect 8536 25100 8542 25112
rect 8573 25109 8585 25112
rect 8619 25109 8631 25143
rect 8680 25140 8708 25180
rect 8754 25168 8760 25220
rect 8812 25208 8818 25220
rect 9674 25208 9680 25220
rect 8812 25180 9680 25208
rect 8812 25168 8818 25180
rect 9674 25168 9680 25180
rect 9732 25208 9738 25220
rect 10321 25211 10379 25217
rect 10321 25208 10333 25211
rect 9732 25180 10333 25208
rect 9732 25168 9738 25180
rect 10321 25177 10333 25180
rect 10367 25208 10379 25211
rect 10962 25208 10968 25220
rect 10367 25180 10968 25208
rect 10367 25177 10379 25180
rect 10321 25171 10379 25177
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 11054 25168 11060 25220
rect 11112 25208 11118 25220
rect 11670 25211 11728 25217
rect 11670 25208 11682 25211
rect 11112 25180 11682 25208
rect 11112 25168 11118 25180
rect 11670 25177 11682 25180
rect 11716 25177 11728 25211
rect 11670 25171 11728 25177
rect 13265 25211 13323 25217
rect 13265 25177 13277 25211
rect 13311 25177 13323 25211
rect 13265 25171 13323 25177
rect 10229 25143 10287 25149
rect 10229 25140 10241 25143
rect 8680 25112 10241 25140
rect 8573 25103 8631 25109
rect 10229 25109 10241 25112
rect 10275 25140 10287 25143
rect 10410 25140 10416 25152
rect 10275 25112 10416 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 10502 25100 10508 25152
rect 10560 25140 10566 25152
rect 12434 25140 12440 25152
rect 10560 25112 12440 25140
rect 10560 25100 10566 25112
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 12805 25143 12863 25149
rect 12805 25109 12817 25143
rect 12851 25140 12863 25143
rect 13170 25140 13176 25152
rect 12851 25112 13176 25140
rect 12851 25109 12863 25112
rect 12805 25103 12863 25109
rect 13170 25100 13176 25112
rect 13228 25100 13234 25152
rect 13280 25140 13308 25171
rect 13722 25168 13728 25220
rect 13780 25208 13786 25220
rect 14292 25208 14320 25248
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 15838 25236 15844 25288
rect 15896 25236 15902 25288
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16850 25276 16856 25288
rect 16163 25248 16856 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16850 25236 16856 25248
rect 16908 25276 16914 25288
rect 16908 25248 17816 25276
rect 16908 25236 16914 25248
rect 13780 25180 14320 25208
rect 14829 25211 14887 25217
rect 13780 25168 13786 25180
rect 14829 25177 14841 25211
rect 14875 25208 14887 25211
rect 15286 25208 15292 25220
rect 14875 25180 15292 25208
rect 14875 25177 14887 25180
rect 14829 25171 14887 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 15396 25208 15424 25236
rect 17497 25211 17555 25217
rect 17497 25208 17509 25211
rect 15396 25180 17509 25208
rect 17497 25177 17509 25180
rect 17543 25177 17555 25211
rect 17497 25171 17555 25177
rect 17678 25168 17684 25220
rect 17736 25168 17742 25220
rect 14090 25140 14096 25152
rect 13280 25112 14096 25140
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14182 25100 14188 25152
rect 14240 25140 14246 25152
rect 15029 25143 15087 25149
rect 15029 25140 15041 25143
rect 14240 25112 15041 25140
rect 14240 25100 14246 25112
rect 15029 25109 15041 25112
rect 15075 25109 15087 25143
rect 15029 25103 15087 25109
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 16482 25140 16488 25152
rect 15243 25112 16488 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 17218 25100 17224 25152
rect 17276 25140 17282 25152
rect 17696 25140 17724 25168
rect 17276 25112 17724 25140
rect 17788 25140 17816 25248
rect 18046 25168 18052 25220
rect 18104 25208 18110 25220
rect 18156 25208 18184 25316
rect 18524 25285 18552 25316
rect 18892 25316 19248 25344
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 18104 25180 18184 25208
rect 18432 25208 18460 25239
rect 18892 25208 18920 25316
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 20622 25304 20628 25356
rect 20680 25344 20686 25356
rect 20680 25316 23520 25344
rect 20680 25304 20686 25316
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 19392 25248 20453 25276
rect 19392 25236 19398 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 21082 25236 21088 25288
rect 21140 25276 21146 25288
rect 21361 25279 21419 25285
rect 21361 25276 21373 25279
rect 21140 25248 21373 25276
rect 21140 25236 21146 25248
rect 21361 25245 21373 25248
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 21913 25279 21971 25285
rect 21913 25245 21925 25279
rect 21959 25276 21971 25279
rect 22462 25276 22468 25288
rect 21959 25248 22468 25276
rect 21959 25245 21971 25248
rect 21913 25239 21971 25245
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 23492 25285 23520 25316
rect 22557 25279 22615 25285
rect 22557 25245 22569 25279
rect 22603 25245 22615 25279
rect 22557 25239 22615 25245
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25245 23535 25279
rect 23477 25239 23535 25245
rect 18432 25180 18920 25208
rect 18104 25168 18110 25180
rect 18966 25168 18972 25220
rect 19024 25208 19030 25220
rect 19429 25211 19487 25217
rect 19429 25208 19441 25211
rect 19024 25180 19441 25208
rect 19024 25168 19030 25180
rect 19429 25177 19441 25180
rect 19475 25177 19487 25211
rect 19429 25171 19487 25177
rect 19613 25211 19671 25217
rect 19613 25177 19625 25211
rect 19659 25208 19671 25211
rect 19886 25208 19892 25220
rect 19659 25180 19892 25208
rect 19659 25177 19671 25180
rect 19613 25171 19671 25177
rect 19886 25168 19892 25180
rect 19944 25168 19950 25220
rect 22572 25208 22600 25239
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25245 24823 25279
rect 24765 25239 24823 25245
rect 22066 25180 23520 25208
rect 22066 25140 22094 25180
rect 17788 25112 22094 25140
rect 23492 25140 23520 25180
rect 23566 25168 23572 25220
rect 23624 25208 23630 25220
rect 24780 25208 24808 25239
rect 26050 25236 26056 25288
rect 26108 25236 26114 25288
rect 23624 25180 24808 25208
rect 26320 25211 26378 25217
rect 23624 25168 23630 25180
rect 26320 25177 26332 25211
rect 26366 25208 26378 25211
rect 26418 25208 26424 25220
rect 26366 25180 26424 25208
rect 26366 25177 26378 25180
rect 26320 25171 26378 25177
rect 26418 25168 26424 25180
rect 26476 25168 26482 25220
rect 23658 25140 23664 25152
rect 23492 25112 23664 25140
rect 17276 25100 17282 25112
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 24670 25100 24676 25152
rect 24728 25100 24734 25152
rect 27430 25100 27436 25152
rect 27488 25100 27494 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 1854 24896 1860 24948
rect 1912 24896 1918 24948
rect 5077 24939 5135 24945
rect 5077 24905 5089 24939
rect 5123 24936 5135 24939
rect 5258 24936 5264 24948
rect 5123 24908 5264 24936
rect 5123 24905 5135 24908
rect 5077 24899 5135 24905
rect 5258 24896 5264 24908
rect 5316 24936 5322 24948
rect 6086 24936 6092 24948
rect 5316 24908 6092 24936
rect 5316 24896 5322 24908
rect 6086 24896 6092 24908
rect 6144 24896 6150 24948
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 6917 24939 6975 24945
rect 6917 24936 6929 24939
rect 6512 24908 6929 24936
rect 6512 24896 6518 24908
rect 6917 24905 6929 24908
rect 6963 24905 6975 24939
rect 6917 24899 6975 24905
rect 2958 24828 2964 24880
rect 3016 24868 3022 24880
rect 5169 24871 5227 24877
rect 5169 24868 5181 24871
rect 3016 24840 4200 24868
rect 3016 24828 3022 24840
rect 1394 24760 1400 24812
rect 1452 24800 1458 24812
rect 1581 24803 1639 24809
rect 1581 24800 1593 24803
rect 1452 24772 1593 24800
rect 1452 24760 1458 24772
rect 1581 24769 1593 24772
rect 1627 24769 1639 24803
rect 1581 24763 1639 24769
rect 1854 24760 1860 24812
rect 1912 24760 1918 24812
rect 2860 24803 2918 24809
rect 2860 24769 2872 24803
rect 2906 24800 2918 24803
rect 4062 24800 4068 24812
rect 2906 24772 4068 24800
rect 2906 24769 2918 24772
rect 2860 24763 2918 24769
rect 4062 24760 4068 24772
rect 4120 24760 4126 24812
rect 4172 24800 4200 24840
rect 4816 24840 5181 24868
rect 4816 24800 4844 24840
rect 5169 24837 5181 24840
rect 5215 24837 5227 24871
rect 5169 24831 5227 24837
rect 5442 24828 5448 24880
rect 5500 24868 5506 24880
rect 5500 24840 5764 24868
rect 5500 24828 5506 24840
rect 4172 24772 4844 24800
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5350 24800 5356 24812
rect 4939 24772 5356 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 5736 24809 5764 24840
rect 5994 24828 6000 24880
rect 6052 24828 6058 24880
rect 6362 24828 6368 24880
rect 6420 24868 6426 24880
rect 6546 24868 6552 24880
rect 6420 24840 6552 24868
rect 6420 24828 6426 24840
rect 6546 24828 6552 24840
rect 6604 24828 6610 24880
rect 6932 24868 6960 24899
rect 7374 24896 7380 24948
rect 7432 24936 7438 24948
rect 7834 24936 7840 24948
rect 7432 24908 7840 24936
rect 7432 24896 7438 24908
rect 7834 24896 7840 24908
rect 7892 24896 7898 24948
rect 8754 24936 8760 24948
rect 7944 24908 8760 24936
rect 7944 24868 7972 24908
rect 8754 24896 8760 24908
rect 8812 24896 8818 24948
rect 9217 24939 9275 24945
rect 9217 24905 9229 24939
rect 9263 24936 9275 24939
rect 9306 24936 9312 24948
rect 9263 24908 9312 24936
rect 9263 24905 9275 24908
rect 9217 24899 9275 24905
rect 9306 24896 9312 24908
rect 9364 24896 9370 24948
rect 10410 24896 10416 24948
rect 10468 24896 10474 24948
rect 10778 24896 10784 24948
rect 10836 24936 10842 24948
rect 11149 24939 11207 24945
rect 11149 24936 11161 24939
rect 10836 24908 11161 24936
rect 10836 24896 10842 24908
rect 11149 24905 11161 24908
rect 11195 24905 11207 24939
rect 11149 24899 11207 24905
rect 11330 24896 11336 24948
rect 11388 24936 11394 24948
rect 12158 24936 12164 24948
rect 11388 24908 12164 24936
rect 11388 24896 11394 24908
rect 12158 24896 12164 24908
rect 12216 24896 12222 24948
rect 12434 24896 12440 24948
rect 12492 24936 12498 24948
rect 19889 24939 19947 24945
rect 12492 24908 17816 24936
rect 12492 24896 12498 24908
rect 8478 24868 8484 24880
rect 6779 24837 6837 24843
rect 6932 24840 7972 24868
rect 8312 24840 8484 24868
rect 6779 24834 6791 24837
rect 5721 24803 5779 24809
rect 5721 24769 5733 24803
rect 5767 24769 5779 24803
rect 5721 24763 5779 24769
rect 5810 24760 5816 24812
rect 5868 24760 5874 24812
rect 6012 24800 6040 24828
rect 6764 24803 6791 24834
rect 6825 24803 6837 24837
rect 6764 24800 6837 24803
rect 6914 24800 6920 24812
rect 6012 24772 6920 24800
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24800 7619 24803
rect 8312 24800 8340 24840
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 8573 24871 8631 24877
rect 8573 24837 8585 24871
rect 8619 24868 8631 24871
rect 8846 24868 8852 24880
rect 8619 24840 8852 24868
rect 8619 24837 8631 24840
rect 8573 24831 8631 24837
rect 8846 24828 8852 24840
rect 8904 24828 8910 24880
rect 10428 24868 10456 24896
rect 11054 24868 11060 24880
rect 9324 24840 9674 24868
rect 10428 24840 11060 24868
rect 9324 24812 9352 24840
rect 7607 24772 8340 24800
rect 8389 24803 8447 24809
rect 7607 24769 7619 24772
rect 7561 24763 7619 24769
rect 8389 24769 8401 24803
rect 8435 24800 8447 24803
rect 8435 24772 8708 24800
rect 8435 24769 8447 24772
rect 8389 24763 8447 24769
rect 2038 24692 2044 24744
rect 2096 24732 2102 24744
rect 2498 24732 2504 24744
rect 2096 24704 2504 24732
rect 2096 24692 2102 24704
rect 2498 24692 2504 24704
rect 2556 24732 2562 24744
rect 2593 24735 2651 24741
rect 2593 24732 2605 24735
rect 2556 24704 2605 24732
rect 2556 24692 2562 24704
rect 2593 24701 2605 24704
rect 2639 24701 2651 24735
rect 5997 24735 6055 24741
rect 5997 24732 6009 24735
rect 2593 24695 2651 24701
rect 3620 24704 6009 24732
rect 3326 24556 3332 24608
rect 3384 24596 3390 24608
rect 3620 24596 3648 24704
rect 5997 24701 6009 24704
rect 6043 24732 6055 24735
rect 7282 24732 7288 24744
rect 6043 24704 7288 24732
rect 6043 24701 6055 24704
rect 5997 24695 6055 24701
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 7374 24692 7380 24744
rect 7432 24732 7438 24744
rect 8404 24732 8432 24763
rect 7432 24704 8432 24732
rect 8680 24732 8708 24772
rect 9306 24760 9312 24812
rect 9364 24760 9370 24812
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 9490 24800 9496 24812
rect 9447 24772 9496 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 9646 24800 9674 24840
rect 11054 24828 11060 24840
rect 11112 24868 11118 24880
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 11112 24840 12081 24868
rect 11112 24828 11118 24840
rect 12069 24837 12081 24840
rect 12115 24837 12127 24871
rect 12894 24868 12900 24880
rect 12069 24831 12127 24837
rect 12544 24840 12900 24868
rect 9861 24803 9919 24809
rect 9861 24800 9873 24803
rect 9646 24772 9873 24800
rect 9861 24769 9873 24772
rect 9907 24800 9919 24803
rect 10321 24803 10379 24809
rect 9907 24772 10288 24800
rect 9907 24769 9919 24772
rect 9861 24763 9919 24769
rect 10042 24732 10048 24744
rect 8680 24704 10048 24732
rect 7432 24692 7438 24704
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 10260 24732 10288 24772
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 10502 24800 10508 24812
rect 10367 24772 10508 24800
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 10502 24760 10508 24772
rect 10560 24760 10566 24812
rect 10594 24760 10600 24812
rect 10652 24760 10658 24812
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 11020 24772 12173 24800
rect 11020 24760 11026 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12544 24800 12572 24840
rect 12894 24828 12900 24840
rect 12952 24828 12958 24880
rect 15286 24828 15292 24880
rect 15344 24868 15350 24880
rect 17405 24871 17463 24877
rect 17405 24868 17417 24871
rect 15344 24840 17417 24868
rect 15344 24828 15350 24840
rect 17405 24837 17417 24840
rect 17451 24837 17463 24871
rect 17788 24868 17816 24908
rect 19889 24905 19901 24939
rect 19935 24936 19947 24939
rect 20070 24936 20076 24948
rect 19935 24908 20076 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 20070 24896 20076 24908
rect 20128 24896 20134 24948
rect 23382 24896 23388 24948
rect 23440 24936 23446 24948
rect 26602 24936 26608 24948
rect 23440 24908 26608 24936
rect 23440 24896 23446 24908
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 24578 24868 24584 24880
rect 17405 24831 17463 24837
rect 17635 24837 17693 24843
rect 17788 24840 24584 24868
rect 17635 24834 17647 24837
rect 12161 24763 12219 24769
rect 12360 24772 12572 24800
rect 10778 24732 10784 24744
rect 10260 24704 10784 24732
rect 10778 24692 10784 24704
rect 10836 24692 10842 24744
rect 12360 24741 12388 24772
rect 12618 24760 12624 24812
rect 12676 24800 12682 24812
rect 13449 24803 13507 24809
rect 13449 24800 13461 24803
rect 12676 24772 13461 24800
rect 12676 24760 12682 24772
rect 13449 24769 13461 24772
rect 13495 24769 13507 24803
rect 13449 24763 13507 24769
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 13705 24803 13763 24809
rect 13705 24800 13717 24803
rect 13596 24772 13717 24800
rect 13596 24760 13602 24772
rect 13705 24769 13717 24772
rect 13751 24769 13763 24803
rect 13705 24763 13763 24769
rect 15654 24760 15660 24812
rect 15712 24760 15718 24812
rect 15746 24760 15752 24812
rect 15804 24800 15810 24812
rect 15804 24772 15849 24800
rect 15804 24760 15810 24772
rect 15930 24760 15936 24812
rect 15988 24760 15994 24812
rect 16022 24760 16028 24812
rect 16080 24760 16086 24812
rect 16114 24760 16120 24812
rect 16172 24809 16178 24812
rect 16172 24800 16180 24809
rect 17620 24803 17647 24834
rect 17681 24812 17693 24837
rect 24578 24828 24584 24840
rect 24636 24828 24642 24880
rect 25038 24828 25044 24880
rect 25096 24868 25102 24880
rect 25470 24871 25528 24877
rect 25470 24868 25482 24871
rect 25096 24840 25482 24868
rect 25096 24828 25102 24840
rect 25470 24837 25482 24840
rect 25516 24837 25528 24871
rect 25470 24831 25528 24837
rect 25590 24828 25596 24880
rect 25648 24828 25654 24880
rect 17681 24803 17684 24812
rect 16172 24772 16217 24800
rect 17620 24772 17684 24803
rect 16172 24763 16180 24772
rect 16172 24760 16178 24763
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 19058 24800 19064 24812
rect 18616 24772 19064 24800
rect 12345 24735 12403 24741
rect 12345 24701 12357 24735
rect 12391 24701 12403 24735
rect 15948 24732 15976 24760
rect 16390 24732 16396 24744
rect 15948 24704 16396 24732
rect 12345 24695 12403 24701
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18233 24735 18291 24741
rect 18233 24732 18245 24735
rect 17828 24704 18245 24732
rect 17828 24692 17834 24704
rect 18233 24701 18245 24704
rect 18279 24701 18291 24735
rect 18233 24695 18291 24701
rect 3973 24667 4031 24673
rect 3973 24633 3985 24667
rect 4019 24664 4031 24667
rect 6362 24664 6368 24676
rect 4019 24636 6368 24664
rect 4019 24633 4031 24636
rect 3973 24627 4031 24633
rect 6362 24624 6368 24636
rect 6420 24624 6426 24676
rect 7837 24667 7895 24673
rect 7837 24633 7849 24667
rect 7883 24664 7895 24667
rect 7926 24664 7932 24676
rect 7883 24636 7932 24664
rect 7883 24633 7895 24636
rect 7837 24627 7895 24633
rect 7926 24624 7932 24636
rect 7984 24624 7990 24676
rect 8846 24624 8852 24676
rect 8904 24664 8910 24676
rect 12802 24664 12808 24676
rect 8904 24636 12808 24664
rect 8904 24624 8910 24636
rect 12802 24624 12808 24636
rect 12860 24624 12866 24676
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 16942 24664 16948 24676
rect 14608 24636 16948 24664
rect 14608 24624 14614 24636
rect 16942 24624 16948 24636
rect 17000 24624 17006 24676
rect 17954 24664 17960 24676
rect 17604 24636 17960 24664
rect 3384 24568 3648 24596
rect 3384 24556 3390 24568
rect 4062 24556 4068 24608
rect 4120 24596 4126 24608
rect 4617 24599 4675 24605
rect 4617 24596 4629 24599
rect 4120 24568 4629 24596
rect 4120 24556 4126 24568
rect 4617 24565 4629 24568
rect 4663 24565 4675 24599
rect 4617 24559 4675 24565
rect 4890 24556 4896 24608
rect 4948 24596 4954 24608
rect 5905 24599 5963 24605
rect 5905 24596 5917 24599
rect 4948 24568 5917 24596
rect 4948 24556 4954 24568
rect 5905 24565 5917 24568
rect 5951 24565 5963 24599
rect 5905 24559 5963 24565
rect 5994 24556 6000 24608
rect 6052 24596 6058 24608
rect 6733 24599 6791 24605
rect 6733 24596 6745 24599
rect 6052 24568 6745 24596
rect 6052 24556 6058 24568
rect 6733 24565 6745 24568
rect 6779 24596 6791 24599
rect 8662 24596 8668 24608
rect 6779 24568 8668 24596
rect 6779 24565 6791 24568
rect 6733 24559 6791 24565
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 8754 24556 8760 24608
rect 8812 24556 8818 24608
rect 9030 24556 9036 24608
rect 9088 24596 9094 24608
rect 11330 24596 11336 24608
rect 9088 24568 11336 24596
rect 9088 24556 9094 24568
rect 11330 24556 11336 24568
rect 11388 24556 11394 24608
rect 11514 24556 11520 24608
rect 11572 24596 11578 24608
rect 11701 24599 11759 24605
rect 11701 24596 11713 24599
rect 11572 24568 11713 24596
rect 11572 24556 11578 24568
rect 11701 24565 11713 24568
rect 11747 24565 11759 24599
rect 11701 24559 11759 24565
rect 12894 24556 12900 24608
rect 12952 24596 12958 24608
rect 14829 24599 14887 24605
rect 14829 24596 14841 24599
rect 12952 24568 14841 24596
rect 12952 24556 12958 24568
rect 14829 24565 14841 24568
rect 14875 24565 14887 24599
rect 14829 24559 14887 24565
rect 15562 24556 15568 24608
rect 15620 24596 15626 24608
rect 17604 24605 17632 24636
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 16301 24599 16359 24605
rect 16301 24596 16313 24599
rect 15620 24568 16313 24596
rect 15620 24556 15626 24568
rect 16301 24565 16313 24568
rect 16347 24565 16359 24599
rect 16301 24559 16359 24565
rect 17589 24599 17647 24605
rect 17589 24565 17601 24599
rect 17635 24565 17647 24599
rect 17589 24559 17647 24565
rect 17770 24556 17776 24608
rect 17828 24556 17834 24608
rect 18248 24596 18276 24695
rect 18616 24673 18644 24772
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 20533 24803 20591 24809
rect 20533 24800 20545 24803
rect 20128 24772 20545 24800
rect 20128 24760 20134 24772
rect 20533 24769 20545 24772
rect 20579 24769 20591 24803
rect 20533 24763 20591 24769
rect 21177 24803 21235 24809
rect 21177 24769 21189 24803
rect 21223 24800 21235 24803
rect 21358 24800 21364 24812
rect 21223 24772 21364 24800
rect 21223 24769 21235 24772
rect 21177 24763 21235 24769
rect 21358 24760 21364 24772
rect 21416 24760 21422 24812
rect 22261 24803 22319 24809
rect 22261 24800 22273 24803
rect 21468 24772 22273 24800
rect 18693 24735 18751 24741
rect 18693 24701 18705 24735
rect 18739 24732 18751 24735
rect 19334 24732 19340 24744
rect 18739 24704 19340 24732
rect 18739 24701 18751 24704
rect 18693 24695 18751 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 19429 24735 19487 24741
rect 19429 24701 19441 24735
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 18601 24667 18659 24673
rect 18601 24633 18613 24667
rect 18647 24633 18659 24667
rect 18601 24627 18659 24633
rect 18782 24624 18788 24676
rect 18840 24664 18846 24676
rect 19444 24664 19472 24695
rect 19518 24692 19524 24744
rect 19576 24732 19582 24744
rect 21468 24732 21496 24772
rect 22261 24769 22273 24772
rect 22307 24769 22319 24803
rect 22261 24763 22319 24769
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 24029 24803 24087 24809
rect 24029 24800 24041 24803
rect 23072 24772 24041 24800
rect 23072 24760 23078 24772
rect 24029 24769 24041 24772
rect 24075 24769 24087 24803
rect 24029 24763 24087 24769
rect 24673 24803 24731 24809
rect 24673 24769 24685 24803
rect 24719 24769 24731 24803
rect 24673 24763 24731 24769
rect 25225 24803 25283 24809
rect 25225 24769 25237 24803
rect 25271 24800 25283 24803
rect 25608 24800 25636 24828
rect 25271 24772 25636 24800
rect 25271 24769 25283 24772
rect 25225 24763 25283 24769
rect 19576 24704 21496 24732
rect 19576 24692 19582 24704
rect 21542 24692 21548 24744
rect 21600 24732 21606 24744
rect 22002 24732 22008 24744
rect 21600 24704 22008 24732
rect 21600 24692 21606 24704
rect 22002 24692 22008 24704
rect 22060 24692 22066 24744
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 24688 24732 24716 24763
rect 23808 24704 24716 24732
rect 23808 24692 23814 24704
rect 18840 24636 19564 24664
rect 18840 24624 18846 24636
rect 18966 24596 18972 24608
rect 18248 24568 18972 24596
rect 18966 24556 18972 24568
rect 19024 24556 19030 24608
rect 19536 24596 19564 24636
rect 19610 24624 19616 24676
rect 19668 24664 19674 24676
rect 19705 24667 19763 24673
rect 19705 24664 19717 24667
rect 19668 24636 19717 24664
rect 19668 24624 19674 24636
rect 19705 24633 19717 24636
rect 19751 24633 19763 24667
rect 19705 24627 19763 24633
rect 20349 24667 20407 24673
rect 20349 24633 20361 24667
rect 20395 24664 20407 24667
rect 23474 24664 23480 24676
rect 20395 24636 21220 24664
rect 20395 24633 20407 24636
rect 20349 24627 20407 24633
rect 20898 24596 20904 24608
rect 19536 24568 20904 24596
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 20990 24556 20996 24608
rect 21048 24556 21054 24608
rect 21192 24596 21220 24636
rect 23124 24636 23480 24664
rect 23124 24596 23152 24636
rect 23474 24624 23480 24636
rect 23532 24624 23538 24676
rect 23845 24667 23903 24673
rect 23845 24633 23857 24667
rect 23891 24664 23903 24667
rect 24854 24664 24860 24676
rect 23891 24636 24860 24664
rect 23891 24633 23903 24636
rect 23845 24627 23903 24633
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 21192 24568 23152 24596
rect 23382 24556 23388 24608
rect 23440 24556 23446 24608
rect 24486 24556 24492 24608
rect 24544 24556 24550 24608
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 26605 24599 26663 24605
rect 26605 24596 26617 24599
rect 25924 24568 26617 24596
rect 25924 24556 25930 24568
rect 26605 24565 26617 24568
rect 26651 24565 26663 24599
rect 26605 24559 26663 24565
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 3510 24352 3516 24404
rect 3568 24392 3574 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 3568 24364 4077 24392
rect 3568 24352 3574 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4065 24355 4123 24361
rect 5442 24352 5448 24404
rect 5500 24392 5506 24404
rect 5626 24392 5632 24404
rect 5500 24364 5632 24392
rect 5500 24352 5506 24364
rect 5626 24352 5632 24364
rect 5684 24392 5690 24404
rect 6917 24395 6975 24401
rect 6917 24392 6929 24395
rect 5684 24364 6929 24392
rect 5684 24352 5690 24364
rect 6917 24361 6929 24364
rect 6963 24361 6975 24395
rect 6917 24355 6975 24361
rect 7650 24352 7656 24404
rect 7708 24392 7714 24404
rect 7745 24395 7803 24401
rect 7745 24392 7757 24395
rect 7708 24364 7757 24392
rect 7708 24352 7714 24364
rect 7745 24361 7757 24364
rect 7791 24361 7803 24395
rect 7745 24355 7803 24361
rect 7834 24352 7840 24404
rect 7892 24392 7898 24404
rect 8389 24395 8447 24401
rect 8389 24392 8401 24395
rect 7892 24364 8401 24392
rect 7892 24352 7898 24364
rect 8389 24361 8401 24364
rect 8435 24361 8447 24395
rect 8389 24355 8447 24361
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 9582 24392 9588 24404
rect 8628 24364 9588 24392
rect 8628 24352 8634 24364
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 10962 24392 10968 24404
rect 10704 24364 10968 24392
rect 5368 24296 7696 24324
rect 5368 24256 5396 24296
rect 7668 24268 7696 24296
rect 10502 24284 10508 24336
rect 10560 24284 10566 24336
rect 10594 24284 10600 24336
rect 10652 24324 10658 24336
rect 10704 24324 10732 24364
rect 10962 24352 10968 24364
rect 11020 24392 11026 24404
rect 17310 24392 17316 24404
rect 11020 24364 17316 24392
rect 11020 24352 11026 24364
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 17770 24352 17776 24404
rect 17828 24352 17834 24404
rect 18693 24395 18751 24401
rect 18693 24361 18705 24395
rect 18739 24392 18751 24395
rect 19518 24392 19524 24404
rect 18739 24364 19524 24392
rect 18739 24361 18751 24364
rect 18693 24355 18751 24361
rect 19518 24352 19524 24364
rect 19576 24352 19582 24404
rect 20441 24395 20499 24401
rect 19628 24364 20392 24392
rect 10652 24296 10732 24324
rect 11701 24327 11759 24333
rect 10652 24284 10658 24296
rect 11701 24293 11713 24327
rect 11747 24324 11759 24327
rect 13725 24327 13783 24333
rect 11747 24296 13216 24324
rect 11747 24293 11759 24296
rect 11701 24287 11759 24293
rect 5445 24259 5503 24265
rect 5445 24256 5457 24259
rect 5368 24228 5457 24256
rect 5445 24225 5457 24228
rect 5491 24225 5503 24259
rect 5902 24256 5908 24268
rect 5445 24219 5503 24225
rect 5690 24228 5908 24256
rect 2038 24148 2044 24200
rect 2096 24148 2102 24200
rect 2130 24148 2136 24200
rect 2188 24188 2194 24200
rect 2297 24191 2355 24197
rect 2297 24188 2309 24191
rect 2188 24160 2309 24188
rect 2188 24148 2194 24160
rect 2297 24157 2309 24160
rect 2343 24157 2355 24191
rect 2297 24151 2355 24157
rect 3878 24148 3884 24200
rect 3936 24188 3942 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 3936 24160 4629 24188
rect 3936 24148 3942 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 4706 24148 4712 24200
rect 4764 24188 4770 24200
rect 4982 24188 4988 24200
rect 4764 24160 4988 24188
rect 4764 24148 4770 24160
rect 4982 24148 4988 24160
rect 5040 24188 5046 24200
rect 5169 24191 5227 24197
rect 5169 24188 5181 24191
rect 5040 24160 5181 24188
rect 5040 24148 5046 24160
rect 5169 24157 5181 24160
rect 5215 24157 5227 24191
rect 5169 24151 5227 24157
rect 5258 24148 5264 24200
rect 5316 24186 5322 24200
rect 5353 24191 5411 24197
rect 5353 24186 5365 24191
rect 5316 24158 5365 24186
rect 5316 24148 5322 24158
rect 5353 24157 5365 24158
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5690 24197 5718 24228
rect 5902 24216 5908 24228
rect 5960 24216 5966 24268
rect 7650 24216 7656 24268
rect 7708 24216 7714 24268
rect 8846 24216 8852 24268
rect 8904 24256 8910 24268
rect 10520 24256 10548 24284
rect 8904 24228 10732 24256
rect 8904 24216 8910 24228
rect 5676 24191 5734 24197
rect 5676 24157 5688 24191
rect 5722 24157 5734 24191
rect 5676 24151 5734 24157
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 7561 24191 7619 24197
rect 7561 24157 7573 24191
rect 7607 24188 7619 24191
rect 9030 24188 9036 24200
rect 7607 24160 9036 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 9030 24148 9036 24160
rect 9088 24148 9094 24200
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 9180 24160 9229 24188
rect 9180 24148 9186 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9401 24191 9459 24197
rect 9401 24157 9413 24191
rect 9447 24188 9459 24191
rect 10413 24191 10471 24197
rect 9447 24160 10364 24188
rect 9447 24157 9459 24160
rect 9401 24151 9459 24157
rect 4338 24080 4344 24132
rect 4396 24080 4402 24132
rect 4525 24123 4583 24129
rect 4525 24089 4537 24123
rect 4571 24120 4583 24123
rect 5994 24120 6000 24132
rect 4571 24092 6000 24120
rect 4571 24089 4583 24092
rect 4525 24083 4583 24089
rect 5994 24080 6000 24092
rect 6052 24080 6058 24132
rect 6086 24080 6092 24132
rect 6144 24120 6150 24132
rect 6546 24120 6552 24132
rect 6144 24092 6552 24120
rect 6144 24080 6150 24092
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 6733 24123 6791 24129
rect 6733 24089 6745 24123
rect 6779 24089 6791 24123
rect 6733 24083 6791 24089
rect 3050 24012 3056 24064
rect 3108 24052 3114 24064
rect 3421 24055 3479 24061
rect 3421 24052 3433 24055
rect 3108 24024 3433 24052
rect 3108 24012 3114 24024
rect 3421 24021 3433 24024
rect 3467 24021 3479 24055
rect 3421 24015 3479 24021
rect 4798 24012 4804 24064
rect 4856 24052 4862 24064
rect 5905 24055 5963 24061
rect 5905 24052 5917 24055
rect 4856 24024 5917 24052
rect 4856 24012 4862 24024
rect 5905 24021 5917 24024
rect 5951 24021 5963 24055
rect 5905 24015 5963 24021
rect 6454 24012 6460 24064
rect 6512 24052 6518 24064
rect 6748 24052 6776 24083
rect 8294 24080 8300 24132
rect 8352 24080 8358 24132
rect 9582 24080 9588 24132
rect 9640 24080 9646 24132
rect 10336 24120 10364 24160
rect 10413 24157 10425 24191
rect 10459 24188 10471 24191
rect 10502 24188 10508 24200
rect 10459 24160 10508 24188
rect 10459 24157 10471 24160
rect 10413 24151 10471 24157
rect 10502 24148 10508 24160
rect 10560 24148 10566 24200
rect 10704 24197 10732 24228
rect 10689 24191 10747 24197
rect 10689 24157 10701 24191
rect 10735 24157 10747 24191
rect 10689 24151 10747 24157
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 11149 24191 11207 24197
rect 11149 24188 11161 24191
rect 10836 24160 11161 24188
rect 10836 24148 10842 24160
rect 11149 24157 11161 24160
rect 11195 24188 11207 24191
rect 11330 24188 11336 24200
rect 11195 24160 11336 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 11606 24120 11612 24132
rect 10336 24092 11612 24120
rect 11606 24080 11612 24092
rect 11664 24080 11670 24132
rect 8386 24052 8392 24064
rect 6512 24024 8392 24052
rect 6512 24012 6518 24024
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8478 24012 8484 24064
rect 8536 24052 8542 24064
rect 11716 24052 11744 24287
rect 12066 24216 12072 24268
rect 12124 24256 12130 24268
rect 13188 24256 13216 24296
rect 13725 24293 13737 24327
rect 13771 24324 13783 24327
rect 15194 24324 15200 24336
rect 13771 24296 15200 24324
rect 13771 24293 13783 24296
rect 13725 24287 13783 24293
rect 15194 24284 15200 24296
rect 15252 24284 15258 24336
rect 17402 24284 17408 24336
rect 17460 24324 17466 24336
rect 18230 24324 18236 24336
rect 17460 24296 18236 24324
rect 17460 24284 17466 24296
rect 18230 24284 18236 24296
rect 18288 24284 18294 24336
rect 18322 24284 18328 24336
rect 18380 24324 18386 24336
rect 18874 24324 18880 24336
rect 18380 24296 18880 24324
rect 18380 24284 18386 24296
rect 18874 24284 18880 24296
rect 18932 24284 18938 24336
rect 19058 24284 19064 24336
rect 19116 24324 19122 24336
rect 19628 24324 19656 24364
rect 19116 24296 19656 24324
rect 19116 24284 19122 24296
rect 19794 24284 19800 24336
rect 19852 24324 19858 24336
rect 20257 24327 20315 24333
rect 20257 24324 20269 24327
rect 19852 24296 20269 24324
rect 19852 24284 19858 24296
rect 20257 24293 20269 24296
rect 20303 24293 20315 24327
rect 20364 24324 20392 24364
rect 20441 24361 20453 24395
rect 20487 24392 20499 24395
rect 20622 24392 20628 24404
rect 20487 24364 20628 24392
rect 20487 24361 20499 24364
rect 20441 24355 20499 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 24946 24392 24952 24404
rect 20732 24364 24952 24392
rect 20732 24324 20760 24364
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 20364 24296 20760 24324
rect 20257 24287 20315 24293
rect 14645 24259 14703 24265
rect 12124 24228 12480 24256
rect 13188 24228 14412 24256
rect 12124 24216 12130 24228
rect 11882 24148 11888 24200
rect 11940 24188 11946 24200
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 11940 24160 12173 24188
rect 11940 24148 11946 24160
rect 12161 24157 12173 24160
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12452 24197 12480 24228
rect 12437 24191 12495 24197
rect 12308 24160 12353 24188
rect 12308 24148 12314 24160
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 12618 24148 12624 24200
rect 12676 24197 12682 24200
rect 12676 24188 12684 24197
rect 13541 24191 13599 24197
rect 12676 24160 12721 24188
rect 12676 24151 12684 24160
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13906 24188 13912 24200
rect 13587 24160 13912 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 12676 24148 12682 24151
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 12529 24123 12587 24129
rect 12529 24089 12541 24123
rect 12575 24089 12587 24123
rect 12529 24083 12587 24089
rect 8536 24024 11744 24052
rect 8536 24012 8542 24024
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 12544 24052 12572 24083
rect 13262 24080 13268 24132
rect 13320 24120 13326 24132
rect 13357 24123 13415 24129
rect 13357 24120 13369 24123
rect 13320 24092 13369 24120
rect 13320 24080 13326 24092
rect 13357 24089 13369 24092
rect 13403 24120 13415 24123
rect 13722 24120 13728 24132
rect 13403 24092 13728 24120
rect 13403 24089 13415 24092
rect 13357 24083 13415 24089
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 11848 24024 12572 24052
rect 12805 24055 12863 24061
rect 11848 24012 11854 24024
rect 12805 24021 12817 24055
rect 12851 24052 12863 24055
rect 14090 24052 14096 24064
rect 12851 24024 14096 24052
rect 12851 24021 12863 24024
rect 12805 24015 12863 24021
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14384 24052 14412 24228
rect 14645 24225 14657 24259
rect 14691 24256 14703 24259
rect 15378 24256 15384 24268
rect 14691 24228 15384 24256
rect 14691 24225 14703 24228
rect 14645 24219 14703 24225
rect 15378 24216 15384 24228
rect 15436 24216 15442 24268
rect 16942 24216 16948 24268
rect 17000 24256 17006 24268
rect 17000 24228 18368 24256
rect 17000 24216 17006 24228
rect 14550 24148 14556 24200
rect 14608 24148 14614 24200
rect 14734 24148 14740 24200
rect 14792 24148 14798 24200
rect 14826 24148 14832 24200
rect 14884 24148 14890 24200
rect 15010 24148 15016 24200
rect 15068 24148 15074 24200
rect 15657 24191 15715 24197
rect 15657 24157 15669 24191
rect 15703 24188 15715 24191
rect 16206 24188 16212 24200
rect 15703 24160 16212 24188
rect 15703 24157 15715 24160
rect 15657 24151 15715 24157
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 16482 24148 16488 24200
rect 16540 24188 16546 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 16540 24160 17877 24188
rect 16540 24148 16546 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 18138 24188 18144 24200
rect 18095 24160 18144 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18230 24148 18236 24200
rect 18288 24148 18294 24200
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 15902 24123 15960 24129
rect 15902 24120 15914 24123
rect 14516 24092 15914 24120
rect 14516 24080 14522 24092
rect 15902 24089 15914 24092
rect 15948 24089 15960 24123
rect 15902 24083 15960 24089
rect 16114 24080 16120 24132
rect 16172 24120 16178 24132
rect 17497 24123 17555 24129
rect 17497 24120 17509 24123
rect 16172 24092 17509 24120
rect 16172 24080 16178 24092
rect 17497 24089 17509 24092
rect 17543 24089 17555 24123
rect 18340 24120 18368 24228
rect 18966 24216 18972 24268
rect 19024 24256 19030 24268
rect 19426 24256 19432 24268
rect 19024 24228 19432 24256
rect 19024 24216 19030 24228
rect 19426 24216 19432 24228
rect 19484 24256 19490 24268
rect 19981 24259 20039 24265
rect 19981 24256 19993 24259
rect 19484 24228 19993 24256
rect 19484 24216 19490 24228
rect 19981 24225 19993 24228
rect 20027 24225 20039 24259
rect 19981 24219 20039 24225
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 20272 24188 20300 24287
rect 20990 24284 20996 24336
rect 21048 24324 21054 24336
rect 21269 24327 21327 24333
rect 21269 24324 21281 24327
rect 21048 24296 21281 24324
rect 21048 24284 21054 24296
rect 21269 24293 21281 24296
rect 21315 24324 21327 24327
rect 21450 24324 21456 24336
rect 21315 24296 21456 24324
rect 21315 24293 21327 24296
rect 21269 24287 21327 24293
rect 21450 24284 21456 24296
rect 21508 24284 21514 24336
rect 23658 24284 23664 24336
rect 23716 24284 23722 24336
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 21542 24256 21548 24268
rect 20956 24228 21548 24256
rect 20956 24216 20962 24228
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 22002 24216 22008 24268
rect 22060 24256 22066 24268
rect 22281 24259 22339 24265
rect 22281 24256 22293 24259
rect 22060 24228 22293 24256
rect 22060 24216 22066 24228
rect 22281 24225 22293 24228
rect 22327 24225 22339 24259
rect 22281 24219 22339 24225
rect 26050 24216 26056 24268
rect 26108 24256 26114 24268
rect 26421 24259 26479 24265
rect 26421 24256 26433 24259
rect 26108 24228 26433 24256
rect 26108 24216 26114 24228
rect 26421 24225 26433 24228
rect 26467 24225 26479 24259
rect 26421 24219 26479 24225
rect 22830 24188 22836 24200
rect 20272 24160 22836 24188
rect 22830 24148 22836 24160
rect 22888 24148 22894 24200
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 23348 24160 24593 24188
rect 23348 24148 23354 24160
rect 24581 24157 24593 24160
rect 24627 24188 24639 24191
rect 25130 24188 25136 24200
rect 24627 24160 25136 24188
rect 24627 24157 24639 24160
rect 24581 24151 24639 24157
rect 25130 24148 25136 24160
rect 25188 24188 25194 24200
rect 26068 24188 26096 24216
rect 26510 24188 26516 24200
rect 25188 24160 26096 24188
rect 26160 24160 26516 24188
rect 25188 24148 25194 24160
rect 18340 24092 19334 24120
rect 17497 24083 17555 24089
rect 16942 24052 16948 24064
rect 14384 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17037 24055 17095 24061
rect 17037 24021 17049 24055
rect 17083 24052 17095 24055
rect 17402 24052 17408 24064
rect 17083 24024 17408 24052
rect 17083 24021 17095 24024
rect 17037 24015 17095 24021
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 19306 24052 19334 24092
rect 19518 24080 19524 24132
rect 19576 24120 19582 24132
rect 22370 24120 22376 24132
rect 19576 24092 22376 24120
rect 19576 24080 19582 24092
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 22554 24129 22560 24132
rect 22548 24083 22560 24129
rect 22554 24080 22560 24083
rect 22612 24080 22618 24132
rect 23198 24080 23204 24132
rect 23256 24120 23262 24132
rect 23934 24120 23940 24132
rect 23256 24092 23940 24120
rect 23256 24080 23262 24092
rect 23934 24080 23940 24092
rect 23992 24080 23998 24132
rect 24854 24129 24860 24132
rect 24848 24083 24860 24129
rect 24854 24080 24860 24083
rect 24912 24080 24918 24132
rect 26160 24120 26188 24160
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 24964 24092 26188 24120
rect 21266 24052 21272 24064
rect 19306 24024 21272 24052
rect 21266 24012 21272 24024
rect 21324 24012 21330 24064
rect 21358 24012 21364 24064
rect 21416 24012 21422 24064
rect 23106 24012 23112 24064
rect 23164 24052 23170 24064
rect 24964 24052 24992 24092
rect 26234 24080 26240 24132
rect 26292 24120 26298 24132
rect 26666 24123 26724 24129
rect 26666 24120 26678 24123
rect 26292 24092 26678 24120
rect 26292 24080 26298 24092
rect 26666 24089 26678 24092
rect 26712 24089 26724 24123
rect 26666 24083 26724 24089
rect 23164 24024 24992 24052
rect 23164 24012 23170 24024
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 25961 24055 26019 24061
rect 25961 24052 25973 24055
rect 25648 24024 25973 24052
rect 25648 24012 25654 24024
rect 25961 24021 25973 24024
rect 26007 24021 26019 24055
rect 25961 24015 26019 24021
rect 27798 24012 27804 24064
rect 27856 24012 27862 24064
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 1857 23851 1915 23857
rect 1857 23817 1869 23851
rect 1903 23817 1915 23851
rect 1857 23811 1915 23817
rect 1949 23851 2007 23857
rect 1949 23817 1961 23851
rect 1995 23848 2007 23851
rect 1995 23820 2774 23848
rect 1995 23817 2007 23820
rect 1949 23811 2007 23817
rect 1762 23740 1768 23792
rect 1820 23740 1826 23792
rect 1872 23780 1900 23811
rect 1872 23752 2544 23780
rect 2130 23672 2136 23724
rect 2188 23672 2194 23724
rect 2516 23712 2544 23752
rect 2590 23740 2596 23792
rect 2648 23740 2654 23792
rect 2746 23780 2774 23820
rect 2958 23808 2964 23860
rect 3016 23848 3022 23860
rect 3878 23848 3884 23860
rect 3016 23820 3884 23848
rect 3016 23808 3022 23820
rect 3878 23808 3884 23820
rect 3936 23808 3942 23860
rect 4430 23808 4436 23860
rect 4488 23848 4494 23860
rect 4614 23848 4620 23860
rect 4488 23820 4620 23848
rect 4488 23808 4494 23820
rect 4614 23808 4620 23820
rect 4672 23848 4678 23860
rect 5077 23851 5135 23857
rect 5077 23848 5089 23851
rect 4672 23820 5089 23848
rect 4672 23808 4678 23820
rect 5077 23817 5089 23820
rect 5123 23817 5135 23851
rect 5077 23811 5135 23817
rect 5169 23851 5227 23857
rect 5169 23817 5181 23851
rect 5215 23848 5227 23851
rect 6270 23848 6276 23860
rect 5215 23820 6276 23848
rect 5215 23817 5227 23820
rect 5169 23811 5227 23817
rect 2746 23752 3556 23780
rect 3418 23712 3424 23724
rect 2516 23684 3424 23712
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 3528 23644 3556 23752
rect 3970 23740 3976 23792
rect 4028 23780 4034 23792
rect 4801 23783 4859 23789
rect 4801 23780 4813 23783
rect 4028 23752 4813 23780
rect 4028 23740 4034 23752
rect 4801 23749 4813 23752
rect 4847 23749 4859 23783
rect 5184 23780 5212 23811
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 6362 23808 6368 23860
rect 6420 23848 6426 23860
rect 6730 23848 6736 23860
rect 6420 23820 6736 23848
rect 6420 23808 6426 23820
rect 6730 23808 6736 23820
rect 6788 23808 6794 23860
rect 7282 23808 7288 23860
rect 7340 23848 7346 23860
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 7340 23820 7849 23848
rect 7340 23808 7346 23820
rect 7837 23817 7849 23820
rect 7883 23817 7895 23851
rect 7837 23811 7895 23817
rect 9585 23851 9643 23857
rect 9585 23817 9597 23851
rect 9631 23848 9643 23851
rect 9858 23848 9864 23860
rect 9631 23820 9864 23848
rect 9631 23817 9643 23820
rect 9585 23811 9643 23817
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 10594 23808 10600 23860
rect 10652 23848 10658 23860
rect 10981 23851 11039 23857
rect 10981 23848 10993 23851
rect 10652 23820 10993 23848
rect 10652 23808 10658 23820
rect 10981 23817 10993 23820
rect 11027 23817 11039 23851
rect 10981 23811 11039 23817
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 11701 23851 11759 23857
rect 11701 23848 11713 23851
rect 11296 23820 11713 23848
rect 11296 23808 11302 23820
rect 11701 23817 11713 23820
rect 11747 23817 11759 23851
rect 13357 23851 13415 23857
rect 11701 23811 11759 23817
rect 11900 23820 12434 23848
rect 5718 23780 5724 23792
rect 4801 23743 4859 23749
rect 4908 23752 5212 23780
rect 5276 23752 5724 23780
rect 3878 23672 3884 23724
rect 3936 23712 3942 23724
rect 4908 23712 4936 23752
rect 3936 23684 4936 23712
rect 4985 23715 5043 23721
rect 3936 23672 3942 23684
rect 4985 23681 4997 23715
rect 5031 23712 5043 23715
rect 5276 23712 5304 23752
rect 5718 23740 5724 23752
rect 5776 23740 5782 23792
rect 5828 23752 10732 23780
rect 5031 23684 5304 23712
rect 5353 23715 5411 23721
rect 5031 23681 5043 23684
rect 4985 23675 5043 23681
rect 5353 23681 5365 23715
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 4706 23644 4712 23656
rect 3528 23616 4712 23644
rect 4706 23604 4712 23616
rect 4764 23604 4770 23656
rect 474 23536 480 23588
rect 532 23576 538 23588
rect 1581 23579 1639 23585
rect 1581 23576 1593 23579
rect 532 23548 1593 23576
rect 532 23536 538 23548
rect 1581 23545 1593 23548
rect 1627 23545 1639 23579
rect 1581 23539 1639 23545
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 5368 23576 5396 23675
rect 5828 23585 5856 23752
rect 5997 23715 6055 23721
rect 5997 23681 6009 23715
rect 6043 23712 6055 23715
rect 6454 23712 6460 23724
rect 6043 23684 6460 23712
rect 6043 23681 6055 23684
rect 5997 23675 6055 23681
rect 6454 23672 6460 23684
rect 6512 23672 6518 23724
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23712 6975 23715
rect 7006 23712 7012 23724
rect 6963 23684 7012 23712
rect 6963 23681 6975 23684
rect 6917 23675 6975 23681
rect 6362 23604 6368 23656
rect 6420 23644 6426 23656
rect 6656 23644 6684 23675
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 7374 23672 7380 23724
rect 7432 23712 7438 23724
rect 7469 23715 7527 23721
rect 7469 23712 7481 23715
rect 7432 23684 7481 23712
rect 7432 23672 7438 23684
rect 7469 23681 7481 23684
rect 7515 23681 7527 23715
rect 8846 23712 8852 23724
rect 8904 23721 8910 23724
rect 8904 23715 8925 23721
rect 7469 23675 7527 23681
rect 7852 23684 8852 23712
rect 7852 23656 7880 23684
rect 8846 23672 8852 23684
rect 8913 23681 8925 23715
rect 8904 23675 8925 23681
rect 8904 23672 8910 23675
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9824 23684 9965 23712
rect 9824 23672 9830 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 10704 23712 10732 23752
rect 10778 23740 10784 23792
rect 10836 23740 10842 23792
rect 11900 23780 11928 23820
rect 10888 23752 11928 23780
rect 10888 23712 10916 23752
rect 11974 23740 11980 23792
rect 12032 23780 12038 23792
rect 12406 23780 12434 23820
rect 13357 23817 13369 23851
rect 13403 23848 13415 23851
rect 13446 23848 13452 23860
rect 13403 23820 13452 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 13814 23808 13820 23860
rect 13872 23808 13878 23860
rect 14734 23808 14740 23860
rect 14792 23848 14798 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 14792 23820 15025 23848
rect 14792 23808 14798 23820
rect 15013 23817 15025 23820
rect 15059 23817 15071 23851
rect 15841 23851 15899 23857
rect 15013 23811 15071 23817
rect 15120 23820 15793 23848
rect 13538 23780 13544 23792
rect 12032 23752 12204 23780
rect 12406 23752 13544 23780
rect 12032 23740 12038 23752
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 10704 23684 10916 23712
rect 10980 23684 12081 23712
rect 9953 23675 10011 23681
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 6420 23616 7573 23644
rect 6420 23604 6426 23616
rect 7561 23613 7573 23616
rect 7607 23644 7619 23647
rect 7834 23644 7840 23656
rect 7607 23616 7840 23644
rect 7607 23613 7619 23616
rect 7561 23607 7619 23613
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8386 23604 8392 23656
rect 8444 23604 8450 23656
rect 8570 23604 8576 23656
rect 8628 23604 8634 23656
rect 8966 23647 9024 23653
rect 8966 23644 8978 23647
rect 8680 23616 8978 23644
rect 4120 23548 5396 23576
rect 5813 23579 5871 23585
rect 4120 23536 4126 23548
rect 5813 23545 5825 23579
rect 5859 23545 5871 23579
rect 5813 23539 5871 23545
rect 6914 23536 6920 23588
rect 6972 23536 6978 23588
rect 4154 23468 4160 23520
rect 4212 23508 4218 23520
rect 4890 23508 4896 23520
rect 4212 23480 4896 23508
rect 4212 23468 4218 23480
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 7653 23511 7711 23517
rect 7653 23477 7665 23511
rect 7699 23508 7711 23511
rect 7926 23508 7932 23520
rect 7699 23480 7932 23508
rect 7699 23477 7711 23480
rect 7653 23471 7711 23477
rect 7926 23468 7932 23480
rect 7984 23508 7990 23520
rect 8680 23508 8708 23616
rect 8966 23613 8978 23616
rect 9012 23644 9024 23647
rect 9306 23644 9312 23656
rect 9012 23616 9312 23644
rect 9012 23613 9024 23616
rect 8966 23607 9024 23613
rect 9306 23604 9312 23616
rect 9364 23644 9370 23656
rect 9858 23644 9864 23656
rect 9364 23616 9864 23644
rect 9364 23604 9370 23616
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 10042 23604 10048 23656
rect 10100 23604 10106 23656
rect 10226 23604 10232 23656
rect 10284 23604 10290 23656
rect 10980 23644 11008 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12176 23712 12204 23752
rect 13538 23740 13544 23752
rect 13596 23740 13602 23792
rect 14645 23783 14703 23789
rect 14645 23749 14657 23783
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 14861 23783 14919 23789
rect 14861 23749 14873 23783
rect 14907 23780 14919 23783
rect 15120 23780 15148 23820
rect 14907 23752 15148 23780
rect 14907 23749 14919 23752
rect 14861 23743 14919 23749
rect 12894 23712 12900 23724
rect 12176 23684 12900 23712
rect 12069 23675 12127 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 12986 23672 12992 23724
rect 13044 23672 13050 23724
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 10428 23616 11008 23644
rect 9766 23536 9772 23588
rect 9824 23576 9830 23588
rect 10244 23576 10272 23604
rect 9824 23548 10272 23576
rect 9824 23536 9830 23548
rect 7984 23480 8708 23508
rect 7984 23468 7990 23480
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 10428 23508 10456 23616
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11882 23644 11888 23656
rect 11112 23616 11888 23644
rect 11112 23604 11118 23616
rect 11882 23604 11888 23616
rect 11940 23644 11946 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 11940 23616 12173 23644
rect 11940 23604 11946 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 12345 23647 12403 23653
rect 12345 23613 12357 23647
rect 12391 23644 12403 23647
rect 12434 23644 12440 23656
rect 12391 23616 12440 23644
rect 12391 23613 12403 23616
rect 12345 23607 12403 23613
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 13188 23644 13216 23675
rect 13262 23672 13268 23724
rect 13320 23712 13326 23724
rect 14001 23715 14059 23721
rect 14001 23712 14013 23715
rect 13320 23684 14013 23712
rect 13320 23672 13326 23684
rect 14001 23681 14013 23684
rect 14047 23681 14059 23715
rect 14660 23712 14688 23743
rect 15194 23740 15200 23792
rect 15252 23780 15258 23792
rect 15473 23783 15531 23789
rect 15473 23780 15485 23783
rect 15252 23752 15485 23780
rect 15252 23740 15258 23752
rect 15473 23749 15485 23752
rect 15519 23749 15531 23783
rect 15473 23743 15531 23749
rect 15678 23783 15736 23789
rect 15678 23749 15690 23783
rect 15724 23749 15736 23783
rect 15765 23780 15793 23820
rect 15841 23817 15853 23851
rect 15887 23848 15899 23851
rect 17954 23848 17960 23860
rect 15887 23820 17960 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 18690 23848 18696 23860
rect 18196 23820 18696 23848
rect 18196 23808 18202 23820
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 19978 23848 19984 23860
rect 18892 23820 19984 23848
rect 16298 23780 16304 23792
rect 15765 23752 16304 23780
rect 15678 23743 15736 23749
rect 15010 23712 15016 23724
rect 14660 23684 15016 23712
rect 14001 23675 14059 23681
rect 15010 23672 15016 23684
rect 15068 23672 15074 23724
rect 14458 23644 14464 23656
rect 13188 23616 14464 23644
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 14734 23604 14740 23656
rect 14792 23644 14798 23656
rect 15688 23644 15716 23743
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 16850 23740 16856 23792
rect 16908 23780 16914 23792
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 16908 23752 16957 23780
rect 16908 23740 16914 23752
rect 16945 23749 16957 23752
rect 16991 23749 17003 23783
rect 16945 23743 17003 23749
rect 17310 23740 17316 23792
rect 17368 23780 17374 23792
rect 18046 23780 18052 23792
rect 17368 23752 18052 23780
rect 17368 23740 17374 23752
rect 18046 23740 18052 23752
rect 18104 23740 18110 23792
rect 15930 23672 15936 23724
rect 15988 23712 15994 23724
rect 15988 23684 17448 23712
rect 15988 23672 15994 23684
rect 17310 23644 17316 23656
rect 14792 23616 17316 23644
rect 14792 23604 14798 23616
rect 17310 23604 17316 23616
rect 17368 23604 17374 23656
rect 17420 23644 17448 23684
rect 17770 23672 17776 23724
rect 17828 23672 17834 23724
rect 18782 23672 18788 23724
rect 18840 23672 18846 23724
rect 18892 23644 18920 23820
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 20162 23808 20168 23860
rect 20220 23848 20226 23860
rect 20441 23851 20499 23857
rect 20441 23848 20453 23851
rect 20220 23820 20453 23848
rect 20220 23808 20226 23820
rect 20441 23817 20453 23820
rect 20487 23817 20499 23851
rect 20441 23811 20499 23817
rect 21085 23851 21143 23857
rect 21085 23817 21097 23851
rect 21131 23848 21143 23851
rect 22278 23848 22284 23860
rect 21131 23820 22284 23848
rect 21131 23817 21143 23820
rect 21085 23811 21143 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22370 23808 22376 23860
rect 22428 23848 22434 23860
rect 24581 23851 24639 23857
rect 24581 23848 24593 23851
rect 22428 23820 24593 23848
rect 22428 23808 22434 23820
rect 24581 23817 24593 23820
rect 24627 23817 24639 23851
rect 24581 23811 24639 23817
rect 24762 23808 24768 23860
rect 24820 23848 24826 23860
rect 28350 23848 28356 23860
rect 24820 23820 28356 23848
rect 24820 23808 24826 23820
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 19153 23783 19211 23789
rect 19153 23749 19165 23783
rect 19199 23780 19211 23783
rect 23566 23780 23572 23792
rect 19199 23752 21312 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 18966 23672 18972 23724
rect 19024 23672 19030 23724
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 20254 23712 20260 23724
rect 19843 23684 20260 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 20622 23672 20628 23724
rect 20680 23672 20686 23724
rect 21284 23721 21312 23752
rect 23124 23752 23572 23780
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23681 21327 23715
rect 21269 23675 21327 23681
rect 22278 23672 22284 23724
rect 22336 23672 22342 23724
rect 17420 23616 18920 23644
rect 19981 23647 20039 23653
rect 19981 23613 19993 23647
rect 20027 23644 20039 23647
rect 23014 23644 23020 23656
rect 20027 23616 23020 23644
rect 20027 23613 20039 23616
rect 19981 23607 20039 23613
rect 23014 23604 23020 23616
rect 23072 23604 23078 23656
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 12526 23576 12532 23588
rect 11195 23548 12532 23576
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 12894 23536 12900 23588
rect 12952 23576 12958 23588
rect 17589 23579 17647 23585
rect 12952 23548 17152 23576
rect 12952 23536 12958 23548
rect 9640 23480 10456 23508
rect 9640 23468 9646 23480
rect 10502 23468 10508 23520
rect 10560 23508 10566 23520
rect 10965 23511 11023 23517
rect 10965 23508 10977 23511
rect 10560 23480 10977 23508
rect 10560 23468 10566 23480
rect 10965 23477 10977 23480
rect 11011 23477 11023 23511
rect 10965 23471 11023 23477
rect 14826 23468 14832 23520
rect 14884 23468 14890 23520
rect 15654 23468 15660 23520
rect 15712 23468 15718 23520
rect 16206 23468 16212 23520
rect 16264 23508 16270 23520
rect 17037 23511 17095 23517
rect 17037 23508 17049 23511
rect 16264 23480 17049 23508
rect 16264 23468 16270 23480
rect 17037 23477 17049 23480
rect 17083 23477 17095 23511
rect 17124 23508 17152 23548
rect 17589 23545 17601 23579
rect 17635 23576 17647 23579
rect 20438 23576 20444 23588
rect 17635 23548 20444 23576
rect 17635 23545 17647 23548
rect 17589 23539 17647 23545
rect 20438 23536 20444 23548
rect 20496 23536 20502 23588
rect 21266 23536 21272 23588
rect 21324 23576 21330 23588
rect 23124 23576 23152 23752
rect 23566 23740 23572 23752
rect 23624 23740 23630 23792
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23712 23259 23715
rect 23290 23712 23296 23724
rect 23247 23684 23296 23712
rect 23247 23681 23259 23684
rect 23201 23675 23259 23681
rect 23290 23672 23296 23684
rect 23348 23672 23354 23724
rect 23474 23721 23480 23724
rect 23468 23675 23480 23721
rect 23474 23672 23480 23675
rect 23532 23672 23538 23724
rect 24210 23672 24216 23724
rect 24268 23712 24274 23724
rect 25481 23715 25539 23721
rect 25481 23712 25493 23715
rect 24268 23684 25493 23712
rect 24268 23672 24274 23684
rect 25481 23681 25493 23684
rect 25527 23681 25539 23715
rect 25481 23675 25539 23681
rect 25225 23647 25283 23653
rect 25225 23613 25237 23647
rect 25271 23613 25283 23647
rect 25225 23607 25283 23613
rect 21324 23548 23152 23576
rect 21324 23536 21330 23548
rect 20714 23508 20720 23520
rect 17124 23480 20720 23508
rect 17037 23471 17095 23477
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 22097 23511 22155 23517
rect 22097 23477 22109 23511
rect 22143 23508 22155 23511
rect 23934 23508 23940 23520
rect 22143 23480 23940 23508
rect 22143 23477 22155 23480
rect 22097 23471 22155 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24486 23508 24492 23520
rect 24176 23480 24492 23508
rect 24176 23468 24182 23480
rect 24486 23468 24492 23480
rect 24544 23508 24550 23520
rect 25240 23508 25268 23607
rect 26142 23508 26148 23520
rect 24544 23480 26148 23508
rect 24544 23468 24550 23480
rect 26142 23468 26148 23480
rect 26200 23468 26206 23520
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 2501 23307 2559 23313
rect 2501 23304 2513 23307
rect 1912 23276 2513 23304
rect 1912 23264 1918 23276
rect 2501 23273 2513 23276
rect 2547 23273 2559 23307
rect 2501 23267 2559 23273
rect 4062 23264 4068 23316
rect 4120 23264 4126 23316
rect 5810 23304 5816 23316
rect 4356 23276 5816 23304
rect 1673 23239 1731 23245
rect 1673 23205 1685 23239
rect 1719 23236 1731 23239
rect 2406 23236 2412 23248
rect 1719 23208 2412 23236
rect 1719 23205 1731 23208
rect 1673 23199 1731 23205
rect 2406 23196 2412 23208
rect 2464 23196 2470 23248
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 3053 23171 3111 23177
rect 3053 23168 3065 23171
rect 3016 23140 3065 23168
rect 3016 23128 3022 23140
rect 3053 23137 3065 23140
rect 3099 23137 3111 23171
rect 3053 23131 3111 23137
rect 3694 23128 3700 23180
rect 3752 23168 3758 23180
rect 4356 23168 4384 23276
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 6380 23276 7328 23304
rect 6380 23236 6408 23276
rect 3752 23140 4384 23168
rect 3752 23128 3758 23140
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 1854 23100 1860 23112
rect 1719 23072 1860 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 4356 23109 4384 23140
rect 5276 23208 6408 23236
rect 6457 23239 6515 23245
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23069 2007 23103
rect 1949 23063 2007 23069
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 4341 23103 4399 23109
rect 2823 23072 4108 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 1302 22992 1308 23044
rect 1360 23032 1366 23044
rect 1964 23032 1992 23063
rect 1360 23004 1992 23032
rect 1360 22992 1366 23004
rect 2958 22992 2964 23044
rect 3016 22992 3022 23044
rect 4080 23032 4108 23072
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 4430 23060 4436 23112
rect 4488 23060 4494 23112
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23100 4583 23103
rect 4614 23100 4620 23112
rect 4571 23072 4620 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 4709 23103 4767 23109
rect 4709 23069 4721 23103
rect 4755 23100 4767 23103
rect 4982 23100 4988 23112
rect 4755 23072 4988 23100
rect 4755 23069 4767 23072
rect 4709 23063 4767 23069
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 5276 23032 5304 23208
rect 6457 23205 6469 23239
rect 6503 23236 6515 23239
rect 6546 23236 6552 23248
rect 6503 23208 6552 23236
rect 6503 23205 6515 23208
rect 6457 23199 6515 23205
rect 6546 23196 6552 23208
rect 6604 23196 6610 23248
rect 7300 23236 7328 23276
rect 7374 23264 7380 23316
rect 7432 23304 7438 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 7432 23276 7849 23304
rect 7432 23264 7438 23276
rect 7837 23273 7849 23276
rect 7883 23304 7895 23307
rect 8386 23304 8392 23316
rect 7883 23276 8392 23304
rect 7883 23273 7895 23276
rect 7837 23267 7895 23273
rect 8386 23264 8392 23276
rect 8444 23264 8450 23316
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10870 23304 10876 23316
rect 9732 23276 10876 23304
rect 9732 23264 9738 23276
rect 10870 23264 10876 23276
rect 10928 23264 10934 23316
rect 11333 23307 11391 23313
rect 11333 23273 11345 23307
rect 11379 23304 11391 23307
rect 11790 23304 11796 23316
rect 11379 23276 11796 23304
rect 11379 23273 11391 23276
rect 11333 23267 11391 23273
rect 11790 23264 11796 23276
rect 11848 23264 11854 23316
rect 12158 23264 12164 23316
rect 12216 23304 12222 23316
rect 12802 23304 12808 23316
rect 12216 23276 12808 23304
rect 12216 23264 12222 23276
rect 12802 23264 12808 23276
rect 12860 23264 12866 23316
rect 13541 23307 13599 23313
rect 13541 23273 13553 23307
rect 13587 23273 13599 23307
rect 13541 23267 13599 23273
rect 13725 23307 13783 23313
rect 13725 23273 13737 23307
rect 13771 23304 13783 23307
rect 14550 23304 14556 23316
rect 13771 23276 14556 23304
rect 13771 23273 13783 23276
rect 13725 23267 13783 23273
rect 10778 23236 10784 23248
rect 7300 23208 10784 23236
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 11238 23196 11244 23248
rect 11296 23236 11302 23248
rect 12894 23236 12900 23248
rect 11296 23208 12900 23236
rect 11296 23196 11302 23208
rect 12894 23196 12900 23208
rect 12952 23196 12958 23248
rect 13556 23236 13584 23267
rect 14550 23264 14556 23276
rect 14608 23264 14614 23316
rect 15010 23264 15016 23316
rect 15068 23304 15074 23316
rect 15746 23304 15752 23316
rect 15068 23276 15752 23304
rect 15068 23264 15074 23276
rect 15746 23264 15752 23276
rect 15804 23264 15810 23316
rect 16022 23264 16028 23316
rect 16080 23264 16086 23316
rect 16390 23264 16396 23316
rect 16448 23304 16454 23316
rect 17037 23307 17095 23313
rect 17037 23304 17049 23307
rect 16448 23276 17049 23304
rect 16448 23264 16454 23276
rect 17037 23273 17049 23276
rect 17083 23273 17095 23307
rect 17037 23267 17095 23273
rect 17586 23264 17592 23316
rect 17644 23304 17650 23316
rect 17865 23307 17923 23313
rect 17865 23304 17877 23307
rect 17644 23276 17877 23304
rect 17644 23264 17650 23276
rect 17865 23273 17877 23276
rect 17911 23273 17923 23307
rect 17865 23267 17923 23273
rect 18874 23264 18880 23316
rect 18932 23264 18938 23316
rect 19889 23307 19947 23313
rect 19889 23273 19901 23307
rect 19935 23304 19947 23307
rect 20070 23304 20076 23316
rect 19935 23276 20076 23304
rect 19935 23273 19947 23276
rect 19889 23267 19947 23273
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 20548 23276 21925 23304
rect 14366 23236 14372 23248
rect 13556 23208 14372 23236
rect 14366 23196 14372 23208
rect 14424 23196 14430 23248
rect 14642 23196 14648 23248
rect 14700 23196 14706 23248
rect 15197 23239 15255 23245
rect 15197 23205 15209 23239
rect 15243 23205 15255 23239
rect 15197 23199 15255 23205
rect 6638 23168 6644 23180
rect 5368 23140 6644 23168
rect 5368 23109 5396 23140
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 7926 23168 7932 23180
rect 7484 23140 7932 23168
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5534 23060 5540 23112
rect 5592 23060 5598 23112
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5718 23100 5724 23112
rect 5675 23072 5724 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5994 23060 6000 23112
rect 6052 23100 6058 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 6052 23072 6285 23100
rect 6052 23060 6058 23072
rect 6273 23069 6285 23072
rect 6319 23069 6331 23103
rect 6273 23063 6331 23069
rect 6549 23103 6607 23109
rect 6549 23069 6561 23103
rect 6595 23100 6607 23103
rect 6822 23100 6828 23112
rect 6595 23072 6828 23100
rect 6595 23069 6607 23072
rect 6549 23063 6607 23069
rect 4080 23004 5304 23032
rect 5810 22992 5816 23044
rect 5868 23032 5874 23044
rect 6564 23032 6592 23063
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 7484 23109 7512 23140
rect 7926 23128 7932 23140
rect 7984 23128 7990 23180
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9364 23140 9689 23168
rect 9364 23128 9370 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 11054 23168 11060 23180
rect 9677 23131 9735 23137
rect 10260 23140 11060 23168
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23069 7527 23103
rect 7469 23063 7527 23069
rect 7834 23060 7840 23112
rect 7892 23060 7898 23112
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 10260 23100 10288 23140
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 12342 23168 12348 23180
rect 11532 23140 12348 23168
rect 9539 23072 10288 23100
rect 10321 23103 10379 23109
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 10321 23069 10333 23103
rect 10367 23069 10379 23103
rect 10321 23063 10379 23069
rect 5868 23004 6592 23032
rect 5868 22992 5874 23004
rect 7190 22992 7196 23044
rect 7248 23032 7254 23044
rect 10336 23032 10364 23063
rect 10410 23060 10416 23112
rect 10468 23100 10474 23112
rect 10505 23103 10563 23109
rect 10505 23100 10517 23103
rect 10468 23072 10517 23100
rect 10468 23060 10474 23072
rect 10505 23069 10517 23072
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 11532 23109 11560 23140
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 13998 23128 14004 23180
rect 14056 23168 14062 23180
rect 14550 23168 14556 23180
rect 14056 23140 14556 23168
rect 14056 23128 14062 23140
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 14737 23171 14795 23177
rect 14737 23137 14749 23171
rect 14783 23137 14795 23171
rect 15212 23168 15240 23199
rect 15378 23196 15384 23248
rect 15436 23236 15442 23248
rect 16209 23239 16267 23245
rect 16209 23236 16221 23239
rect 15436 23208 16221 23236
rect 15436 23196 15442 23208
rect 16209 23205 16221 23208
rect 16255 23205 16267 23239
rect 16209 23199 16267 23205
rect 18506 23196 18512 23248
rect 18564 23236 18570 23248
rect 19150 23236 19156 23248
rect 18564 23208 19156 23236
rect 18564 23196 18570 23208
rect 19150 23196 19156 23208
rect 19208 23196 19214 23248
rect 19702 23196 19708 23248
rect 19760 23196 19766 23248
rect 19978 23196 19984 23248
rect 20036 23236 20042 23248
rect 20548 23236 20576 23276
rect 21913 23273 21925 23276
rect 21959 23273 21971 23307
rect 21913 23267 21971 23273
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22888 23276 22937 23304
rect 22888 23264 22894 23276
rect 22925 23273 22937 23276
rect 22971 23304 22983 23307
rect 23290 23304 23296 23316
rect 22971 23276 23296 23304
rect 22971 23273 22983 23276
rect 22925 23267 22983 23273
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23304 23535 23307
rect 24854 23304 24860 23316
rect 23523 23276 24860 23304
rect 23523 23273 23535 23276
rect 23477 23267 23535 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 27433 23307 27491 23313
rect 27433 23304 27445 23307
rect 24964 23276 27445 23304
rect 20036 23208 20576 23236
rect 20036 23196 20042 23208
rect 22462 23196 22468 23248
rect 22520 23236 22526 23248
rect 24964 23236 24992 23276
rect 27433 23273 27445 23276
rect 27479 23273 27491 23307
rect 27433 23267 27491 23273
rect 22520 23208 24992 23236
rect 22520 23196 22526 23208
rect 16758 23168 16764 23180
rect 15212 23140 16764 23168
rect 14737 23131 14795 23137
rect 12158 23109 12164 23112
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 11977 23063 12035 23069
rect 12125 23103 12164 23109
rect 12125 23069 12137 23103
rect 12125 23063 12164 23069
rect 10597 23035 10655 23041
rect 10597 23032 10609 23035
rect 7248 23004 10364 23032
rect 7248 22992 7254 23004
rect 10336 22976 10364 23004
rect 10520 23004 10609 23032
rect 10520 22976 10548 23004
rect 10597 23001 10609 23004
rect 10643 23001 10655 23035
rect 11992 23032 12020 23063
rect 12158 23060 12164 23063
rect 12216 23060 12222 23112
rect 12434 23060 12440 23112
rect 12492 23109 12498 23112
rect 12492 23100 12500 23109
rect 12618 23100 12624 23112
rect 12492 23072 12624 23100
rect 12492 23063 12500 23072
rect 12492 23060 12498 23063
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 14752 23100 14780 23131
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 18748 23140 20668 23168
rect 18748 23128 18754 23140
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 13372 23072 14412 23100
rect 14752 23072 15393 23100
rect 10597 22995 10655 23001
rect 10888 23004 12020 23032
rect 12253 23035 12311 23041
rect 1857 22967 1915 22973
rect 1857 22933 1869 22967
rect 1903 22964 1915 22967
rect 2498 22964 2504 22976
rect 1903 22936 2504 22964
rect 1903 22933 1915 22936
rect 1857 22927 1915 22933
rect 2498 22924 2504 22936
rect 2556 22924 2562 22976
rect 3050 22924 3056 22976
rect 3108 22964 3114 22976
rect 4062 22964 4068 22976
rect 3108 22936 4068 22964
rect 3108 22924 3114 22936
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4246 22924 4252 22976
rect 4304 22964 4310 22976
rect 5169 22967 5227 22973
rect 5169 22964 5181 22967
rect 4304 22936 5181 22964
rect 4304 22924 4310 22936
rect 5169 22933 5181 22936
rect 5215 22933 5227 22967
rect 5169 22927 5227 22933
rect 6086 22924 6092 22976
rect 6144 22924 6150 22976
rect 6178 22924 6184 22976
rect 6236 22964 6242 22976
rect 8021 22967 8079 22973
rect 8021 22964 8033 22967
rect 6236 22936 8033 22964
rect 6236 22924 6242 22936
rect 8021 22933 8033 22936
rect 8067 22933 8079 22967
rect 8021 22927 8079 22933
rect 9122 22924 9128 22976
rect 9180 22924 9186 22976
rect 9582 22924 9588 22976
rect 9640 22924 9646 22976
rect 10318 22924 10324 22976
rect 10376 22924 10382 22976
rect 10502 22924 10508 22976
rect 10560 22924 10566 22976
rect 10888 22973 10916 23004
rect 12253 23001 12265 23035
rect 12299 23001 12311 23035
rect 12253 22995 12311 23001
rect 10873 22967 10931 22973
rect 10873 22933 10885 22967
rect 10919 22933 10931 22967
rect 10873 22927 10931 22933
rect 11882 22924 11888 22976
rect 11940 22964 11946 22976
rect 12066 22964 12072 22976
rect 11940 22936 12072 22964
rect 11940 22924 11946 22936
rect 12066 22924 12072 22936
rect 12124 22964 12130 22976
rect 12268 22964 12296 22995
rect 12342 22992 12348 23044
rect 12400 22992 12406 23044
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 13372 23041 13400 23072
rect 13357 23035 13415 23041
rect 13357 23032 13369 23035
rect 13228 23004 13369 23032
rect 13228 22992 13234 23004
rect 13357 23001 13369 23004
rect 13403 23001 13415 23035
rect 13357 22995 13415 23001
rect 14274 22992 14280 23044
rect 14332 22992 14338 23044
rect 14384 23032 14412 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 16206 23100 16212 23112
rect 15381 23063 15439 23069
rect 15488 23072 16212 23100
rect 15488 23032 15516 23072
rect 16206 23060 16212 23072
rect 16264 23100 16270 23112
rect 16669 23103 16727 23109
rect 16669 23100 16681 23103
rect 16264 23072 16681 23100
rect 16264 23060 16270 23072
rect 16669 23069 16681 23072
rect 16715 23069 16727 23103
rect 16853 23103 16911 23109
rect 16853 23100 16865 23103
rect 16669 23063 16727 23069
rect 16756 23072 16865 23100
rect 14384 23004 15516 23032
rect 15746 22992 15752 23044
rect 15804 23032 15810 23044
rect 15841 23035 15899 23041
rect 15841 23032 15853 23035
rect 15804 23004 15853 23032
rect 15804 22992 15810 23004
rect 15841 23001 15853 23004
rect 15887 23001 15899 23035
rect 15841 22995 15899 23001
rect 16574 22992 16580 23044
rect 16632 23032 16638 23044
rect 16756 23032 16784 23072
rect 16853 23069 16865 23072
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 17126 23060 17132 23112
rect 17184 23100 17190 23112
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 17184 23072 17509 23100
rect 17184 23060 17190 23072
rect 17497 23069 17509 23072
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 19334 23100 19340 23112
rect 17920 23072 19340 23100
rect 17920 23060 17926 23072
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20533 23103 20591 23109
rect 20533 23100 20545 23103
rect 20220 23072 20545 23100
rect 20220 23060 20226 23072
rect 20533 23069 20545 23072
rect 20579 23069 20591 23103
rect 20640 23100 20668 23140
rect 22370 23128 22376 23180
rect 22428 23168 22434 23180
rect 22428 23140 25912 23168
rect 22428 23128 22434 23140
rect 22833 23103 22891 23109
rect 20640 23072 22784 23100
rect 20533 23063 20591 23069
rect 18509 23035 18567 23041
rect 18509 23032 18521 23035
rect 16632 23004 16784 23032
rect 16868 23004 18521 23032
rect 16632 22992 16638 23004
rect 16868 22976 16896 23004
rect 18509 23001 18521 23004
rect 18555 23001 18567 23035
rect 18509 22995 18567 23001
rect 12124 22936 12296 22964
rect 12621 22967 12679 22973
rect 12124 22924 12130 22936
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 13446 22964 13452 22976
rect 12667 22936 13452 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 13446 22924 13452 22936
rect 13504 22924 13510 22976
rect 13538 22924 13544 22976
rect 13596 22973 13602 22976
rect 13596 22967 13615 22973
rect 13603 22933 13615 22967
rect 13596 22927 13615 22933
rect 13596 22924 13602 22927
rect 15286 22924 15292 22976
rect 15344 22964 15350 22976
rect 16041 22967 16099 22973
rect 16041 22964 16053 22967
rect 15344 22936 16053 22964
rect 15344 22924 15350 22936
rect 16041 22933 16053 22936
rect 16087 22933 16099 22967
rect 16041 22927 16099 22933
rect 16850 22924 16856 22976
rect 16908 22924 16914 22976
rect 18524 22964 18552 22995
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 18693 23035 18751 23041
rect 18693 23032 18705 23035
rect 18656 23004 18705 23032
rect 18656 22992 18662 23004
rect 18693 23001 18705 23004
rect 18739 23001 18751 23035
rect 18693 22995 18751 23001
rect 19426 22992 19432 23044
rect 19484 22992 19490 23044
rect 20070 22992 20076 23044
rect 20128 23032 20134 23044
rect 20778 23035 20836 23041
rect 20778 23032 20790 23035
rect 20128 23004 20790 23032
rect 20128 22992 20134 23004
rect 20778 23001 20790 23004
rect 20824 23001 20836 23035
rect 20778 22995 20836 23001
rect 18782 22964 18788 22976
rect 18524 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22964 18846 22976
rect 19150 22964 19156 22976
rect 18840 22936 19156 22964
rect 18840 22924 18846 22936
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19886 22964 19892 22976
rect 19392 22936 19892 22964
rect 19392 22924 19398 22936
rect 19886 22924 19892 22936
rect 19944 22924 19950 22976
rect 22756 22964 22784 23072
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23014 23100 23020 23112
rect 22879 23072 23020 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 23014 23060 23020 23072
rect 23072 23060 23078 23112
rect 23661 23103 23719 23109
rect 23661 23100 23673 23103
rect 23584 23072 23673 23100
rect 23290 22992 23296 23044
rect 23348 23032 23354 23044
rect 23584 23032 23612 23072
rect 23661 23069 23673 23072
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23069 24823 23103
rect 24765 23063 24823 23069
rect 23348 23004 23612 23032
rect 23348 22992 23354 23004
rect 24394 22992 24400 23044
rect 24452 23032 24458 23044
rect 24780 23032 24808 23063
rect 24452 23004 24808 23032
rect 24452 22992 24458 23004
rect 24026 22964 24032 22976
rect 22756 22936 24032 22964
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 25774 22964 25780 22976
rect 24627 22936 25780 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 25774 22924 25780 22936
rect 25832 22924 25838 22976
rect 25884 22964 25912 23140
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23100 26111 23103
rect 26142 23100 26148 23112
rect 26099 23072 26148 23100
rect 26099 23069 26111 23072
rect 26053 23063 26111 23069
rect 26142 23060 26148 23072
rect 26200 23060 26206 23112
rect 26320 23035 26378 23041
rect 26320 23001 26332 23035
rect 26366 23032 26378 23035
rect 26510 23032 26516 23044
rect 26366 23004 26516 23032
rect 26366 23001 26378 23004
rect 26320 22995 26378 23001
rect 26510 22992 26516 23004
rect 26568 22992 26574 23044
rect 26418 22964 26424 22976
rect 25884 22936 26424 22964
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 1958 22763 2016 22769
rect 1958 22760 1970 22763
rect 1820 22732 1970 22760
rect 1820 22720 1826 22732
rect 1958 22729 1970 22732
rect 2004 22760 2016 22763
rect 2682 22760 2688 22772
rect 2004 22732 2688 22760
rect 2004 22729 2016 22732
rect 1958 22723 2016 22729
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 3694 22760 3700 22772
rect 3620 22732 3700 22760
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22593 1639 22627
rect 1581 22587 1639 22593
rect 1596 22556 1624 22587
rect 2130 22584 2136 22636
rect 2188 22624 2194 22636
rect 2225 22627 2283 22633
rect 2225 22624 2237 22627
rect 2188 22596 2237 22624
rect 2188 22584 2194 22596
rect 2225 22593 2237 22596
rect 2271 22593 2283 22627
rect 2225 22587 2283 22593
rect 3234 22584 3240 22636
rect 3292 22624 3298 22636
rect 3620 22633 3648 22732
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 4525 22763 4583 22769
rect 4525 22760 4537 22763
rect 3896 22732 4537 22760
rect 3513 22627 3571 22633
rect 3513 22624 3525 22627
rect 3292 22596 3525 22624
rect 3292 22584 3298 22596
rect 3513 22593 3525 22596
rect 3559 22593 3571 22627
rect 3513 22587 3571 22593
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22593 3663 22627
rect 3605 22587 3663 22593
rect 3694 22584 3700 22636
rect 3752 22584 3758 22636
rect 3896 22633 3924 22732
rect 4525 22729 4537 22732
rect 4571 22760 4583 22763
rect 4982 22760 4988 22772
rect 4571 22732 4988 22760
rect 4571 22729 4583 22732
rect 4525 22723 4583 22729
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 5077 22763 5135 22769
rect 5077 22729 5089 22763
rect 5123 22760 5135 22763
rect 5534 22760 5540 22772
rect 5123 22732 5540 22760
rect 5123 22729 5135 22732
rect 5077 22723 5135 22729
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 7285 22763 7343 22769
rect 7285 22729 7297 22763
rect 7331 22760 7343 22763
rect 7742 22760 7748 22772
rect 7331 22732 7748 22760
rect 7331 22729 7343 22732
rect 7285 22723 7343 22729
rect 7742 22720 7748 22732
rect 7800 22720 7806 22772
rect 9125 22763 9183 22769
rect 9125 22729 9137 22763
rect 9171 22729 9183 22763
rect 9125 22723 9183 22729
rect 6178 22692 6184 22704
rect 4356 22664 6184 22692
rect 4356 22633 4384 22664
rect 6178 22652 6184 22664
rect 6236 22652 6242 22704
rect 6454 22652 6460 22704
rect 6512 22692 6518 22704
rect 9140 22692 9168 22723
rect 10318 22720 10324 22772
rect 10376 22760 10382 22772
rect 10965 22763 11023 22769
rect 10965 22760 10977 22763
rect 10376 22732 10977 22760
rect 10376 22720 10382 22732
rect 10965 22729 10977 22732
rect 11011 22729 11023 22763
rect 10965 22723 11023 22729
rect 11790 22720 11796 22772
rect 11848 22760 11854 22772
rect 12342 22760 12348 22772
rect 11848 22732 12348 22760
rect 11848 22720 11854 22732
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 12897 22763 12955 22769
rect 12897 22729 12909 22763
rect 12943 22760 12955 22763
rect 13722 22760 13728 22772
rect 12943 22732 13728 22760
rect 12943 22729 12955 22732
rect 12897 22723 12955 22729
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 14090 22720 14096 22772
rect 14148 22760 14154 22772
rect 15378 22760 15384 22772
rect 14148 22732 15384 22760
rect 14148 22720 14154 22732
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 17770 22760 17776 22772
rect 17267 22732 17776 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 17954 22720 17960 22772
rect 18012 22720 18018 22772
rect 19334 22760 19340 22772
rect 19076 22732 19340 22760
rect 10134 22692 10140 22704
rect 6512 22664 9168 22692
rect 9232 22664 10140 22692
rect 6512 22652 6518 22664
rect 3881 22627 3939 22633
rect 3881 22593 3893 22627
rect 3927 22593 3939 22627
rect 3881 22587 3939 22593
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22593 4399 22627
rect 5445 22627 5503 22633
rect 5445 22624 5457 22627
rect 4341 22587 4399 22593
rect 4448 22596 5457 22624
rect 2038 22556 2044 22568
rect 1596 22528 2044 22556
rect 2038 22516 2044 22528
rect 2096 22556 2102 22568
rect 3970 22556 3976 22568
rect 2096 22528 3976 22556
rect 2096 22516 2102 22528
rect 3970 22516 3976 22528
rect 4028 22516 4034 22568
rect 4062 22516 4068 22568
rect 4120 22556 4126 22568
rect 4448 22556 4476 22596
rect 5445 22593 5457 22596
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22624 6883 22627
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 6871 22596 8677 22624
rect 6871 22593 6883 22596
rect 6825 22587 6883 22593
rect 8665 22593 8677 22596
rect 8711 22624 8723 22627
rect 9030 22624 9036 22636
rect 8711 22596 9036 22624
rect 8711 22593 8723 22596
rect 8665 22587 8723 22593
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 4120 22528 4476 22556
rect 4120 22516 4126 22528
rect 4982 22516 4988 22568
rect 5040 22556 5046 22568
rect 5537 22559 5595 22565
rect 5537 22556 5549 22559
rect 5040 22528 5549 22556
rect 5040 22516 5046 22528
rect 5537 22525 5549 22528
rect 5583 22525 5595 22559
rect 5537 22519 5595 22525
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22556 5687 22559
rect 5994 22556 6000 22568
rect 5675 22528 6000 22556
rect 5675 22525 5687 22528
rect 5629 22519 5687 22525
rect 4338 22488 4344 22500
rect 1964 22460 4344 22488
rect 1964 22429 1992 22460
rect 4338 22448 4344 22460
rect 4396 22448 4402 22500
rect 4448 22460 5396 22488
rect 1949 22423 2007 22429
rect 1949 22389 1961 22423
rect 1995 22389 2007 22423
rect 1949 22383 2007 22389
rect 2406 22380 2412 22432
rect 2464 22420 2470 22432
rect 2866 22420 2872 22432
rect 2464 22392 2872 22420
rect 2464 22380 2470 22392
rect 2866 22380 2872 22392
rect 2924 22380 2930 22432
rect 3234 22380 3240 22432
rect 3292 22380 3298 22432
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 4448 22420 4476 22460
rect 3568 22392 4476 22420
rect 5368 22420 5396 22460
rect 5442 22448 5448 22500
rect 5500 22488 5506 22500
rect 5644 22488 5672 22519
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7374 22556 7380 22568
rect 7024 22528 7380 22556
rect 5500 22460 5672 22488
rect 6012 22488 6040 22516
rect 7024 22488 7052 22528
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 7742 22516 7748 22568
rect 7800 22516 7806 22568
rect 9232 22556 9260 22664
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 10686 22652 10692 22704
rect 10744 22692 10750 22704
rect 13354 22692 13360 22704
rect 10744 22664 13360 22692
rect 10744 22652 10750 22664
rect 9585 22627 9643 22633
rect 9585 22593 9597 22627
rect 9631 22624 9643 22627
rect 9674 22624 9680 22636
rect 9631 22596 9680 22624
rect 9631 22593 9643 22596
rect 9585 22587 9643 22593
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 9852 22627 9910 22633
rect 9852 22593 9864 22627
rect 9898 22624 9910 22627
rect 10870 22624 10876 22636
rect 9898 22596 10876 22624
rect 9898 22593 9910 22596
rect 9852 22587 9910 22593
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 13004 22633 13032 22664
rect 13354 22652 13360 22664
rect 13412 22652 13418 22704
rect 13630 22652 13636 22704
rect 13688 22652 13694 22704
rect 13849 22695 13907 22701
rect 13849 22661 13861 22695
rect 13895 22692 13907 22695
rect 14182 22692 14188 22704
rect 13895 22664 14188 22692
rect 13895 22661 13907 22664
rect 13849 22655 13907 22661
rect 14182 22652 14188 22664
rect 14240 22692 14246 22704
rect 16574 22692 16580 22704
rect 14240 22664 16580 22692
rect 14240 22652 14246 22664
rect 16574 22652 16580 22664
rect 16632 22652 16638 22704
rect 17494 22652 17500 22704
rect 17552 22692 17558 22704
rect 17681 22695 17739 22701
rect 17681 22692 17693 22695
rect 17552 22664 17693 22692
rect 17552 22652 17558 22664
rect 17681 22661 17693 22664
rect 17727 22661 17739 22695
rect 17972 22692 18000 22720
rect 17681 22655 17739 22661
rect 17896 22664 18000 22692
rect 17896 22661 17969 22664
rect 12621 22627 12679 22633
rect 12621 22624 12633 22627
rect 12584 22596 12633 22624
rect 12584 22584 12590 22596
rect 12621 22593 12633 22596
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22593 13047 22627
rect 13372 22624 13400 22652
rect 14458 22624 14464 22636
rect 13372 22596 14464 22624
rect 12989 22587 13047 22593
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22624 15623 22627
rect 15654 22624 15660 22636
rect 15611 22596 15660 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 15749 22627 15807 22633
rect 15749 22593 15761 22627
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 8036 22528 9260 22556
rect 12253 22559 12311 22565
rect 6012 22460 7052 22488
rect 5500 22448 5506 22460
rect 7190 22448 7196 22500
rect 7248 22448 7254 22500
rect 8036 22497 8064 22528
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 13354 22556 13360 22568
rect 12299 22528 13360 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 13814 22516 13820 22568
rect 13872 22556 13878 22568
rect 15289 22559 15347 22565
rect 15289 22556 15301 22559
rect 13872 22528 15301 22556
rect 13872 22516 13878 22528
rect 15289 22525 15301 22528
rect 15335 22525 15347 22559
rect 15764 22556 15792 22587
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16390 22624 16396 22636
rect 16080 22596 16396 22624
rect 16080 22584 16086 22596
rect 16390 22584 16396 22596
rect 16448 22584 16454 22636
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 17770 22624 17776 22636
rect 17092 22596 17776 22624
rect 17092 22584 17098 22596
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 17896 22630 17923 22661
rect 17911 22627 17923 22630
rect 17957 22627 17969 22661
rect 18046 22652 18052 22704
rect 18104 22692 18110 22704
rect 18690 22692 18696 22704
rect 18104 22664 18696 22692
rect 18104 22652 18110 22664
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 17911 22621 17969 22627
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18288 22596 18521 22624
rect 18288 22584 18294 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18874 22584 18880 22636
rect 18932 22584 18938 22636
rect 17402 22556 17408 22568
rect 15289 22519 15347 22525
rect 15488 22528 15700 22556
rect 15764 22528 17408 22556
rect 8021 22491 8079 22497
rect 8021 22457 8033 22491
rect 8067 22457 8079 22491
rect 8021 22451 8079 22457
rect 9033 22491 9091 22497
rect 9033 22457 9045 22491
rect 9079 22457 9091 22491
rect 9033 22451 9091 22457
rect 6730 22420 6736 22432
rect 5368 22392 6736 22420
rect 3568 22380 3574 22392
rect 6730 22380 6736 22392
rect 6788 22380 6794 22432
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 8205 22423 8263 22429
rect 8205 22420 8217 22423
rect 7156 22392 8217 22420
rect 7156 22380 7162 22392
rect 8205 22389 8217 22392
rect 8251 22389 8263 22423
rect 9048 22420 9076 22451
rect 10686 22448 10692 22500
rect 10744 22488 10750 22500
rect 15488 22497 15516 22528
rect 12713 22491 12771 22497
rect 12713 22488 12725 22491
rect 10744 22460 12725 22488
rect 10744 22448 10750 22460
rect 12713 22457 12725 22460
rect 12759 22457 12771 22491
rect 12713 22451 12771 22457
rect 14001 22491 14059 22497
rect 14001 22457 14013 22491
rect 14047 22488 14059 22491
rect 15381 22491 15439 22497
rect 15381 22488 15393 22491
rect 14047 22460 15393 22488
rect 14047 22457 14059 22460
rect 14001 22451 14059 22457
rect 15381 22457 15393 22460
rect 15427 22457 15439 22491
rect 15381 22451 15439 22457
rect 15473 22491 15531 22497
rect 15473 22457 15485 22491
rect 15519 22457 15531 22491
rect 15672 22488 15700 22528
rect 17402 22516 17408 22528
rect 17460 22516 17466 22568
rect 19076 22556 19104 22732
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 19705 22763 19763 22769
rect 19705 22729 19717 22763
rect 19751 22760 19763 22763
rect 20622 22760 20628 22772
rect 19751 22732 20628 22760
rect 19751 22729 19763 22732
rect 19705 22723 19763 22729
rect 20622 22720 20628 22732
rect 20680 22720 20686 22772
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22760 21051 22763
rect 22554 22760 22560 22772
rect 21039 22732 22560 22760
rect 21039 22729 21051 22732
rect 20993 22723 21051 22729
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 22830 22720 22836 22772
rect 22888 22760 22894 22772
rect 23106 22760 23112 22772
rect 22888 22732 23112 22760
rect 22888 22720 22894 22732
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 26605 22763 26663 22769
rect 26605 22760 26617 22763
rect 23492 22732 26617 22760
rect 19521 22695 19579 22701
rect 19521 22692 19533 22695
rect 19444 22664 19533 22692
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 19208 22596 19349 22624
rect 19208 22584 19214 22596
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 17788 22528 19104 22556
rect 17586 22488 17592 22500
rect 15672 22460 17592 22488
rect 15473 22451 15531 22457
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 9950 22420 9956 22432
rect 9048 22392 9956 22420
rect 8205 22383 8263 22389
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 12526 22380 12532 22432
rect 12584 22380 12590 22432
rect 13817 22423 13875 22429
rect 13817 22389 13829 22423
rect 13863 22420 13875 22423
rect 13906 22420 13912 22432
rect 13863 22392 13912 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 15010 22380 15016 22432
rect 15068 22380 15074 22432
rect 15654 22380 15660 22432
rect 15712 22420 15718 22432
rect 17788 22420 17816 22528
rect 18506 22488 18512 22500
rect 17880 22460 18512 22488
rect 17880 22429 17908 22460
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 19150 22488 19156 22500
rect 18800 22460 19156 22488
rect 15712 22392 17816 22420
rect 17865 22423 17923 22429
rect 15712 22380 15718 22392
rect 17865 22389 17877 22423
rect 17911 22389 17923 22423
rect 17865 22383 17923 22389
rect 18046 22380 18052 22432
rect 18104 22380 18110 22432
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 18800 22420 18828 22460
rect 19150 22448 19156 22460
rect 19208 22448 19214 22500
rect 19444 22488 19472 22664
rect 19521 22661 19533 22664
rect 19567 22661 19579 22695
rect 19521 22655 19579 22661
rect 19610 22652 19616 22704
rect 19668 22692 19674 22704
rect 20165 22695 20223 22701
rect 20165 22692 20177 22695
rect 19668 22664 20177 22692
rect 19668 22652 19674 22664
rect 20165 22661 20177 22664
rect 20211 22692 20223 22695
rect 20438 22692 20444 22704
rect 20211 22664 20444 22692
rect 20211 22661 20223 22664
rect 20165 22655 20223 22661
rect 20438 22652 20444 22664
rect 20496 22652 20502 22704
rect 20530 22652 20536 22704
rect 20588 22652 20594 22704
rect 21634 22652 21640 22704
rect 21692 22692 21698 22704
rect 23492 22692 23520 22732
rect 26605 22729 26617 22732
rect 26651 22729 26663 22763
rect 26605 22723 26663 22729
rect 21692 22664 23520 22692
rect 21692 22652 21698 22664
rect 23566 22652 23572 22704
rect 23624 22692 23630 22704
rect 25470 22695 25528 22701
rect 25470 22692 25482 22695
rect 23624 22664 25482 22692
rect 23624 22652 23630 22664
rect 25470 22661 25482 22664
rect 25516 22661 25528 22695
rect 25470 22655 25528 22661
rect 19702 22584 19708 22636
rect 19760 22624 19766 22636
rect 20349 22627 20407 22633
rect 20349 22624 20361 22627
rect 19760 22596 20361 22624
rect 19760 22584 19766 22596
rect 20349 22593 20361 22596
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 21177 22627 21235 22633
rect 21177 22624 21189 22627
rect 20772 22596 21189 22624
rect 20772 22584 20778 22596
rect 21177 22593 21189 22596
rect 21223 22593 21235 22627
rect 21177 22587 21235 22593
rect 22186 22584 22192 22636
rect 22244 22584 22250 22636
rect 22554 22584 22560 22636
rect 22612 22624 22618 22636
rect 22997 22627 23055 22633
rect 22997 22624 23009 22627
rect 22612 22596 23009 22624
rect 22612 22584 22618 22596
rect 22997 22593 23009 22596
rect 23043 22593 23055 22627
rect 22997 22587 23055 22593
rect 24578 22584 24584 22636
rect 24636 22584 24642 22636
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 25225 22627 25283 22633
rect 25225 22624 25237 22627
rect 25188 22596 25237 22624
rect 25188 22584 25194 22596
rect 25225 22593 25237 22596
rect 25271 22593 25283 22627
rect 25958 22624 25964 22636
rect 25225 22587 25283 22593
rect 25332 22596 25964 22624
rect 22738 22516 22744 22568
rect 22796 22516 22802 22568
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25332 22556 25360 22596
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 24912 22528 25360 22556
rect 24912 22516 24918 22528
rect 19306 22460 22508 22488
rect 18196 22392 18828 22420
rect 18196 22380 18202 22392
rect 19058 22380 19064 22432
rect 19116 22420 19122 22432
rect 19306 22420 19334 22460
rect 19116 22392 19334 22420
rect 22005 22423 22063 22429
rect 19116 22380 19122 22392
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22370 22420 22376 22432
rect 22051 22392 22376 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 22480 22420 22508 22460
rect 24670 22448 24676 22500
rect 24728 22448 24734 22500
rect 23382 22420 23388 22432
rect 22480 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 24121 22423 24179 22429
rect 24121 22389 24133 22423
rect 24167 22420 24179 22423
rect 24302 22420 24308 22432
rect 24167 22392 24308 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 24302 22380 24308 22392
rect 24360 22380 24366 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 2866 22176 2872 22228
rect 2924 22176 2930 22228
rect 3237 22219 3295 22225
rect 3237 22185 3249 22219
rect 3283 22216 3295 22219
rect 3694 22216 3700 22228
rect 3283 22188 3700 22216
rect 3283 22185 3295 22188
rect 3237 22179 3295 22185
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 5074 22216 5080 22228
rect 4764 22188 5080 22216
rect 4764 22176 4770 22188
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 6914 22216 6920 22228
rect 5408 22188 6920 22216
rect 5408 22176 5414 22188
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 8113 22219 8171 22225
rect 8113 22216 8125 22219
rect 7708 22188 8125 22216
rect 7708 22176 7714 22188
rect 8113 22185 8125 22188
rect 8159 22185 8171 22219
rect 8113 22179 8171 22185
rect 8386 22176 8392 22228
rect 8444 22216 8450 22228
rect 9585 22219 9643 22225
rect 9585 22216 9597 22219
rect 8444 22188 9597 22216
rect 8444 22176 8450 22188
rect 9585 22185 9597 22188
rect 9631 22185 9643 22219
rect 9585 22179 9643 22185
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 1544 22052 1992 22080
rect 1544 22040 1550 22052
rect 1762 21972 1768 22024
rect 1820 21972 1826 22024
rect 1854 21972 1860 22024
rect 1912 21972 1918 22024
rect 1964 22021 1992 22052
rect 1964 22015 2047 22021
rect 1964 21984 2001 22015
rect 1989 21981 2001 21984
rect 2035 21981 2047 22015
rect 1989 21975 2047 21981
rect 2130 21972 2136 22024
rect 2188 21972 2194 22024
rect 2593 22015 2651 22021
rect 2593 22012 2605 22015
rect 2332 21984 2605 22012
rect 566 21904 572 21956
rect 624 21944 630 21956
rect 1581 21947 1639 21953
rect 1581 21944 1593 21947
rect 624 21916 1593 21944
rect 624 21904 630 21916
rect 1581 21913 1593 21916
rect 1627 21913 1639 21947
rect 1872 21944 1900 21972
rect 2332 21944 2360 21984
rect 2593 21981 2605 21984
rect 2639 21981 2651 22015
rect 2593 21975 2651 21981
rect 2682 21972 2688 22024
rect 2740 21972 2746 22024
rect 2884 21953 2912 22176
rect 7193 22151 7251 22157
rect 7193 22117 7205 22151
rect 7239 22148 7251 22151
rect 7374 22148 7380 22160
rect 7239 22120 7380 22148
rect 7239 22117 7251 22120
rect 7193 22111 7251 22117
rect 7374 22108 7380 22120
rect 7432 22148 7438 22160
rect 9600 22148 9628 22179
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 11330 22216 11336 22228
rect 10836 22188 11336 22216
rect 10836 22176 10842 22188
rect 11330 22176 11336 22188
rect 11388 22176 11394 22228
rect 13078 22176 13084 22228
rect 13136 22216 13142 22228
rect 13357 22219 13415 22225
rect 13357 22216 13369 22219
rect 13136 22188 13369 22216
rect 13136 22176 13142 22188
rect 13357 22185 13369 22188
rect 13403 22185 13415 22219
rect 13357 22179 13415 22185
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17405 22219 17463 22225
rect 17405 22216 17417 22219
rect 17276 22188 17417 22216
rect 17276 22176 17282 22188
rect 17405 22185 17417 22188
rect 17451 22185 17463 22219
rect 17405 22179 17463 22185
rect 17586 22176 17592 22228
rect 17644 22176 17650 22228
rect 18138 22216 18144 22228
rect 17972 22188 18144 22216
rect 10318 22148 10324 22160
rect 7432 22120 8708 22148
rect 9600 22120 10324 22148
rect 7432 22108 7438 22120
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 4249 22083 4307 22089
rect 4249 22080 4261 22083
rect 3844 22052 4261 22080
rect 3844 22040 3850 22052
rect 4249 22049 4261 22052
rect 4295 22049 4307 22083
rect 5350 22080 5356 22092
rect 4249 22043 4307 22049
rect 4356 22052 5356 22080
rect 3099 22015 3157 22021
rect 3099 21981 3111 22015
rect 3145 22012 3157 22015
rect 4356 22012 4384 22052
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 5629 22083 5687 22089
rect 5629 22049 5641 22083
rect 5675 22080 5687 22083
rect 5902 22080 5908 22092
rect 5675 22052 5908 22080
rect 5675 22049 5687 22052
rect 5629 22043 5687 22049
rect 5902 22040 5908 22052
rect 5960 22040 5966 22092
rect 6914 22040 6920 22092
rect 6972 22080 6978 22092
rect 6972 22052 8616 22080
rect 6972 22040 6978 22052
rect 3145 21984 4384 22012
rect 4433 22015 4491 22021
rect 3145 21981 3157 21984
rect 3099 21975 3157 21981
rect 3252 21956 3280 21984
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4798 22012 4804 22024
rect 4479 21984 4804 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 5132 21984 5549 22012
rect 5132 21972 5138 21984
rect 5537 21981 5549 21984
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 1872 21916 2360 21944
rect 2869 21947 2927 21953
rect 1581 21907 1639 21913
rect 2869 21913 2881 21947
rect 2915 21913 2927 21947
rect 2869 21907 2927 21913
rect 2961 21947 3019 21953
rect 2961 21913 2973 21947
rect 3007 21944 3019 21947
rect 3007 21916 3096 21944
rect 3007 21913 3019 21916
rect 2961 21907 3019 21913
rect 3068 21888 3096 21916
rect 3234 21904 3240 21956
rect 3292 21904 3298 21956
rect 4338 21904 4344 21956
rect 4396 21944 4402 21956
rect 4617 21947 4675 21953
rect 4617 21944 4629 21947
rect 4396 21916 4629 21944
rect 4396 21904 4402 21916
rect 4617 21913 4629 21916
rect 4663 21913 4675 21947
rect 4617 21907 4675 21913
rect 4709 21947 4767 21953
rect 4709 21913 4721 21947
rect 4755 21944 4767 21947
rect 4890 21944 4896 21956
rect 4755 21916 4896 21944
rect 4755 21913 4767 21916
rect 4709 21907 4767 21913
rect 4890 21904 4896 21916
rect 4948 21904 4954 21956
rect 1857 21879 1915 21885
rect 1857 21845 1869 21879
rect 1903 21876 1915 21879
rect 2222 21876 2228 21888
rect 1903 21848 2228 21876
rect 1903 21845 1915 21848
rect 1857 21839 1915 21845
rect 2222 21836 2228 21848
rect 2280 21836 2286 21888
rect 3050 21836 3056 21888
rect 3108 21836 3114 21888
rect 5350 21836 5356 21888
rect 5408 21836 5414 21888
rect 5534 21836 5540 21888
rect 5592 21876 5598 21888
rect 5736 21876 5764 21975
rect 5810 21972 5816 22024
rect 5868 21972 5874 22024
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 22012 6883 22015
rect 7098 22012 7104 22024
rect 6871 21984 7104 22012
rect 6871 21981 6883 21984
rect 6825 21975 6883 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8386 22012 8392 22024
rect 8343 21984 8392 22012
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 8588 22021 8616 22052
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 6454 21904 6460 21956
rect 6512 21944 6518 21956
rect 6638 21944 6644 21956
rect 6512 21916 6644 21944
rect 6512 21904 6518 21916
rect 6638 21904 6644 21916
rect 6696 21944 6702 21956
rect 7009 21947 7067 21953
rect 7009 21944 7021 21947
rect 6696 21916 7021 21944
rect 6696 21904 6702 21916
rect 7009 21913 7021 21916
rect 7055 21913 7067 21947
rect 8680 21944 8708 22120
rect 10318 22108 10324 22120
rect 10376 22148 10382 22160
rect 10962 22148 10968 22160
rect 10376 22120 10968 22148
rect 10376 22108 10382 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 14734 22108 14740 22160
rect 14792 22108 14798 22160
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 17972 22148 18000 22188
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 18598 22176 18604 22228
rect 18656 22216 18662 22228
rect 18966 22216 18972 22228
rect 18656 22188 18972 22216
rect 18656 22176 18662 22188
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 19092 22188 19380 22216
rect 19092 22148 19120 22188
rect 15160 22120 18000 22148
rect 18892 22120 19120 22148
rect 19352 22148 19380 22188
rect 19426 22176 19432 22228
rect 19484 22176 19490 22228
rect 19518 22176 19524 22228
rect 19576 22176 19582 22228
rect 19702 22176 19708 22228
rect 19760 22216 19766 22228
rect 24854 22216 24860 22228
rect 19760 22188 24860 22216
rect 19760 22176 19766 22188
rect 24854 22176 24860 22188
rect 24912 22176 24918 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 25188 22188 25912 22216
rect 25188 22176 25194 22188
rect 19536 22148 19564 22176
rect 19352 22120 19564 22148
rect 15160 22108 15166 22120
rect 18892 22094 18920 22120
rect 21634 22108 21640 22160
rect 21692 22148 21698 22160
rect 21913 22151 21971 22157
rect 21913 22148 21925 22151
rect 21692 22120 21925 22148
rect 21692 22108 21698 22120
rect 21913 22117 21925 22120
rect 21959 22117 21971 22151
rect 25884 22148 25912 22188
rect 25884 22120 26004 22148
rect 21913 22111 21971 22117
rect 8846 22040 8852 22092
rect 8904 22080 8910 22092
rect 9125 22083 9183 22089
rect 9125 22080 9137 22083
rect 8904 22052 9137 22080
rect 8904 22040 8910 22052
rect 9125 22049 9137 22052
rect 9171 22080 9183 22083
rect 12713 22083 12771 22089
rect 9171 22052 10180 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 10152 22024 10180 22052
rect 12713 22049 12725 22083
rect 12759 22080 12771 22083
rect 13262 22080 13268 22092
rect 12759 22052 13268 22080
rect 12759 22049 12771 22052
rect 12713 22043 12771 22049
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 16022 22040 16028 22092
rect 16080 22080 16086 22092
rect 18616 22080 18920 22094
rect 16080 22052 16436 22080
rect 16080 22040 16086 22052
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 22012 9551 22015
rect 9858 22012 9864 22024
rect 9539 21984 9864 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 10192 21984 10425 22012
rect 10192 21972 10198 21984
rect 10413 21981 10425 21984
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 9766 21944 9772 21956
rect 8680 21916 9772 21944
rect 7009 21907 7067 21913
rect 9766 21904 9772 21916
rect 9824 21904 9830 21956
rect 9876 21944 9904 21972
rect 10612 21944 10640 21975
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11057 22015 11115 22021
rect 11057 22012 11069 22015
rect 11020 21984 11069 22012
rect 11020 21972 11026 21984
rect 11057 21981 11069 21984
rect 11103 21981 11115 22015
rect 12986 22012 12992 22024
rect 11057 21975 11115 21981
rect 12360 21984 12992 22012
rect 9876 21916 10640 21944
rect 12158 21904 12164 21956
rect 12216 21944 12222 21956
rect 12360 21953 12388 21984
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 13596 21984 14565 22012
rect 13596 21972 13602 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 16408 22021 16436 22052
rect 16500 22066 18920 22080
rect 16500 22052 18644 22066
rect 16500 22021 16528 22052
rect 18966 22040 18972 22092
rect 19024 22080 19030 22092
rect 20806 22080 20812 22092
rect 19024 22052 20812 22080
rect 19024 22040 19030 22052
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 21082 22040 21088 22092
rect 21140 22040 21146 22092
rect 22572 22052 22784 22080
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 14700 21984 16221 22012
rect 14700 21972 14706 21984
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12216 21916 12357 21944
rect 12216 21904 12222 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 12529 21947 12587 21953
rect 12529 21913 12541 21947
rect 12575 21944 12587 21947
rect 12802 21944 12808 21956
rect 12575 21916 12808 21944
rect 12575 21913 12587 21916
rect 12529 21907 12587 21913
rect 12802 21904 12808 21916
rect 12860 21904 12866 21956
rect 13173 21947 13231 21953
rect 13173 21913 13185 21947
rect 13219 21944 13231 21947
rect 15381 21947 15439 21953
rect 13219 21916 15240 21944
rect 13219 21913 13231 21916
rect 13173 21907 13231 21913
rect 15212 21888 15240 21916
rect 15381 21913 15393 21947
rect 15427 21944 15439 21947
rect 15746 21944 15752 21956
rect 15427 21916 15752 21944
rect 15427 21913 15439 21916
rect 15381 21907 15439 21913
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 16224 21944 16252 21975
rect 16574 21972 16580 22024
rect 16632 21972 16638 22024
rect 16684 21984 17356 22012
rect 16684 21944 16712 21984
rect 16224 21916 16712 21944
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 17221 21947 17279 21953
rect 17221 21944 17233 21947
rect 17184 21916 17233 21944
rect 17184 21904 17190 21916
rect 17221 21913 17233 21916
rect 17267 21913 17279 21947
rect 17328 21944 17356 21984
rect 18230 21972 18236 22024
rect 18288 21972 18294 22024
rect 18874 21972 18880 22024
rect 18932 21972 18938 22024
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 19392 21984 19625 22012
rect 19392 21972 19398 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 20257 22015 20315 22021
rect 20257 22012 20269 22015
rect 19760 21984 20269 22012
rect 19760 21972 19766 21984
rect 20257 21981 20269 21984
rect 20303 21981 20315 22015
rect 22572 22012 22600 22052
rect 20257 21975 20315 21981
rect 20364 21984 22600 22012
rect 18598 21944 18604 21956
rect 17328 21916 18604 21944
rect 17221 21907 17279 21913
rect 18598 21904 18604 21916
rect 18656 21904 18662 21956
rect 20364 21944 20392 21984
rect 22646 21972 22652 22024
rect 22704 21972 22710 22024
rect 22756 22012 22784 22052
rect 24118 22040 24124 22092
rect 24176 22080 24182 22092
rect 25976 22080 26004 22120
rect 26789 22083 26847 22089
rect 26789 22080 26801 22083
rect 24176 22052 25084 22080
rect 25976 22052 26801 22080
rect 24176 22040 24182 22052
rect 22756 21984 23040 22012
rect 18708 21916 20392 21944
rect 5592 21848 5764 21876
rect 5592 21836 5598 21848
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 9306 21876 9312 21888
rect 6604 21848 9312 21876
rect 6604 21836 6610 21848
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 9548 21848 10609 21876
rect 9548 21836 9554 21848
rect 10597 21845 10609 21848
rect 10643 21845 10655 21879
rect 10597 21839 10655 21845
rect 13354 21836 13360 21888
rect 13412 21885 13418 21888
rect 13412 21879 13431 21885
rect 13419 21845 13431 21879
rect 13412 21839 13431 21845
rect 13541 21879 13599 21885
rect 13541 21845 13553 21879
rect 13587 21876 13599 21879
rect 13814 21876 13820 21888
rect 13587 21848 13820 21876
rect 13587 21845 13599 21848
rect 13541 21839 13599 21845
rect 13412 21836 13418 21839
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 15102 21876 15108 21888
rect 14700 21848 15108 21876
rect 14700 21836 14706 21848
rect 15102 21836 15108 21848
rect 15160 21836 15166 21888
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 15252 21848 15485 21876
rect 15252 21836 15258 21848
rect 15473 21845 15485 21848
rect 15519 21876 15531 21879
rect 16022 21876 16028 21888
rect 15519 21848 16028 21876
rect 15519 21845 15531 21848
rect 15473 21839 15531 21845
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 16758 21836 16764 21888
rect 16816 21836 16822 21888
rect 17402 21836 17408 21888
rect 17460 21885 17466 21888
rect 17460 21879 17479 21885
rect 17467 21845 17479 21879
rect 17460 21839 17479 21845
rect 18049 21879 18107 21885
rect 18049 21845 18061 21879
rect 18095 21876 18107 21879
rect 18322 21876 18328 21888
rect 18095 21848 18328 21876
rect 18095 21845 18107 21848
rect 18049 21839 18107 21845
rect 17460 21836 17466 21839
rect 18322 21836 18328 21848
rect 18380 21836 18386 21888
rect 18708 21885 18736 21916
rect 20438 21904 20444 21956
rect 20496 21944 20502 21956
rect 20717 21947 20775 21953
rect 20717 21944 20729 21947
rect 20496 21916 20729 21944
rect 20496 21904 20502 21916
rect 20717 21913 20729 21916
rect 20763 21913 20775 21947
rect 20717 21907 20775 21913
rect 20898 21904 20904 21956
rect 20956 21904 20962 21956
rect 21450 21904 21456 21956
rect 21508 21944 21514 21956
rect 21637 21947 21695 21953
rect 21637 21944 21649 21947
rect 21508 21916 21649 21944
rect 21508 21904 21514 21916
rect 21637 21913 21649 21916
rect 21683 21913 21695 21947
rect 22894 21947 22952 21953
rect 22894 21944 22906 21947
rect 21637 21907 21695 21913
rect 21744 21916 22906 21944
rect 18693 21879 18751 21885
rect 18693 21845 18705 21879
rect 18739 21845 18751 21879
rect 18693 21839 18751 21845
rect 20073 21879 20131 21885
rect 20073 21845 20085 21879
rect 20119 21876 20131 21879
rect 21744 21876 21772 21916
rect 22894 21913 22906 21916
rect 22940 21913 22952 21947
rect 23012 21944 23040 21984
rect 24946 21972 24952 22024
rect 25004 21972 25010 22024
rect 25056 22012 25084 22052
rect 26789 22049 26801 22052
rect 26835 22049 26847 22083
rect 26789 22043 26847 22049
rect 27045 22015 27103 22021
rect 27045 22012 27057 22015
rect 25056 21984 27057 22012
rect 27045 21981 27057 21984
rect 27091 21981 27103 22015
rect 27045 21975 27103 21981
rect 25194 21947 25252 21953
rect 25194 21944 25206 21947
rect 23012 21916 25206 21944
rect 22894 21907 22952 21913
rect 25194 21913 25206 21916
rect 25240 21913 25252 21947
rect 25194 21907 25252 21913
rect 20119 21848 21772 21876
rect 22097 21879 22155 21885
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 23750 21876 23756 21888
rect 22143 21848 23756 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 23842 21836 23848 21888
rect 23900 21876 23906 21888
rect 24029 21879 24087 21885
rect 24029 21876 24041 21879
rect 23900 21848 24041 21876
rect 23900 21836 23906 21848
rect 24029 21845 24041 21848
rect 24075 21845 24087 21879
rect 24029 21839 24087 21845
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 26329 21879 26387 21885
rect 26329 21876 26341 21879
rect 24728 21848 26341 21876
rect 24728 21836 24734 21848
rect 26329 21845 26341 21848
rect 26375 21845 26387 21879
rect 26329 21839 26387 21845
rect 28166 21836 28172 21888
rect 28224 21836 28230 21888
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 3602 21632 3608 21684
rect 3660 21672 3666 21684
rect 3789 21675 3847 21681
rect 3789 21672 3801 21675
rect 3660 21644 3801 21672
rect 3660 21632 3666 21644
rect 3789 21641 3801 21644
rect 3835 21641 3847 21675
rect 3789 21635 3847 21641
rect 4985 21675 5043 21681
rect 4985 21641 4997 21675
rect 5031 21672 5043 21675
rect 5258 21672 5264 21684
rect 5031 21644 5264 21672
rect 5031 21641 5043 21644
rect 4985 21635 5043 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 6270 21632 6276 21684
rect 6328 21672 6334 21684
rect 7650 21672 7656 21684
rect 6328 21644 7656 21672
rect 6328 21632 6334 21644
rect 7650 21632 7656 21644
rect 7708 21672 7714 21684
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 7708 21644 7941 21672
rect 7708 21632 7714 21644
rect 7929 21641 7941 21644
rect 7975 21641 7987 21675
rect 9950 21672 9956 21684
rect 7929 21635 7987 21641
rect 9048 21644 9956 21672
rect 1762 21564 1768 21616
rect 1820 21564 1826 21616
rect 4890 21564 4896 21616
rect 4948 21604 4954 21616
rect 6638 21604 6644 21616
rect 4948 21576 6644 21604
rect 4948 21564 4954 21576
rect 6638 21564 6644 21576
rect 6696 21564 6702 21616
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 7837 21607 7895 21613
rect 7837 21604 7849 21607
rect 6788 21576 7849 21604
rect 6788 21564 6794 21576
rect 7837 21573 7849 21576
rect 7883 21573 7895 21607
rect 7837 21567 7895 21573
rect 1780 21536 1808 21564
rect 2041 21539 2099 21545
rect 2041 21536 2053 21539
rect 1780 21508 2053 21536
rect 2041 21505 2053 21508
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 2222 21496 2228 21548
rect 2280 21496 2286 21548
rect 2498 21496 2504 21548
rect 2556 21496 2562 21548
rect 3050 21496 3056 21548
rect 3108 21496 3114 21548
rect 4154 21496 4160 21548
rect 4212 21496 4218 21548
rect 4246 21496 4252 21548
rect 4304 21496 4310 21548
rect 5166 21496 5172 21548
rect 5224 21536 5230 21548
rect 5261 21539 5319 21545
rect 5261 21536 5273 21539
rect 5224 21508 5273 21536
rect 5224 21496 5230 21508
rect 5261 21505 5273 21508
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 474 21428 480 21480
rect 532 21468 538 21480
rect 1581 21471 1639 21477
rect 1581 21468 1593 21471
rect 532 21440 1593 21468
rect 532 21428 538 21440
rect 1581 21437 1593 21440
rect 1627 21437 1639 21471
rect 1581 21431 1639 21437
rect 1762 21428 1768 21480
rect 1820 21468 1826 21480
rect 2685 21471 2743 21477
rect 2685 21468 2697 21471
rect 1820 21440 2697 21468
rect 1820 21428 1826 21440
rect 2685 21437 2697 21440
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 3970 21428 3976 21480
rect 4028 21428 4034 21480
rect 5368 21468 5396 21499
rect 5442 21496 5448 21548
rect 5500 21496 5506 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 5810 21536 5816 21548
rect 5675 21508 5816 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 6914 21496 6920 21548
rect 6972 21496 6978 21548
rect 7098 21496 7104 21548
rect 7156 21496 7162 21548
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 8754 21536 8760 21548
rect 7800 21508 8760 21536
rect 7800 21496 7806 21508
rect 8754 21496 8760 21508
rect 8812 21536 8818 21548
rect 9048 21545 9076 21644
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10413 21675 10471 21681
rect 10060 21644 10364 21672
rect 10060 21613 10088 21644
rect 10045 21607 10103 21613
rect 10045 21573 10057 21607
rect 10091 21573 10103 21607
rect 10245 21607 10303 21613
rect 10245 21604 10257 21607
rect 10045 21567 10103 21573
rect 10244 21573 10257 21604
rect 10291 21573 10303 21607
rect 10336 21604 10364 21644
rect 10413 21641 10425 21675
rect 10459 21672 10471 21675
rect 10686 21672 10692 21684
rect 10459 21644 10692 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 10778 21632 10784 21684
rect 10836 21672 10842 21684
rect 10836 21644 12434 21672
rect 10836 21632 10842 21644
rect 11054 21604 11060 21616
rect 10336 21576 11060 21604
rect 10244 21567 10303 21573
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8812 21508 9045 21536
rect 8812 21496 8818 21508
rect 9033 21505 9045 21508
rect 9079 21505 9091 21539
rect 10244 21536 10272 21567
rect 11054 21564 11060 21576
rect 11112 21564 11118 21616
rect 11146 21564 11152 21616
rect 11204 21604 11210 21616
rect 11977 21607 12035 21613
rect 11977 21604 11989 21607
rect 11204 21576 11989 21604
rect 11204 21564 11210 21576
rect 11977 21573 11989 21576
rect 12023 21573 12035 21607
rect 12406 21604 12434 21644
rect 12710 21632 12716 21684
rect 12768 21632 12774 21684
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 14737 21675 14795 21681
rect 14737 21672 14749 21675
rect 12952 21644 14749 21672
rect 12952 21632 12958 21644
rect 14737 21641 14749 21644
rect 14783 21641 14795 21675
rect 14737 21635 14795 21641
rect 15838 21632 15844 21684
rect 15896 21632 15902 21684
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 18414 21672 18420 21684
rect 16264 21644 17264 21672
rect 16264 21632 16270 21644
rect 17236 21616 17264 21644
rect 17972 21644 18420 21672
rect 14274 21604 14280 21616
rect 12406 21576 14280 21604
rect 11977 21567 12035 21573
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 15746 21564 15752 21616
rect 15804 21604 15810 21616
rect 16853 21607 16911 21613
rect 16853 21604 16865 21607
rect 15804 21576 16865 21604
rect 15804 21564 15810 21576
rect 16853 21573 16865 21576
rect 16899 21573 16911 21607
rect 16853 21567 16911 21573
rect 16942 21564 16948 21616
rect 17000 21604 17006 21616
rect 17053 21607 17111 21613
rect 17053 21604 17065 21607
rect 17000 21576 17065 21604
rect 17000 21564 17006 21576
rect 17053 21573 17065 21576
rect 17099 21573 17111 21607
rect 17053 21567 17111 21573
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17681 21607 17739 21613
rect 17681 21604 17693 21607
rect 17276 21576 17693 21604
rect 17276 21564 17282 21576
rect 17681 21573 17693 21576
rect 17727 21573 17739 21607
rect 17681 21567 17739 21573
rect 17881 21607 17939 21613
rect 17881 21573 17893 21607
rect 17927 21604 17939 21607
rect 17972 21604 18000 21644
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19702 21632 19708 21684
rect 19760 21632 19766 21684
rect 20625 21675 20683 21681
rect 20625 21641 20637 21675
rect 20671 21672 20683 21675
rect 22186 21672 22192 21684
rect 20671 21644 22192 21672
rect 20671 21641 20683 21644
rect 20625 21635 20683 21641
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22336 21644 22477 21672
rect 22336 21632 22342 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 22925 21675 22983 21681
rect 22925 21641 22937 21675
rect 22971 21672 22983 21675
rect 26234 21672 26240 21684
rect 22971 21644 26240 21672
rect 22971 21641 22983 21644
rect 22925 21635 22983 21641
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 17927 21576 18000 21604
rect 17927 21573 17939 21576
rect 17881 21567 17939 21573
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 18509 21607 18567 21613
rect 18509 21604 18521 21607
rect 18196 21576 18521 21604
rect 18196 21564 18202 21576
rect 18509 21573 18521 21576
rect 18555 21573 18567 21607
rect 18709 21607 18767 21613
rect 18709 21604 18721 21607
rect 18509 21567 18567 21573
rect 18616 21576 18721 21604
rect 10686 21536 10692 21548
rect 10244 21508 10692 21536
rect 9033 21499 9091 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 10873 21539 10931 21545
rect 10873 21536 10885 21539
rect 10836 21508 10885 21536
rect 10836 21496 10842 21508
rect 10873 21505 10885 21508
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 11848 21508 11897 21536
rect 11848 21496 11854 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 12434 21536 12440 21548
rect 12115 21508 12440 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 12434 21496 12440 21508
rect 12492 21536 12498 21548
rect 12618 21536 12624 21548
rect 12492 21508 12624 21536
rect 12492 21496 12498 21508
rect 12618 21496 12624 21508
rect 12676 21496 12682 21548
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21505 12955 21539
rect 12897 21499 12955 21505
rect 5534 21468 5540 21480
rect 5368 21440 5540 21468
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21468 9551 21471
rect 12912 21468 12940 21499
rect 12986 21496 12992 21548
rect 13044 21536 13050 21548
rect 13613 21539 13671 21545
rect 13613 21536 13625 21539
rect 13044 21508 13625 21536
rect 13044 21496 13050 21508
rect 13613 21505 13625 21508
rect 13659 21505 13671 21539
rect 13613 21499 13671 21505
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16482 21536 16488 21548
rect 15979 21508 16488 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 17310 21496 17316 21548
rect 17368 21536 17374 21548
rect 18616 21536 18644 21576
rect 18709 21573 18721 21576
rect 18755 21573 18767 21607
rect 18709 21567 18767 21573
rect 19521 21607 19579 21613
rect 19521 21573 19533 21607
rect 19567 21604 19579 21607
rect 19886 21604 19892 21616
rect 19567 21576 19892 21604
rect 19567 21573 19579 21576
rect 19521 21567 19579 21573
rect 19886 21564 19892 21576
rect 19944 21564 19950 21616
rect 23934 21613 23940 21616
rect 23928 21604 23940 21613
rect 23895 21576 23940 21604
rect 23928 21567 23940 21576
rect 23934 21564 23940 21567
rect 23992 21564 23998 21616
rect 24026 21564 24032 21616
rect 24084 21604 24090 21616
rect 25038 21604 25044 21616
rect 24084 21576 25044 21604
rect 24084 21564 24090 21576
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 17368 21508 18644 21536
rect 19337 21539 19395 21545
rect 17368 21496 17374 21508
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 19383 21508 20269 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 20257 21505 20269 21508
rect 20303 21536 20315 21539
rect 20346 21536 20352 21548
rect 20303 21508 20352 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20438 21496 20444 21548
rect 20496 21496 20502 21548
rect 21266 21496 21272 21548
rect 21324 21496 21330 21548
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 23109 21539 23167 21545
rect 23109 21536 23121 21539
rect 21784 21508 23121 21536
rect 21784 21496 21790 21508
rect 23109 21505 23121 21508
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 23348 21508 25697 21536
rect 23348 21496 23354 21508
rect 25685 21505 25697 21508
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 9539 21440 12940 21468
rect 13357 21471 13415 21477
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 13357 21437 13369 21471
rect 13403 21437 13415 21471
rect 13357 21431 13415 21437
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 20990 21468 20996 21480
rect 15611 21440 18092 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 1946 21360 1952 21412
rect 2004 21400 2010 21412
rect 7285 21403 7343 21409
rect 7285 21400 7297 21403
rect 2004 21372 7297 21400
rect 2004 21360 2010 21372
rect 7285 21369 7297 21372
rect 7331 21369 7343 21403
rect 7285 21363 7343 21369
rect 8757 21403 8815 21409
rect 8757 21369 8769 21403
rect 8803 21400 8815 21403
rect 9398 21400 9404 21412
rect 8803 21372 9404 21400
rect 8803 21369 8815 21372
rect 8757 21363 8815 21369
rect 9398 21360 9404 21372
rect 9456 21360 9462 21412
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 9950 21400 9956 21412
rect 9732 21372 9956 21400
rect 9732 21360 9738 21372
rect 9950 21360 9956 21372
rect 10008 21400 10014 21412
rect 13372 21400 13400 21431
rect 18064 21409 18092 21440
rect 18616 21440 20996 21468
rect 15473 21403 15531 21409
rect 15473 21400 15485 21403
rect 10008 21372 13400 21400
rect 14292 21372 15485 21400
rect 10008 21360 10014 21372
rect 1670 21292 1676 21344
rect 1728 21332 1734 21344
rect 6086 21332 6092 21344
rect 1728 21304 6092 21332
rect 1728 21292 1734 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 8294 21332 8300 21344
rect 6972 21304 8300 21332
rect 6972 21292 6978 21304
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 9490 21332 9496 21344
rect 8996 21304 9496 21332
rect 8996 21292 9002 21304
rect 9490 21292 9496 21304
rect 9548 21292 9554 21344
rect 10226 21292 10232 21344
rect 10284 21292 10290 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 10962 21332 10968 21344
rect 10744 21304 10968 21332
rect 10744 21292 10750 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 12066 21332 12072 21344
rect 11112 21304 12072 21332
rect 11112 21292 11118 21304
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 14292 21332 14320 21372
rect 15473 21369 15485 21372
rect 15519 21369 15531 21403
rect 15473 21363 15531 21369
rect 15657 21403 15715 21409
rect 15657 21369 15669 21403
rect 15703 21400 15715 21403
rect 17221 21403 17279 21409
rect 17221 21400 17233 21403
rect 15703 21372 17233 21400
rect 15703 21369 15715 21372
rect 15657 21363 15715 21369
rect 17221 21369 17233 21372
rect 17267 21369 17279 21403
rect 17221 21363 17279 21369
rect 18049 21403 18107 21409
rect 18049 21369 18061 21403
rect 18095 21369 18107 21403
rect 18049 21363 18107 21369
rect 13780 21304 14320 21332
rect 13780 21292 13786 21304
rect 15194 21292 15200 21344
rect 15252 21292 15258 21344
rect 17034 21292 17040 21344
rect 17092 21292 17098 21344
rect 17865 21335 17923 21341
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 18616 21332 18644 21440
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 22005 21471 22063 21477
rect 22005 21437 22017 21471
rect 22051 21468 22063 21471
rect 22094 21468 22100 21480
rect 22051 21440 22100 21468
rect 22051 21437 22063 21440
rect 22005 21431 22063 21437
rect 22094 21428 22100 21440
rect 22152 21428 22158 21480
rect 22204 21440 22416 21468
rect 19150 21400 19156 21412
rect 18708 21372 19156 21400
rect 18708 21341 18736 21372
rect 19150 21360 19156 21372
rect 19208 21360 19214 21412
rect 21085 21403 21143 21409
rect 21085 21369 21097 21403
rect 21131 21400 21143 21403
rect 22204 21400 22232 21440
rect 21131 21372 22232 21400
rect 21131 21369 21143 21372
rect 21085 21363 21143 21369
rect 22278 21360 22284 21412
rect 22336 21360 22342 21412
rect 22388 21400 22416 21440
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 22704 21440 23673 21468
rect 22704 21428 22710 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23474 21400 23480 21412
rect 22388 21372 23480 21400
rect 23474 21360 23480 21372
rect 23532 21360 23538 21412
rect 25590 21400 25596 21412
rect 24964 21372 25596 21400
rect 17911 21304 18644 21332
rect 18693 21335 18751 21341
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 18693 21301 18705 21335
rect 18739 21301 18751 21335
rect 18693 21295 18751 21301
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18840 21304 18889 21332
rect 18840 21292 18846 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 22830 21332 22836 21344
rect 20496 21304 22836 21332
rect 20496 21292 20502 21304
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 23106 21292 23112 21344
rect 23164 21332 23170 21344
rect 24964 21332 24992 21372
rect 25590 21360 25596 21372
rect 25648 21360 25654 21412
rect 23164 21304 24992 21332
rect 23164 21292 23170 21304
rect 25038 21292 25044 21344
rect 25096 21292 25102 21344
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25501 21335 25559 21341
rect 25501 21332 25513 21335
rect 25188 21304 25513 21332
rect 25188 21292 25194 21304
rect 25501 21301 25513 21304
rect 25547 21301 25559 21335
rect 25501 21295 25559 21301
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 2225 21131 2283 21137
rect 2225 21097 2237 21131
rect 2271 21128 2283 21131
rect 2590 21128 2596 21140
rect 2271 21100 2596 21128
rect 2271 21097 2283 21100
rect 2225 21091 2283 21097
rect 2590 21088 2596 21100
rect 2648 21088 2654 21140
rect 3418 21088 3424 21140
rect 3476 21088 3482 21140
rect 4356 21100 5396 21128
rect 2038 21020 2044 21072
rect 2096 21060 2102 21072
rect 3234 21060 3240 21072
rect 2096 21032 3240 21060
rect 2096 21020 2102 21032
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 4154 21020 4160 21072
rect 4212 21060 4218 21072
rect 4356 21069 4384 21100
rect 4341 21063 4399 21069
rect 4341 21060 4353 21063
rect 4212 21032 4353 21060
rect 4212 21020 4218 21032
rect 4341 21029 4353 21032
rect 4387 21029 4399 21063
rect 4341 21023 4399 21029
rect 5258 21020 5264 21072
rect 5316 21020 5322 21072
rect 5368 21060 5396 21100
rect 5442 21088 5448 21140
rect 5500 21088 5506 21140
rect 5997 21131 6055 21137
rect 5997 21097 6009 21131
rect 6043 21128 6055 21131
rect 7006 21128 7012 21140
rect 6043 21100 7012 21128
rect 6043 21097 6055 21100
rect 5997 21091 6055 21097
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 7745 21131 7803 21137
rect 7745 21128 7757 21131
rect 7616 21100 7757 21128
rect 7616 21088 7622 21100
rect 7745 21097 7757 21100
rect 7791 21097 7803 21131
rect 7745 21091 7803 21097
rect 9585 21131 9643 21137
rect 9585 21097 9597 21131
rect 9631 21128 9643 21131
rect 10042 21128 10048 21140
rect 9631 21100 10048 21128
rect 9631 21097 9643 21100
rect 9585 21091 9643 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 12986 21128 12992 21140
rect 10827 21100 12992 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13357 21131 13415 21137
rect 13357 21128 13369 21131
rect 13136 21100 13369 21128
rect 13136 21088 13142 21100
rect 13357 21097 13369 21100
rect 13403 21128 13415 21131
rect 13630 21128 13636 21140
rect 13403 21100 13636 21128
rect 13403 21097 13415 21100
rect 13357 21091 13415 21097
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 14550 21088 14556 21140
rect 14608 21088 14614 21140
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15654 21128 15660 21140
rect 15344 21100 15660 21128
rect 15344 21088 15350 21100
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 16482 21088 16488 21140
rect 16540 21088 16546 21140
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 17954 21128 17960 21140
rect 17635 21100 17960 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 18693 21131 18751 21137
rect 18693 21097 18705 21131
rect 18739 21128 18751 21131
rect 18874 21128 18880 21140
rect 18739 21100 18880 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 21726 21088 21732 21140
rect 21784 21088 21790 21140
rect 22189 21131 22247 21137
rect 22189 21097 22201 21131
rect 22235 21128 22247 21131
rect 22235 21100 23244 21128
rect 22235 21097 22247 21100
rect 22189 21091 22247 21097
rect 5534 21060 5540 21072
rect 5368 21032 5540 21060
rect 5534 21020 5540 21032
rect 5592 21060 5598 21072
rect 6546 21060 6552 21072
rect 5592 21032 6552 21060
rect 5592 21020 5598 21032
rect 6546 21020 6552 21032
rect 6604 21020 6610 21072
rect 7101 21063 7159 21069
rect 7101 21029 7113 21063
rect 7147 21060 7159 21063
rect 9490 21060 9496 21072
rect 7147 21032 9496 21060
rect 7147 21029 7159 21032
rect 7101 21023 7159 21029
rect 9490 21020 9496 21032
rect 9548 21020 9554 21072
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 11793 21063 11851 21069
rect 11793 21060 11805 21063
rect 9732 21032 11805 21060
rect 9732 21020 9738 21032
rect 11793 21029 11805 21032
rect 11839 21029 11851 21063
rect 11793 21023 11851 21029
rect 12618 21020 12624 21072
rect 12676 21020 12682 21072
rect 12802 21020 12808 21072
rect 12860 21060 12866 21072
rect 15473 21063 15531 21069
rect 12860 21032 14044 21060
rect 12860 21020 12866 21032
rect 3050 20992 3056 21004
rect 1872 20964 3056 20992
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20893 1639 20927
rect 1581 20887 1639 20893
rect 1596 20788 1624 20887
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 1872 20933 1900 20964
rect 3050 20952 3056 20964
rect 3108 20952 3114 21004
rect 3973 20995 4031 21001
rect 3973 20992 3985 20995
rect 3160 20964 3985 20992
rect 1857 20927 1915 20933
rect 1728 20896 1773 20924
rect 1728 20884 1734 20896
rect 1857 20893 1869 20927
rect 1903 20893 1915 20927
rect 1857 20887 1915 20893
rect 2038 20884 2044 20936
rect 2096 20933 2102 20936
rect 2096 20924 2104 20933
rect 2777 20927 2835 20933
rect 2096 20896 2141 20924
rect 2096 20887 2104 20896
rect 2777 20893 2789 20927
rect 2823 20893 2835 20927
rect 2777 20887 2835 20893
rect 2925 20927 2983 20933
rect 2925 20893 2937 20927
rect 2971 20924 2983 20927
rect 3160 20924 3188 20964
rect 3973 20961 3985 20964
rect 4019 20961 4031 20995
rect 5276 20992 5304 21020
rect 3973 20955 4031 20961
rect 4172 20964 5304 20992
rect 2971 20896 3188 20924
rect 2971 20893 2983 20896
rect 2925 20887 2983 20893
rect 2096 20884 2102 20887
rect 1949 20859 2007 20865
rect 1949 20825 1961 20859
rect 1995 20856 2007 20859
rect 2222 20856 2228 20868
rect 1995 20828 2228 20856
rect 1995 20825 2007 20828
rect 1949 20819 2007 20825
rect 2222 20816 2228 20828
rect 2280 20816 2286 20868
rect 2792 20856 2820 20887
rect 3234 20884 3240 20936
rect 3292 20933 3298 20936
rect 3292 20924 3300 20933
rect 3292 20896 3337 20924
rect 3292 20887 3300 20896
rect 3292 20884 3298 20887
rect 3510 20884 3516 20936
rect 3568 20924 3574 20936
rect 4172 20933 4200 20964
rect 6638 20952 6644 21004
rect 6696 20952 6702 21004
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 10137 20995 10195 21001
rect 10137 20992 10149 20995
rect 9364 20964 10149 20992
rect 9364 20952 9370 20964
rect 10137 20961 10149 20964
rect 10183 20961 10195 20995
rect 10137 20955 10195 20961
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 10778 20992 10784 21004
rect 10376 20964 10784 20992
rect 10376 20952 10382 20964
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 13906 20992 13912 21004
rect 11624 20964 13912 20992
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 3568 20896 4169 20924
rect 3568 20884 3574 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4157 20887 4215 20893
rect 4430 20884 4436 20936
rect 4488 20924 4494 20936
rect 5074 20924 5080 20936
rect 4488 20896 5080 20924
rect 4488 20884 4494 20896
rect 5074 20884 5080 20896
rect 5132 20884 5138 20936
rect 5258 20884 5264 20936
rect 5316 20884 5322 20936
rect 5442 20884 5448 20936
rect 5500 20924 5506 20936
rect 6122 20927 6180 20933
rect 6122 20924 6134 20927
rect 5500 20896 6134 20924
rect 5500 20884 5506 20896
rect 6122 20893 6134 20896
rect 6168 20893 6180 20927
rect 6122 20887 6180 20893
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20924 7987 20927
rect 8386 20924 8392 20936
rect 7975 20896 8392 20924
rect 7975 20893 7987 20896
rect 7929 20887 7987 20893
rect 3053 20859 3111 20865
rect 2792 20828 2912 20856
rect 2884 20800 2912 20828
rect 3053 20825 3065 20859
rect 3099 20825 3111 20859
rect 3053 20819 3111 20825
rect 3145 20859 3203 20865
rect 3145 20825 3157 20859
rect 3191 20856 3203 20859
rect 3694 20856 3700 20868
rect 3191 20828 3700 20856
rect 3191 20825 3203 20828
rect 3145 20819 3203 20825
rect 2314 20788 2320 20800
rect 1596 20760 2320 20788
rect 2314 20748 2320 20760
rect 2372 20788 2378 20800
rect 2866 20788 2872 20800
rect 2372 20760 2872 20788
rect 2372 20748 2378 20760
rect 2866 20748 2872 20760
rect 2924 20748 2930 20800
rect 3068 20788 3096 20819
rect 3694 20816 3700 20828
rect 3752 20816 3758 20868
rect 7300 20856 7328 20887
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 8570 20884 8576 20936
rect 8628 20884 8634 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 11624 20933 11652 20964
rect 13906 20952 13912 20964
rect 13964 20952 13970 21004
rect 14016 20992 14044 21032
rect 15473 21029 15485 21063
rect 15519 21060 15531 21063
rect 17770 21060 17776 21072
rect 15519 21032 17776 21060
rect 15519 21029 15531 21032
rect 15473 21023 15531 21029
rect 17770 21020 17776 21032
rect 17828 21020 17834 21072
rect 23106 21020 23112 21072
rect 23164 21020 23170 21072
rect 23216 21060 23244 21100
rect 23290 21088 23296 21140
rect 23348 21088 23354 21140
rect 27798 21128 27804 21140
rect 24504 21100 27804 21128
rect 23566 21060 23572 21072
rect 23216 21032 23572 21060
rect 23566 21020 23572 21032
rect 23624 21020 23630 21072
rect 19702 20992 19708 21004
rect 14016 20964 16344 20992
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 9732 20896 10977 20924
rect 9732 20884 9738 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20893 11667 20927
rect 11609 20887 11667 20893
rect 12345 20927 12403 20933
rect 12345 20893 12357 20927
rect 12391 20893 12403 20927
rect 12345 20887 12403 20893
rect 8294 20856 8300 20868
rect 7300 20828 8300 20856
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 8662 20816 8668 20868
rect 8720 20856 8726 20868
rect 9306 20856 9312 20868
rect 8720 20828 9312 20856
rect 8720 20816 8726 20828
rect 9306 20816 9312 20828
rect 9364 20856 9370 20868
rect 9953 20859 10011 20865
rect 9953 20856 9965 20859
rect 9364 20828 9965 20856
rect 9364 20816 9370 20828
rect 9953 20825 9965 20828
rect 9999 20825 10011 20859
rect 9953 20819 10011 20825
rect 11422 20816 11428 20868
rect 11480 20816 11486 20868
rect 12360 20856 12388 20887
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 13354 20924 13360 20936
rect 12492 20896 13360 20924
rect 12492 20884 12498 20896
rect 13354 20884 13360 20896
rect 13412 20924 13418 20936
rect 13412 20896 14612 20924
rect 13412 20884 13418 20896
rect 13170 20856 13176 20868
rect 12360 20828 13176 20856
rect 13170 20816 13176 20828
rect 13228 20816 13234 20868
rect 13265 20859 13323 20865
rect 13265 20825 13277 20859
rect 13311 20856 13323 20859
rect 13998 20856 14004 20868
rect 13311 20828 14004 20856
rect 13311 20825 13323 20828
rect 13265 20819 13323 20825
rect 4062 20788 4068 20800
rect 3068 20760 4068 20788
rect 4062 20748 4068 20760
rect 4120 20748 4126 20800
rect 4338 20748 4344 20800
rect 4396 20788 4402 20800
rect 6181 20791 6239 20797
rect 6181 20788 6193 20791
rect 4396 20760 6193 20788
rect 4396 20748 4402 20760
rect 6181 20757 6193 20760
rect 6227 20757 6239 20791
rect 6181 20751 6239 20757
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 9582 20788 9588 20800
rect 8435 20760 9588 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 10042 20748 10048 20800
rect 10100 20748 10106 20800
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 13280 20788 13308 20819
rect 13998 20816 14004 20828
rect 14056 20816 14062 20868
rect 14584 20865 14612 20896
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 16316 20933 16344 20964
rect 19444 20964 19708 20992
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 15804 20896 16129 20924
rect 15804 20884 15810 20896
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17862 20924 17868 20936
rect 17092 20896 17868 20924
rect 17092 20884 17098 20896
rect 17862 20884 17868 20896
rect 17920 20924 17926 20936
rect 19242 20924 19248 20936
rect 17920 20896 18644 20924
rect 17920 20884 17926 20896
rect 14369 20859 14427 20865
rect 14369 20825 14381 20859
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 14569 20859 14627 20865
rect 14569 20825 14581 20859
rect 14615 20825 14627 20859
rect 15102 20856 15108 20868
rect 14569 20819 14627 20825
rect 14660 20828 15108 20856
rect 10836 20760 13308 20788
rect 10836 20748 10842 20760
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14384 20788 14412 20819
rect 14660 20788 14688 20828
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 15289 20859 15347 20865
rect 15289 20825 15301 20859
rect 15335 20856 15347 20859
rect 15930 20856 15936 20868
rect 15335 20828 15936 20856
rect 15335 20825 15347 20828
rect 15289 20819 15347 20825
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 17405 20859 17463 20865
rect 17405 20856 17417 20859
rect 16080 20828 17417 20856
rect 16080 20816 16086 20828
rect 17405 20825 17417 20828
rect 17451 20856 17463 20859
rect 17494 20856 17500 20868
rect 17451 20828 17500 20856
rect 17451 20825 17463 20828
rect 17405 20819 17463 20825
rect 17494 20816 17500 20828
rect 17552 20816 17558 20868
rect 17678 20865 17684 20868
rect 17621 20859 17684 20865
rect 17621 20825 17633 20859
rect 17667 20825 17684 20859
rect 17621 20819 17684 20825
rect 17678 20816 17684 20819
rect 17736 20856 17742 20868
rect 18322 20856 18328 20868
rect 17736 20828 18328 20856
rect 17736 20816 17742 20828
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20825 18567 20859
rect 18616 20856 18644 20896
rect 18800 20896 19248 20924
rect 18709 20859 18767 20865
rect 18709 20856 18721 20859
rect 18616 20828 18721 20856
rect 18509 20819 18567 20825
rect 18709 20825 18721 20828
rect 18755 20825 18767 20859
rect 18709 20819 18767 20825
rect 13964 20760 14688 20788
rect 14737 20791 14795 20797
rect 13964 20748 13970 20760
rect 14737 20757 14749 20791
rect 14783 20788 14795 20791
rect 16298 20788 16304 20800
rect 14783 20760 16304 20788
rect 14783 20757 14795 20760
rect 14737 20751 14795 20757
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 17770 20748 17776 20800
rect 17828 20748 17834 20800
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 18524 20788 18552 20819
rect 18800 20788 18828 20896
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 19444 20933 19472 20964
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 24394 20992 24400 21004
rect 20947 20964 24400 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 24394 20952 24400 20964
rect 24452 20952 24458 21004
rect 19610 20933 19616 20936
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19577 20927 19616 20933
rect 19577 20893 19589 20927
rect 19577 20887 19616 20893
rect 19610 20884 19616 20887
rect 19668 20884 19674 20936
rect 19794 20884 19800 20936
rect 19852 20884 19858 20936
rect 19886 20884 19892 20936
rect 19944 20933 19950 20936
rect 19944 20924 19952 20933
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 19944 20896 19989 20924
rect 20548 20896 21373 20924
rect 19944 20887 19952 20896
rect 19944 20884 19950 20887
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 19705 20859 19763 20865
rect 19705 20856 19717 20859
rect 19208 20828 19717 20856
rect 19208 20816 19214 20828
rect 19705 20825 19717 20828
rect 19751 20825 19763 20859
rect 19705 20819 19763 20825
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 20548 20865 20576 20896
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 20533 20859 20591 20865
rect 20533 20856 20545 20859
rect 20496 20828 20545 20856
rect 20496 20816 20502 20828
rect 20533 20825 20545 20828
rect 20579 20825 20591 20859
rect 20533 20819 20591 20825
rect 20717 20859 20775 20865
rect 20717 20825 20729 20859
rect 20763 20856 20775 20859
rect 20806 20856 20812 20868
rect 20763 20828 20812 20856
rect 20763 20825 20775 20828
rect 20717 20819 20775 20825
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 21542 20816 21548 20868
rect 21600 20816 21606 20868
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 22833 20859 22891 20865
rect 22833 20856 22845 20859
rect 22152 20828 22845 20856
rect 22152 20816 22158 20828
rect 22833 20825 22845 20828
rect 22879 20856 22891 20859
rect 23014 20856 23020 20868
rect 22879 20828 23020 20856
rect 22879 20825 22891 20828
rect 22833 20819 22891 20825
rect 23014 20816 23020 20828
rect 23072 20816 23078 20868
rect 18012 20760 18828 20788
rect 18877 20791 18935 20797
rect 18012 20748 18018 20760
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 19610 20788 19616 20800
rect 18923 20760 19616 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 20070 20748 20076 20800
rect 20128 20748 20134 20800
rect 20824 20788 20852 20816
rect 24504 20788 24532 21100
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 24578 20952 24584 21004
rect 24636 20952 24642 21004
rect 24848 20927 24906 20933
rect 24848 20893 24860 20927
rect 24894 20924 24906 20927
rect 25130 20924 25136 20936
rect 24894 20896 25136 20924
rect 24894 20893 24906 20896
rect 24848 20887 24906 20893
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 24946 20816 24952 20868
rect 25004 20856 25010 20868
rect 27034 20859 27092 20865
rect 27034 20856 27046 20859
rect 25004 20828 27046 20856
rect 25004 20816 25010 20828
rect 27034 20825 27046 20828
rect 27080 20825 27092 20859
rect 27034 20819 27092 20825
rect 20824 20760 24532 20788
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25924 20760 25973 20788
rect 25924 20748 25930 20760
rect 25961 20757 25973 20760
rect 26007 20757 26019 20791
rect 25961 20751 26019 20757
rect 26326 20748 26332 20800
rect 26384 20788 26390 20800
rect 28169 20791 28227 20797
rect 28169 20788 28181 20791
rect 26384 20760 28181 20788
rect 26384 20748 26390 20760
rect 28169 20757 28181 20760
rect 28215 20757 28227 20791
rect 28169 20751 28227 20757
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 1302 20544 1308 20596
rect 1360 20584 1366 20596
rect 2406 20584 2412 20596
rect 1360 20556 2412 20584
rect 1360 20544 1366 20556
rect 2406 20544 2412 20556
rect 2464 20544 2470 20596
rect 3510 20584 3516 20596
rect 3068 20556 3516 20584
rect 2866 20516 2872 20528
rect 1596 20488 2872 20516
rect 1596 20457 1624 20488
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20417 1639 20451
rect 1581 20411 1639 20417
rect 1670 20408 1676 20460
rect 1728 20448 1734 20460
rect 1765 20451 1823 20457
rect 1765 20448 1777 20451
rect 1728 20420 1777 20448
rect 1728 20408 1734 20420
rect 1765 20417 1777 20420
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 2130 20408 2136 20460
rect 2188 20448 2194 20460
rect 3068 20457 3096 20556
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 3620 20556 4936 20584
rect 3620 20516 3648 20556
rect 3160 20488 3648 20516
rect 2317 20451 2375 20457
rect 2317 20448 2329 20451
rect 2188 20420 2329 20448
rect 2188 20408 2194 20420
rect 2317 20417 2329 20420
rect 2363 20417 2375 20451
rect 2317 20411 2375 20417
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 1118 20340 1124 20392
rect 1176 20380 1182 20392
rect 3160 20380 3188 20488
rect 3234 20408 3240 20460
rect 3292 20408 3298 20460
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20448 3387 20451
rect 3510 20448 3516 20460
rect 3375 20420 3516 20448
rect 3375 20417 3387 20420
rect 3329 20411 3387 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 3620 20457 3648 20488
rect 4246 20476 4252 20528
rect 4304 20516 4310 20528
rect 4617 20519 4675 20525
rect 4617 20516 4629 20519
rect 4304 20488 4629 20516
rect 4304 20476 4310 20488
rect 4617 20485 4629 20488
rect 4663 20485 4675 20519
rect 4617 20479 4675 20485
rect 4706 20476 4712 20528
rect 4764 20476 4770 20528
rect 4908 20516 4936 20556
rect 4982 20544 4988 20596
rect 5040 20544 5046 20596
rect 5074 20544 5080 20596
rect 5132 20584 5138 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 5132 20556 5825 20584
rect 5132 20544 5138 20556
rect 5813 20553 5825 20556
rect 5859 20584 5871 20587
rect 8665 20587 8723 20593
rect 8665 20584 8677 20587
rect 5859 20556 8677 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 8665 20553 8677 20556
rect 8711 20584 8723 20587
rect 12529 20587 12587 20593
rect 8711 20556 12434 20584
rect 8711 20553 8723 20556
rect 8665 20547 8723 20553
rect 5629 20519 5687 20525
rect 5629 20516 5641 20519
rect 4908 20488 5641 20516
rect 5629 20485 5641 20488
rect 5675 20516 5687 20519
rect 5902 20516 5908 20528
rect 5675 20488 5908 20516
rect 5675 20485 5687 20488
rect 5629 20479 5687 20485
rect 5902 20476 5908 20488
rect 5960 20516 5966 20528
rect 5960 20488 6224 20516
rect 5960 20476 5966 20488
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 4430 20408 4436 20460
rect 4488 20408 4494 20460
rect 4982 20458 4988 20460
rect 4816 20457 4988 20458
rect 4801 20451 4988 20457
rect 4801 20417 4813 20451
rect 4847 20430 4988 20451
rect 4847 20417 4859 20430
rect 4801 20411 4859 20417
rect 4982 20408 4988 20430
rect 5040 20408 5046 20460
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 6196 20448 6224 20488
rect 6730 20476 6736 20528
rect 6788 20516 6794 20528
rect 7653 20519 7711 20525
rect 7653 20516 7665 20519
rect 6788 20488 7665 20516
rect 6788 20476 6794 20488
rect 7653 20485 7665 20488
rect 7699 20485 7711 20519
rect 10226 20516 10232 20528
rect 7653 20479 7711 20485
rect 9646 20488 10232 20516
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 6196 20420 6929 20448
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20448 7159 20451
rect 7374 20448 7380 20460
rect 7147 20420 7380 20448
rect 7147 20417 7159 20420
rect 7101 20411 7159 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 9646 20448 9674 20488
rect 10226 20476 10232 20488
rect 10284 20516 10290 20528
rect 11793 20519 11851 20525
rect 10284 20488 10364 20516
rect 10284 20476 10290 20488
rect 7616 20420 9674 20448
rect 7616 20408 7622 20420
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 9916 20420 10057 20448
rect 9916 20408 9922 20420
rect 1176 20352 3188 20380
rect 3421 20383 3479 20389
rect 1176 20340 1182 20352
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 4154 20380 4160 20392
rect 3467 20352 4160 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 5442 20340 5448 20392
rect 5500 20340 5506 20392
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 5552 20352 8769 20380
rect 1581 20315 1639 20321
rect 1581 20281 1593 20315
rect 1627 20312 1639 20315
rect 1627 20284 2636 20312
rect 1627 20281 1639 20284
rect 1581 20275 1639 20281
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 2501 20247 2559 20253
rect 2501 20244 2513 20247
rect 1544 20216 2513 20244
rect 1544 20204 1550 20216
rect 2501 20213 2513 20216
rect 2547 20213 2559 20247
rect 2608 20244 2636 20284
rect 4798 20272 4804 20324
rect 4856 20312 4862 20324
rect 5552 20312 5580 20352
rect 8757 20349 8769 20352
rect 8803 20349 8815 20383
rect 8757 20343 8815 20349
rect 8846 20340 8852 20392
rect 8904 20340 8910 20392
rect 4856 20284 5580 20312
rect 4856 20272 4862 20284
rect 6086 20272 6092 20324
rect 6144 20312 6150 20324
rect 7009 20315 7067 20321
rect 7009 20312 7021 20315
rect 6144 20284 7021 20312
rect 6144 20272 6150 20284
rect 7009 20281 7021 20284
rect 7055 20312 7067 20315
rect 9766 20312 9772 20324
rect 7055 20284 9772 20312
rect 7055 20281 7067 20284
rect 7009 20275 7067 20281
rect 9766 20272 9772 20284
rect 9824 20272 9830 20324
rect 9968 20312 9996 20420
rect 10045 20417 10057 20420
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10134 20408 10140 20460
rect 10192 20408 10198 20460
rect 10336 20457 10364 20488
rect 11793 20485 11805 20519
rect 11839 20516 11851 20519
rect 11882 20516 11888 20528
rect 11839 20488 11888 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 11146 20448 11152 20460
rect 10367 20420 11152 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 12406 20448 12434 20556
rect 12529 20553 12541 20587
rect 12575 20584 12587 20587
rect 13538 20584 13544 20596
rect 12575 20556 13544 20584
rect 12575 20553 12587 20556
rect 12529 20547 12587 20553
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 14369 20587 14427 20593
rect 14369 20553 14381 20587
rect 14415 20584 14427 20587
rect 14458 20584 14464 20596
rect 14415 20556 14464 20584
rect 14415 20553 14427 20556
rect 14369 20547 14427 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 17221 20587 17279 20593
rect 17221 20553 17233 20587
rect 17267 20584 17279 20587
rect 18230 20584 18236 20596
rect 17267 20556 18236 20584
rect 17267 20553 17279 20556
rect 17221 20547 17279 20553
rect 18230 20544 18236 20556
rect 18288 20544 18294 20596
rect 20070 20584 20076 20596
rect 18340 20556 20076 20584
rect 13446 20476 13452 20528
rect 13504 20516 13510 20528
rect 15289 20519 15347 20525
rect 15289 20516 15301 20519
rect 13504 20488 15301 20516
rect 13504 20476 13510 20488
rect 15289 20485 15301 20488
rect 15335 20485 15347 20519
rect 18340 20516 18368 20556
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 21269 20587 21327 20593
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 24210 20584 24216 20596
rect 21315 20556 24216 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 24210 20544 24216 20556
rect 24268 20544 24274 20596
rect 25682 20544 25688 20596
rect 25740 20584 25746 20596
rect 26605 20587 26663 20593
rect 26605 20584 26617 20587
rect 25740 20556 26617 20584
rect 25740 20544 25746 20556
rect 26605 20553 26617 20556
rect 26651 20553 26663 20587
rect 26605 20547 26663 20553
rect 21542 20516 21548 20528
rect 15289 20479 15347 20485
rect 15488 20488 18368 20516
rect 19076 20488 21548 20516
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 12406 20420 13185 20448
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13320 20420 14197 20448
rect 13320 20408 13326 20420
rect 14185 20417 14197 20420
rect 14231 20448 14243 20451
rect 14826 20448 14832 20460
rect 14231 20420 14832 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 15488 20457 15516 20488
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 16482 20448 16488 20460
rect 15611 20420 16488 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20448 17095 20451
rect 17494 20448 17500 20460
rect 17083 20420 17500 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 17862 20408 17868 20460
rect 17920 20408 17926 20460
rect 18874 20408 18880 20460
rect 18932 20408 18938 20460
rect 19076 20457 19104 20488
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 21726 20476 21732 20528
rect 21784 20516 21790 20528
rect 24762 20516 24768 20528
rect 21784 20488 24768 20516
rect 21784 20476 21790 20488
rect 24762 20476 24768 20488
rect 24820 20476 24826 20528
rect 19025 20451 19104 20457
rect 19025 20417 19037 20451
rect 19071 20420 19104 20451
rect 19071 20417 19083 20420
rect 19025 20411 19083 20417
rect 19150 20408 19156 20460
rect 19208 20408 19214 20460
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19342 20451 19400 20457
rect 19342 20417 19354 20451
rect 19388 20448 19400 20451
rect 19886 20448 19892 20460
rect 19388 20420 19892 20448
rect 19388 20417 19400 20420
rect 19342 20411 19400 20417
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 11112 20352 12265 20380
rect 11112 20340 11118 20352
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 12434 20380 12440 20392
rect 12391 20352 12440 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 13078 20340 13084 20392
rect 13136 20340 13142 20392
rect 13998 20340 14004 20392
rect 14056 20380 14062 20392
rect 15286 20380 15292 20392
rect 14056 20352 15292 20380
rect 14056 20340 14062 20352
rect 15286 20340 15292 20352
rect 15344 20380 15350 20392
rect 15746 20380 15752 20392
rect 15344 20352 15752 20380
rect 15344 20340 15350 20352
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 16868 20380 16896 20408
rect 17586 20380 17592 20392
rect 16868 20352 17592 20380
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 17681 20383 17739 20389
rect 17681 20349 17693 20383
rect 17727 20380 17739 20383
rect 17954 20380 17960 20392
rect 17727 20352 17960 20380
rect 17727 20349 17739 20352
rect 17681 20343 17739 20349
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 19352 20380 19380 20411
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 20438 20408 20444 20460
rect 20496 20408 20502 20460
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 21453 20451 21511 20457
rect 21453 20448 21465 20451
rect 20855 20420 21465 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 21453 20417 21465 20420
rect 21499 20417 21511 20451
rect 22445 20451 22503 20457
rect 22445 20448 22457 20451
rect 21453 20411 21511 20417
rect 22066 20420 22457 20448
rect 18095 20352 19380 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 19518 20340 19524 20392
rect 19576 20380 19582 20392
rect 19794 20380 19800 20392
rect 19576 20352 19800 20380
rect 19576 20340 19582 20352
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 22066 20380 22094 20420
rect 22445 20417 22457 20420
rect 22491 20417 22503 20451
rect 22445 20411 22503 20417
rect 22738 20408 22744 20460
rect 22796 20448 22802 20460
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 22796 20420 24225 20448
rect 22796 20408 22802 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 25130 20448 25136 20460
rect 24636 20420 25136 20448
rect 24636 20408 24642 20420
rect 25130 20408 25136 20420
rect 25188 20448 25194 20460
rect 25225 20451 25283 20457
rect 25225 20448 25237 20451
rect 25188 20420 25237 20448
rect 25188 20408 25194 20420
rect 25225 20417 25237 20420
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 25492 20451 25550 20457
rect 25492 20417 25504 20451
rect 25538 20448 25550 20451
rect 26234 20448 26240 20460
rect 25538 20420 26240 20448
rect 25538 20417 25550 20420
rect 25492 20411 25550 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 20036 20352 22094 20380
rect 22189 20383 22247 20389
rect 20036 20340 20042 20352
rect 22189 20349 22201 20383
rect 22235 20349 22247 20383
rect 22189 20343 22247 20349
rect 10686 20312 10692 20324
rect 9968 20284 10692 20312
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 10778 20272 10784 20324
rect 10836 20312 10842 20324
rect 11793 20315 11851 20321
rect 11793 20312 11805 20315
rect 10836 20284 11805 20312
rect 10836 20272 10842 20284
rect 11793 20281 11805 20284
rect 11839 20281 11851 20315
rect 19886 20312 19892 20324
rect 11793 20275 11851 20281
rect 19444 20284 19892 20312
rect 3142 20244 3148 20256
rect 2608 20216 3148 20244
rect 2501 20207 2559 20213
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 3786 20204 3792 20256
rect 3844 20204 3850 20256
rect 4706 20204 4712 20256
rect 4764 20244 4770 20256
rect 5534 20244 5540 20256
rect 4764 20216 5540 20244
rect 4764 20204 4770 20216
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6270 20244 6276 20256
rect 6043 20216 6276 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7745 20247 7803 20253
rect 7745 20244 7757 20247
rect 7432 20216 7757 20244
rect 7432 20204 7438 20216
rect 7745 20213 7757 20216
rect 7791 20213 7803 20247
rect 7745 20207 7803 20213
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 8297 20247 8355 20253
rect 8297 20244 8309 20247
rect 7892 20216 8309 20244
rect 7892 20204 7898 20216
rect 8297 20213 8309 20216
rect 8343 20213 8355 20247
rect 8297 20207 8355 20213
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 8904 20216 10149 20244
rect 8904 20204 8910 20216
rect 10137 20213 10149 20216
rect 10183 20213 10195 20247
rect 10137 20207 10195 20213
rect 10226 20204 10232 20256
rect 10284 20244 10290 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 10284 20216 13461 20244
rect 10284 20204 10290 20216
rect 13449 20213 13461 20216
rect 13495 20213 13507 20247
rect 13449 20207 13507 20213
rect 13998 20204 14004 20256
rect 14056 20244 14062 20256
rect 14182 20244 14188 20256
rect 14056 20216 14188 20244
rect 14056 20204 14062 20216
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 15562 20204 15568 20256
rect 15620 20204 15626 20256
rect 15746 20204 15752 20256
rect 15804 20204 15810 20256
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 19444 20244 19472 20284
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 20622 20272 20628 20324
rect 20680 20312 20686 20324
rect 21726 20312 21732 20324
rect 20680 20284 21732 20312
rect 20680 20272 20686 20284
rect 21726 20272 21732 20284
rect 21784 20272 21790 20324
rect 16080 20216 19472 20244
rect 16080 20204 16086 20216
rect 19518 20204 19524 20256
rect 19576 20204 19582 20256
rect 22204 20244 22232 20343
rect 22830 20244 22836 20256
rect 22204 20216 22836 20244
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 23566 20204 23572 20256
rect 23624 20204 23630 20256
rect 24029 20247 24087 20253
rect 24029 20213 24041 20247
rect 24075 20244 24087 20247
rect 26510 20244 26516 20256
rect 24075 20216 26516 20244
rect 24075 20213 24087 20216
rect 24029 20207 24087 20213
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 2409 20043 2467 20049
rect 2409 20009 2421 20043
rect 2455 20040 2467 20043
rect 3970 20040 3976 20052
rect 2455 20012 3976 20040
rect 2455 20009 2467 20012
rect 2409 20003 2467 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4890 20040 4896 20052
rect 4387 20012 4896 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 4985 20043 5043 20049
rect 4985 20009 4997 20043
rect 5031 20040 5043 20043
rect 7834 20040 7840 20052
rect 5031 20012 7840 20040
rect 5031 20009 5043 20012
rect 4985 20003 5043 20009
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8294 20000 8300 20052
rect 8352 20000 8358 20052
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 9493 20043 9551 20049
rect 9493 20040 9505 20043
rect 8444 20012 9505 20040
rect 8444 20000 8450 20012
rect 9493 20009 9505 20012
rect 9539 20009 9551 20043
rect 11698 20040 11704 20052
rect 9493 20003 9551 20009
rect 9968 20012 11704 20040
rect 2590 19932 2596 19984
rect 2648 19972 2654 19984
rect 5077 19975 5135 19981
rect 5077 19972 5089 19975
rect 2648 19944 5089 19972
rect 2648 19932 2654 19944
rect 5077 19941 5089 19944
rect 5123 19941 5135 19975
rect 5077 19935 5135 19941
rect 5442 19932 5448 19984
rect 5500 19972 5506 19984
rect 8205 19975 8263 19981
rect 5500 19944 6224 19972
rect 5500 19932 5506 19944
rect 5166 19864 5172 19916
rect 5224 19864 5230 19916
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 5684 19876 6040 19904
rect 5684 19864 5690 19876
rect 2585 19849 2643 19855
rect 1946 19796 1952 19848
rect 2004 19796 2010 19848
rect 2585 19846 2597 19849
rect 2424 19818 2597 19846
rect 1854 19728 1860 19780
rect 1912 19768 1918 19780
rect 2424 19768 2452 19818
rect 2585 19815 2597 19818
rect 2631 19815 2643 19849
rect 2585 19809 2643 19815
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19805 2743 19839
rect 2685 19799 2743 19805
rect 2700 19768 2728 19799
rect 2866 19796 2872 19848
rect 2924 19796 2930 19848
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3326 19836 3332 19848
rect 3007 19808 3332 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 3602 19796 3608 19848
rect 3660 19836 3666 19848
rect 3970 19836 3976 19848
rect 3660 19808 3976 19836
rect 3660 19796 3666 19808
rect 3970 19796 3976 19808
rect 4028 19836 4034 19848
rect 4065 19839 4123 19845
rect 4065 19836 4077 19839
rect 4028 19808 4077 19836
rect 4028 19796 4034 19808
rect 4065 19805 4077 19808
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4706 19836 4712 19848
rect 4212 19808 4712 19836
rect 4212 19796 4218 19808
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19836 5871 19839
rect 5902 19836 5908 19848
rect 5859 19808 5908 19836
rect 5859 19805 5871 19808
rect 5813 19799 5871 19805
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 6012 19845 6040 19876
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 6196 19836 6224 19944
rect 8205 19941 8217 19975
rect 8251 19972 8263 19975
rect 9968 19972 9996 20012
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12069 20043 12127 20049
rect 12069 20040 12081 20043
rect 12032 20012 12081 20040
rect 12032 20000 12038 20012
rect 12069 20009 12081 20012
rect 12115 20009 12127 20043
rect 12069 20003 12127 20009
rect 12253 20043 12311 20049
rect 12253 20009 12265 20043
rect 12299 20040 12311 20043
rect 12526 20040 12532 20052
rect 12299 20012 12532 20040
rect 12299 20009 12311 20012
rect 12253 20003 12311 20009
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 12989 20043 13047 20049
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13078 20040 13084 20052
rect 13035 20012 13084 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13630 20000 13636 20052
rect 13688 20000 13694 20052
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 8251 19944 9996 19972
rect 8251 19941 8263 19944
rect 8205 19935 8263 19941
rect 12618 19932 12624 19984
rect 12676 19972 12682 19984
rect 12894 19972 12900 19984
rect 12676 19944 12900 19972
rect 12676 19932 12682 19944
rect 12894 19932 12900 19944
rect 12952 19932 12958 19984
rect 14936 19972 14964 20003
rect 15470 20000 15476 20052
rect 15528 20040 15534 20052
rect 15565 20043 15623 20049
rect 15565 20040 15577 20043
rect 15528 20012 15577 20040
rect 15528 20000 15534 20012
rect 15565 20009 15577 20012
rect 15611 20009 15623 20043
rect 15565 20003 15623 20009
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16206 20040 16212 20052
rect 16071 20012 16212 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 17770 20040 17776 20052
rect 17359 20012 17776 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 17920 20012 18337 20040
rect 17920 20000 17926 20012
rect 18325 20009 18337 20012
rect 18371 20040 18383 20043
rect 18966 20040 18972 20052
rect 18371 20012 18972 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 18966 20000 18972 20012
rect 19024 20040 19030 20052
rect 19889 20043 19947 20049
rect 19024 20012 19840 20040
rect 19024 20000 19030 20012
rect 16666 19972 16672 19984
rect 14936 19944 16672 19972
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 17405 19975 17463 19981
rect 17405 19941 17417 19975
rect 17451 19972 17463 19975
rect 18046 19972 18052 19984
rect 17451 19944 18052 19972
rect 17451 19941 17463 19944
rect 17405 19935 17463 19941
rect 18046 19932 18052 19944
rect 18104 19932 18110 19984
rect 19426 19932 19432 19984
rect 19484 19972 19490 19984
rect 19705 19975 19763 19981
rect 19705 19972 19717 19975
rect 19484 19944 19717 19972
rect 19484 19932 19490 19944
rect 19705 19941 19717 19944
rect 19751 19941 19763 19975
rect 19812 19972 19840 20012
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20714 20040 20720 20052
rect 19935 20012 20720 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 21177 20043 21235 20049
rect 21177 20009 21189 20043
rect 21223 20040 21235 20043
rect 21266 20040 21272 20052
rect 21223 20012 21272 20040
rect 21223 20009 21235 20012
rect 21177 20003 21235 20009
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 22925 20043 22983 20049
rect 22925 20009 22937 20043
rect 22971 20040 22983 20043
rect 24946 20040 24952 20052
rect 22971 20012 24952 20040
rect 22971 20009 22983 20012
rect 22925 20003 22983 20009
rect 24946 20000 24952 20012
rect 25004 20000 25010 20052
rect 22186 19972 22192 19984
rect 19812 19944 22192 19972
rect 19705 19935 19763 19941
rect 22186 19932 22192 19944
rect 22244 19932 22250 19984
rect 22281 19975 22339 19981
rect 22281 19941 22293 19975
rect 22327 19972 22339 19975
rect 26418 19972 26424 19984
rect 22327 19944 26424 19972
rect 22327 19941 22339 19944
rect 22281 19935 22339 19941
rect 26418 19932 26424 19944
rect 26476 19932 26482 19984
rect 6730 19864 6736 19916
rect 6788 19864 6794 19916
rect 9950 19864 9956 19916
rect 10008 19864 10014 19916
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 11882 19904 11888 19916
rect 11388 19876 11888 19904
rect 11388 19864 11394 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 15749 19907 15807 19913
rect 12400 19876 13584 19904
rect 12400 19864 12406 19876
rect 6917 19839 6975 19845
rect 6917 19836 6929 19839
rect 6196 19808 6929 19836
rect 6917 19805 6929 19808
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7098 19796 7104 19848
rect 7156 19796 7162 19848
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9214 19836 9220 19848
rect 9171 19808 9220 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 1912 19740 2452 19768
rect 2611 19740 2728 19768
rect 1912 19728 1918 19740
rect 842 19660 848 19712
rect 900 19700 906 19712
rect 1765 19703 1823 19709
rect 1765 19700 1777 19703
rect 900 19672 1777 19700
rect 900 19660 906 19672
rect 1765 19669 1777 19672
rect 1811 19669 1823 19703
rect 1765 19663 1823 19669
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 2611 19700 2639 19740
rect 2774 19728 2780 19780
rect 2832 19768 2838 19780
rect 4798 19768 4804 19780
rect 2832 19740 4804 19768
rect 2832 19728 2838 19740
rect 4798 19728 4804 19740
rect 4856 19728 4862 19780
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 7208 19768 7236 19799
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 12526 19836 12532 19848
rect 10152 19808 12532 19836
rect 6236 19740 7236 19768
rect 7837 19771 7895 19777
rect 6236 19728 6242 19740
rect 7837 19737 7849 19771
rect 7883 19768 7895 19771
rect 8662 19768 8668 19780
rect 7883 19740 8668 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 8662 19728 8668 19740
rect 8720 19728 8726 19780
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 10152 19768 10180 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12676 19808 12817 19836
rect 12676 19796 12682 19808
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13446 19836 13452 19848
rect 13228 19808 13452 19836
rect 13228 19796 13234 19808
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 13556 19845 13584 19876
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 19518 19904 19524 19916
rect 15795 19876 19524 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 21082 19864 21088 19916
rect 21140 19904 21146 19916
rect 23566 19904 23572 19916
rect 21140 19876 23572 19904
rect 21140 19864 21146 19876
rect 23566 19864 23572 19876
rect 23624 19864 23630 19916
rect 26786 19864 26792 19916
rect 26844 19904 26850 19916
rect 26973 19907 27031 19913
rect 26973 19904 26985 19907
rect 26844 19876 26985 19904
rect 26844 19864 26850 19876
rect 26973 19873 26985 19876
rect 27019 19873 27031 19907
rect 26973 19867 27031 19873
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 14366 19796 14372 19848
rect 14424 19836 14430 19848
rect 14918 19836 14924 19848
rect 14424 19808 14924 19836
rect 14424 19796 14430 19808
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15436 19808 15577 19836
rect 15436 19796 15442 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 15838 19796 15844 19848
rect 15896 19796 15902 19848
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16298 19836 16304 19848
rect 15988 19808 16304 19836
rect 15988 19796 15994 19808
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17402 19836 17408 19848
rect 17267 19808 17408 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17494 19796 17500 19848
rect 17552 19796 17558 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 17681 19799 17739 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19836 19487 19839
rect 19794 19836 19800 19848
rect 19475 19808 19800 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 9355 19740 10180 19768
rect 10220 19771 10278 19777
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 10220 19737 10232 19771
rect 10266 19737 10278 19771
rect 10220 19731 10278 19737
rect 2280 19672 2639 19700
rect 2280 19660 2286 19672
rect 5626 19660 5632 19712
rect 5684 19660 5690 19712
rect 9490 19660 9496 19712
rect 9548 19700 9554 19712
rect 10244 19700 10272 19731
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 11296 19740 11897 19768
rect 11296 19728 11302 19740
rect 11885 19737 11897 19740
rect 11931 19768 11943 19771
rect 14274 19768 14280 19780
rect 11931 19740 14280 19768
rect 11931 19737 11943 19740
rect 11885 19731 11943 19737
rect 14274 19728 14280 19740
rect 14332 19728 14338 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 14384 19740 14749 19768
rect 9548 19672 10272 19700
rect 11333 19703 11391 19709
rect 9548 19660 9554 19672
rect 11333 19669 11345 19703
rect 11379 19700 11391 19703
rect 11790 19700 11796 19712
rect 11379 19672 11796 19700
rect 11379 19669 11391 19672
rect 11333 19663 11391 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 12066 19660 12072 19712
rect 12124 19709 12130 19712
rect 12124 19703 12143 19709
rect 12131 19669 12143 19703
rect 12124 19663 12143 19669
rect 12124 19660 12130 19663
rect 12986 19660 12992 19712
rect 13044 19700 13050 19712
rect 14384 19700 14412 19740
rect 14737 19737 14749 19740
rect 14783 19737 14795 19771
rect 15654 19768 15660 19780
rect 14737 19731 14795 19737
rect 14844 19740 15660 19768
rect 13044 19672 14412 19700
rect 13044 19660 13050 19672
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 14844 19700 14872 19740
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16945 19771 17003 19777
rect 16945 19768 16957 19771
rect 15804 19740 16957 19768
rect 15804 19728 15810 19740
rect 16945 19737 16957 19740
rect 16991 19737 17003 19771
rect 16945 19731 17003 19737
rect 17310 19728 17316 19780
rect 17368 19768 17374 19780
rect 17696 19768 17724 19799
rect 17368 19740 17724 19768
rect 17368 19728 17374 19740
rect 14516 19672 14872 19700
rect 14516 19660 14522 19672
rect 14918 19660 14924 19712
rect 14976 19709 14982 19712
rect 14976 19703 14995 19709
rect 14983 19669 14995 19703
rect 14976 19663 14995 19669
rect 14976 19660 14982 19663
rect 15102 19660 15108 19712
rect 15160 19660 15166 19712
rect 15672 19700 15700 19728
rect 18156 19700 18184 19799
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 20772 19808 21833 19836
rect 20772 19796 20778 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 22465 19839 22523 19845
rect 22465 19836 22477 19839
rect 22336 19808 22477 19836
rect 22336 19796 22342 19808
rect 22465 19805 22477 19808
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 19518 19728 19524 19780
rect 19576 19768 19582 19780
rect 20438 19768 20444 19780
rect 19576 19740 20444 19768
rect 19576 19728 19582 19740
rect 20438 19728 20444 19740
rect 20496 19768 20502 19780
rect 20809 19771 20867 19777
rect 20809 19768 20821 19771
rect 20496 19740 20821 19768
rect 20496 19728 20502 19740
rect 20809 19737 20821 19740
rect 20855 19737 20867 19771
rect 20809 19731 20867 19737
rect 20993 19771 21051 19777
rect 20993 19737 21005 19771
rect 21039 19737 21051 19771
rect 20993 19731 21051 19737
rect 15672 19672 18184 19700
rect 21008 19700 21036 19731
rect 21174 19728 21180 19780
rect 21232 19768 21238 19780
rect 23124 19768 23152 19799
rect 24026 19796 24032 19848
rect 24084 19796 24090 19848
rect 21232 19740 23152 19768
rect 21232 19728 21238 19740
rect 24210 19728 24216 19780
rect 24268 19768 24274 19780
rect 27218 19771 27276 19777
rect 27218 19768 27230 19771
rect 24268 19740 27230 19768
rect 24268 19728 24274 19740
rect 27218 19737 27230 19740
rect 27264 19737 27276 19771
rect 27218 19731 27276 19737
rect 21542 19700 21548 19712
rect 21008 19672 21548 19700
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 21637 19703 21695 19709
rect 21637 19669 21649 19703
rect 21683 19700 21695 19703
rect 22554 19700 22560 19712
rect 21683 19672 22560 19700
rect 21683 19669 21695 19672
rect 21637 19663 21695 19669
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 23845 19703 23903 19709
rect 23845 19669 23857 19703
rect 23891 19700 23903 19703
rect 26050 19700 26056 19712
rect 23891 19672 26056 19700
rect 23891 19669 23903 19672
rect 23845 19663 23903 19669
rect 26050 19660 26056 19672
rect 26108 19660 26114 19712
rect 28350 19660 28356 19712
rect 28408 19660 28414 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 2498 19496 2504 19508
rect 2148 19468 2504 19496
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 2041 19363 2099 19369
rect 2041 19329 2053 19363
rect 2087 19360 2099 19363
rect 2148 19360 2176 19468
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 2774 19456 2780 19508
rect 2832 19456 2838 19508
rect 2961 19499 3019 19505
rect 2961 19465 2973 19499
rect 3007 19496 3019 19499
rect 3142 19496 3148 19508
rect 3007 19468 3148 19496
rect 3007 19465 3019 19468
rect 2961 19459 3019 19465
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 4163 19499 4221 19505
rect 4163 19496 4175 19499
rect 3292 19468 4175 19496
rect 3292 19456 3298 19468
rect 4163 19465 4175 19468
rect 4209 19465 4221 19499
rect 4163 19459 4221 19465
rect 4249 19499 4307 19505
rect 4249 19465 4261 19499
rect 4295 19496 4307 19499
rect 4430 19496 4436 19508
rect 4295 19468 4436 19496
rect 4295 19465 4307 19468
rect 4249 19459 4307 19465
rect 4430 19456 4436 19468
rect 4488 19496 4494 19508
rect 4798 19496 4804 19508
rect 4488 19468 4804 19496
rect 4488 19456 4494 19468
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 9039 19499 9097 19505
rect 9039 19496 9051 19499
rect 5224 19468 9051 19496
rect 5224 19456 5230 19468
rect 9039 19465 9051 19468
rect 9085 19465 9097 19499
rect 9039 19459 9097 19465
rect 9950 19456 9956 19508
rect 10008 19456 10014 19508
rect 10778 19456 10784 19508
rect 10836 19496 10842 19508
rect 11238 19496 11244 19508
rect 10836 19468 11244 19496
rect 10836 19456 10842 19468
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 12529 19499 12587 19505
rect 12529 19465 12541 19499
rect 12575 19496 12587 19499
rect 14458 19496 14464 19508
rect 12575 19468 14464 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 14608 19468 15117 19496
rect 14608 19456 14614 19468
rect 15105 19465 15117 19468
rect 15151 19465 15163 19499
rect 15105 19459 15163 19465
rect 16206 19456 16212 19508
rect 16264 19456 16270 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 17589 19499 17647 19505
rect 17589 19496 17601 19499
rect 16724 19468 17601 19496
rect 16724 19456 16730 19468
rect 17589 19465 17601 19468
rect 17635 19465 17647 19499
rect 17589 19459 17647 19465
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 18012 19468 19257 19496
rect 18012 19456 18018 19468
rect 19245 19465 19257 19468
rect 19291 19465 19303 19499
rect 19245 19459 19303 19465
rect 20349 19499 20407 19505
rect 20349 19465 20361 19499
rect 20395 19496 20407 19499
rect 22370 19496 22376 19508
rect 20395 19468 22376 19496
rect 20395 19465 20407 19468
rect 20349 19459 20407 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 22465 19499 22523 19505
rect 22465 19465 22477 19499
rect 22511 19496 22523 19499
rect 22738 19496 22744 19508
rect 22511 19468 22744 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 23382 19456 23388 19508
rect 23440 19456 23446 19508
rect 3786 19428 3792 19440
rect 2240 19400 3792 19428
rect 2240 19369 2268 19400
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 3970 19388 3976 19440
rect 4028 19428 4034 19440
rect 5074 19428 5080 19440
rect 4028 19400 4384 19428
rect 4028 19388 4034 19400
rect 2087 19332 2176 19360
rect 2225 19363 2283 19369
rect 2087 19329 2099 19332
rect 2041 19323 2099 19329
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 2314 19320 2320 19372
rect 2372 19320 2378 19372
rect 2682 19320 2688 19372
rect 2740 19360 2746 19372
rect 2902 19363 2960 19369
rect 2902 19360 2914 19363
rect 2740 19332 2914 19360
rect 2740 19320 2746 19332
rect 2902 19329 2914 19332
rect 2948 19329 2960 19363
rect 2902 19323 2960 19329
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4154 19360 4160 19372
rect 4111 19332 4160 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4356 19369 4384 19400
rect 4816 19400 5080 19428
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 1762 19252 1768 19304
rect 1820 19252 1826 19304
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 2648 19264 3433 19292
rect 2648 19252 2654 19264
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3421 19255 3479 19261
rect 2038 19184 2044 19236
rect 2096 19224 2102 19236
rect 3329 19227 3387 19233
rect 3329 19224 3341 19227
rect 2096 19196 3341 19224
rect 2096 19184 2102 19196
rect 3329 19193 3341 19196
rect 3375 19193 3387 19227
rect 4816 19224 4844 19400
rect 5074 19388 5080 19400
rect 5132 19388 5138 19440
rect 5721 19431 5779 19437
rect 5721 19397 5733 19431
rect 5767 19428 5779 19431
rect 6086 19428 6092 19440
rect 5767 19400 6092 19428
rect 5767 19397 5779 19400
rect 5721 19391 5779 19397
rect 6086 19388 6092 19400
rect 6144 19388 6150 19440
rect 7374 19388 7380 19440
rect 7432 19428 7438 19440
rect 9766 19428 9772 19440
rect 7432 19400 9772 19428
rect 7432 19388 7438 19400
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 9861 19431 9919 19437
rect 9861 19397 9873 19431
rect 9907 19428 9919 19431
rect 13081 19431 13139 19437
rect 9907 19400 13032 19428
rect 9907 19397 9919 19400
rect 9861 19391 9919 19397
rect 4982 19320 4988 19372
rect 5040 19320 5046 19372
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 5184 19292 5212 19323
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 5442 19360 5448 19372
rect 5316 19332 5448 19360
rect 5316 19320 5322 19332
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5905 19363 5963 19369
rect 5905 19360 5917 19363
rect 5592 19332 5917 19360
rect 5592 19320 5598 19332
rect 5905 19329 5917 19332
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6178 19360 6184 19372
rect 6043 19332 6184 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6178 19320 6184 19332
rect 6236 19320 6242 19372
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7466 19360 7472 19372
rect 7055 19332 7472 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 7650 19320 7656 19372
rect 7708 19360 7714 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7708 19332 7849 19360
rect 7708 19320 7714 19332
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 8938 19320 8944 19372
rect 8996 19320 9002 19372
rect 9122 19320 9128 19372
rect 9180 19320 9186 19372
rect 9214 19320 9220 19372
rect 9272 19320 9278 19372
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 9456 19332 10517 19360
rect 9456 19320 9462 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10686 19360 10692 19372
rect 10505 19323 10563 19329
rect 10612 19332 10692 19360
rect 6546 19292 6552 19304
rect 5184 19264 6552 19292
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 10318 19292 10324 19304
rect 8159 19264 10324 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 4985 19227 5043 19233
rect 4985 19224 4997 19227
rect 4816 19196 4997 19224
rect 3329 19187 3387 19193
rect 4985 19193 4997 19196
rect 5031 19193 5043 19227
rect 7193 19227 7251 19233
rect 7193 19224 7205 19227
rect 4985 19187 5043 19193
rect 5460 19196 7205 19224
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3602 19156 3608 19168
rect 3016 19128 3608 19156
rect 3016 19116 3022 19128
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3694 19116 3700 19168
rect 3752 19156 3758 19168
rect 5074 19156 5080 19168
rect 3752 19128 5080 19156
rect 3752 19116 3758 19128
rect 5074 19116 5080 19128
rect 5132 19156 5138 19168
rect 5460 19156 5488 19196
rect 7193 19193 7205 19196
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 7466 19184 7472 19236
rect 7524 19224 7530 19236
rect 7524 19196 9352 19224
rect 7524 19184 7530 19196
rect 5132 19128 5488 19156
rect 5132 19116 5138 19128
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5721 19159 5779 19165
rect 5721 19156 5733 19159
rect 5592 19128 5733 19156
rect 5592 19116 5598 19128
rect 5721 19125 5733 19128
rect 5767 19125 5779 19159
rect 5721 19119 5779 19125
rect 6086 19116 6092 19168
rect 6144 19156 6150 19168
rect 8202 19156 8208 19168
rect 6144 19128 8208 19156
rect 6144 19116 6150 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 9324 19156 9352 19196
rect 9398 19184 9404 19236
rect 9456 19224 9462 19236
rect 10612 19224 10640 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11011 19332 11045 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 10778 19252 10784 19304
rect 10836 19252 10842 19304
rect 10980 19292 11008 19323
rect 11606 19320 11612 19372
rect 11664 19360 11670 19372
rect 12253 19363 12311 19369
rect 12253 19360 12265 19363
rect 11664 19332 12265 19360
rect 11664 19320 11670 19332
rect 12253 19329 12265 19332
rect 12299 19329 12311 19363
rect 13004 19360 13032 19400
rect 13081 19397 13093 19431
rect 13127 19428 13139 19431
rect 13170 19428 13176 19440
rect 13127 19400 13176 19428
rect 13127 19397 13139 19400
rect 13081 19391 13139 19397
rect 13170 19388 13176 19400
rect 13228 19388 13234 19440
rect 13262 19388 13268 19440
rect 13320 19437 13326 19440
rect 13320 19431 13339 19437
rect 13327 19397 13339 19431
rect 13320 19391 13339 19397
rect 13320 19388 13326 19391
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 13906 19428 13912 19440
rect 13596 19400 13912 19428
rect 13596 19388 13602 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 13998 19388 14004 19440
rect 14056 19428 14062 19440
rect 14114 19431 14172 19437
rect 14114 19428 14126 19431
rect 14056 19400 14126 19428
rect 14056 19388 14062 19400
rect 14114 19397 14126 19400
rect 14160 19397 14172 19431
rect 14114 19391 14172 19397
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 14737 19431 14795 19437
rect 14737 19428 14749 19431
rect 14700 19400 14749 19428
rect 14700 19388 14706 19400
rect 14737 19397 14749 19400
rect 14783 19397 14795 19431
rect 14737 19391 14795 19397
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 14953 19431 15011 19437
rect 14953 19428 14965 19431
rect 14884 19400 14965 19428
rect 14884 19388 14890 19400
rect 14953 19397 14965 19400
rect 14999 19428 15011 19431
rect 15470 19428 15476 19440
rect 14999 19400 15476 19428
rect 14999 19397 15011 19400
rect 14953 19391 15011 19397
rect 15470 19388 15476 19400
rect 15528 19388 15534 19440
rect 16390 19388 16396 19440
rect 16448 19428 16454 19440
rect 17126 19428 17132 19440
rect 16448 19400 17132 19428
rect 16448 19388 16454 19400
rect 17126 19388 17132 19400
rect 17184 19428 17190 19440
rect 17221 19431 17279 19437
rect 17221 19428 17233 19431
rect 17184 19400 17233 19428
rect 17184 19388 17190 19400
rect 17221 19397 17233 19400
rect 17267 19397 17279 19431
rect 17221 19391 17279 19397
rect 17437 19431 17495 19437
rect 17437 19397 17449 19431
rect 17483 19428 17495 19431
rect 17862 19428 17868 19440
rect 17483 19400 17868 19428
rect 17483 19397 17495 19400
rect 17437 19391 17495 19397
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 18138 19388 18144 19440
rect 18196 19428 18202 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 18196 19400 18889 19428
rect 18196 19388 18202 19400
rect 18877 19397 18889 19400
rect 18923 19397 18935 19431
rect 18877 19391 18935 19397
rect 18966 19388 18972 19440
rect 19024 19428 19030 19440
rect 19077 19431 19135 19437
rect 19077 19428 19089 19431
rect 19024 19400 19089 19428
rect 19024 19388 19030 19400
rect 19077 19397 19089 19400
rect 19123 19397 19135 19431
rect 19077 19391 19135 19397
rect 19886 19388 19892 19440
rect 19944 19428 19950 19440
rect 21450 19428 21456 19440
rect 19944 19400 21456 19428
rect 19944 19388 19950 19400
rect 21450 19388 21456 19400
rect 21508 19428 21514 19440
rect 22005 19431 22063 19437
rect 22005 19428 22017 19431
rect 21508 19400 22017 19428
rect 21508 19388 21514 19400
rect 22005 19397 22017 19400
rect 22051 19397 22063 19431
rect 22005 19391 22063 19397
rect 22925 19431 22983 19437
rect 22925 19397 22937 19431
rect 22971 19428 22983 19431
rect 23014 19428 23020 19440
rect 22971 19400 23020 19428
rect 22971 19397 22983 19400
rect 22925 19391 22983 19397
rect 23014 19388 23020 19400
rect 23072 19428 23078 19440
rect 23750 19428 23756 19440
rect 23072 19400 23756 19428
rect 23072 19388 23078 19400
rect 23750 19388 23756 19400
rect 23808 19388 23814 19440
rect 26786 19428 26792 19440
rect 24044 19400 26792 19428
rect 15654 19360 15660 19372
rect 13004 19332 15660 19360
rect 12253 19323 12311 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16206 19360 16212 19372
rect 15856 19332 16212 19360
rect 11146 19292 11152 19304
rect 10980 19264 11152 19292
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11296 19264 11897 19292
rect 11296 19252 11302 19264
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 11885 19255 11943 19261
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 12176 19224 12204 19255
rect 12342 19252 12348 19304
rect 12400 19301 12406 19304
rect 12400 19295 12428 19301
rect 12416 19261 12428 19295
rect 15856 19292 15884 19332
rect 16206 19320 16212 19332
rect 16264 19320 16270 19372
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 17586 19360 17592 19372
rect 16347 19332 17592 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18046 19360 18052 19372
rect 17828 19332 18052 19360
rect 17828 19320 17834 19332
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 18231 19363 18289 19369
rect 18231 19329 18243 19363
rect 18277 19329 18289 19363
rect 18231 19323 18289 19329
rect 12400 19255 12428 19261
rect 14200 19264 15884 19292
rect 12400 19252 12406 19255
rect 9456 19196 10640 19224
rect 11348 19196 12204 19224
rect 9456 19184 9462 19196
rect 11348 19168 11376 19196
rect 12894 19184 12900 19236
rect 12952 19224 12958 19236
rect 14200 19224 14228 19264
rect 15930 19252 15936 19304
rect 15988 19252 15994 19304
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18248 19292 18276 19323
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 18656 19332 20821 19360
rect 18656 19320 18662 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21082 19360 21088 19372
rect 21039 19332 21088 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21928 19332 22094 19360
rect 18196 19264 18276 19292
rect 18196 19252 18202 19264
rect 12952 19196 14228 19224
rect 14277 19227 14335 19233
rect 12952 19184 12958 19196
rect 14277 19193 14289 19227
rect 14323 19224 14335 19227
rect 16025 19227 16083 19233
rect 16025 19224 16037 19227
rect 14323 19196 16037 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 16025 19193 16037 19196
rect 16071 19193 16083 19227
rect 18248 19224 18276 19264
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19292 18475 19295
rect 19334 19292 19340 19304
rect 18463 19264 19340 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 20622 19292 20628 19304
rect 20088 19264 20628 19292
rect 20088 19224 20116 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 21174 19252 21180 19304
rect 21232 19252 21238 19304
rect 21266 19252 21272 19304
rect 21324 19292 21330 19304
rect 21928 19292 21956 19332
rect 21324 19264 21956 19292
rect 22066 19292 22094 19332
rect 24044 19301 24072 19400
rect 26786 19388 26792 19400
rect 26844 19388 26850 19440
rect 24302 19369 24308 19372
rect 24285 19363 24308 19369
rect 24285 19329 24297 19363
rect 24285 19323 24308 19329
rect 24302 19320 24308 19323
rect 24360 19320 24366 19372
rect 24029 19295 24087 19301
rect 22066 19264 23336 19292
rect 21324 19252 21330 19264
rect 23308 19236 23336 19264
rect 24029 19261 24041 19295
rect 24075 19261 24087 19295
rect 24029 19255 24087 19261
rect 18248 19196 20116 19224
rect 16025 19187 16083 19193
rect 20162 19184 20168 19236
rect 20220 19184 20226 19236
rect 22281 19227 22339 19233
rect 22281 19193 22293 19227
rect 22327 19193 22339 19227
rect 22281 19187 22339 19193
rect 9490 19156 9496 19168
rect 9324 19128 9496 19156
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 11330 19156 11336 19168
rect 10744 19128 11336 19156
rect 10744 19116 10750 19128
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 13262 19116 13268 19168
rect 13320 19116 13326 19168
rect 13446 19116 13452 19168
rect 13504 19116 13510 19168
rect 14090 19116 14096 19168
rect 14148 19116 14154 19168
rect 14918 19116 14924 19168
rect 14976 19116 14982 19168
rect 15562 19116 15568 19168
rect 15620 19116 15626 19168
rect 15838 19116 15844 19168
rect 15896 19116 15902 19168
rect 17405 19159 17463 19165
rect 17405 19125 17417 19159
rect 17451 19156 17463 19159
rect 17494 19156 17500 19168
rect 17451 19128 17500 19156
rect 17451 19125 17463 19128
rect 17405 19119 17463 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18598 19156 18604 19168
rect 18104 19128 18604 19156
rect 18104 19116 18110 19128
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 20898 19156 20904 19168
rect 19107 19128 20904 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 22296 19156 22324 19187
rect 23290 19184 23296 19236
rect 23348 19184 23354 19236
rect 23566 19184 23572 19236
rect 23624 19224 23630 19236
rect 28166 19224 28172 19236
rect 23624 19196 24072 19224
rect 23624 19184 23630 19196
rect 23842 19156 23848 19168
rect 21048 19128 23848 19156
rect 21048 19116 21054 19128
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 24044 19156 24072 19196
rect 24964 19196 28172 19224
rect 24964 19156 24992 19196
rect 28166 19184 28172 19196
rect 28224 19184 28230 19236
rect 24044 19128 24992 19156
rect 25038 19116 25044 19168
rect 25096 19156 25102 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 25096 19128 25421 19156
rect 25096 19116 25102 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25409 19119 25467 19125
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 2915 18924 3740 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 3712 18884 3740 18924
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 4212 18924 5365 18952
rect 4212 18912 4218 18924
rect 5353 18921 5365 18924
rect 5399 18921 5411 18955
rect 7466 18952 7472 18964
rect 5353 18915 5411 18921
rect 6764 18924 7472 18952
rect 4246 18884 4252 18896
rect 1627 18856 3188 18884
rect 3712 18856 4252 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 2222 18816 2228 18828
rect 1872 18788 2228 18816
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 1872 18757 1900 18788
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2590 18748 2596 18760
rect 2179 18720 2596 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 1872 18624 1900 18711
rect 1854 18572 1860 18624
rect 1912 18572 1918 18624
rect 2056 18612 2084 18711
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 3050 18708 3056 18760
rect 3108 18708 3114 18760
rect 3160 18757 3188 18856
rect 4246 18844 4252 18856
rect 4304 18844 4310 18896
rect 4338 18844 4344 18896
rect 4396 18844 4402 18896
rect 4430 18844 4436 18896
rect 4488 18884 4494 18896
rect 4982 18884 4988 18896
rect 4488 18856 4988 18884
rect 4488 18844 4494 18856
rect 4982 18844 4988 18856
rect 5040 18884 5046 18896
rect 6764 18884 6792 18924
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 7742 18912 7748 18964
rect 7800 18912 7806 18964
rect 9674 18912 9680 18964
rect 9732 18912 9738 18964
rect 10318 18912 10324 18964
rect 10376 18952 10382 18964
rect 13081 18955 13139 18961
rect 13081 18952 13093 18955
rect 10376 18924 13093 18952
rect 10376 18912 10382 18924
rect 13081 18921 13093 18924
rect 13127 18952 13139 18955
rect 13814 18952 13820 18964
rect 13127 18924 13820 18952
rect 13127 18921 13139 18924
rect 13081 18915 13139 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14645 18955 14703 18961
rect 14645 18921 14657 18955
rect 14691 18952 14703 18955
rect 16758 18952 16764 18964
rect 14691 18924 16764 18952
rect 14691 18921 14703 18924
rect 14645 18915 14703 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 21174 18952 21180 18964
rect 19300 18924 21180 18952
rect 19300 18912 19306 18924
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 21634 18912 21640 18964
rect 21692 18912 21698 18964
rect 24946 18952 24952 18964
rect 22066 18924 24952 18952
rect 5040 18856 6792 18884
rect 5040 18844 5046 18856
rect 6822 18844 6828 18896
rect 6880 18844 6886 18896
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 8846 18884 8852 18896
rect 7892 18856 8852 18884
rect 7892 18844 7898 18856
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 11333 18887 11391 18893
rect 11333 18853 11345 18887
rect 11379 18884 11391 18887
rect 11606 18884 11612 18896
rect 11379 18856 11612 18884
rect 11379 18853 11391 18856
rect 11333 18847 11391 18853
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 11974 18844 11980 18896
rect 12032 18884 12038 18896
rect 12069 18887 12127 18893
rect 12069 18884 12081 18887
rect 12032 18856 12081 18884
rect 12032 18844 12038 18856
rect 12069 18853 12081 18856
rect 12115 18853 12127 18887
rect 12069 18847 12127 18853
rect 16206 18844 16212 18896
rect 16264 18884 16270 18896
rect 16577 18887 16635 18893
rect 16577 18884 16589 18887
rect 16264 18856 16589 18884
rect 16264 18844 16270 18856
rect 16577 18853 16589 18856
rect 16623 18884 16635 18887
rect 16850 18884 16856 18896
rect 16623 18856 16856 18884
rect 16623 18853 16635 18856
rect 16577 18847 16635 18853
rect 16850 18844 16856 18856
rect 16908 18884 16914 18896
rect 18598 18884 18604 18896
rect 16908 18856 18604 18884
rect 16908 18844 16914 18856
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 22066 18884 22094 18924
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 26789 18955 26847 18961
rect 26789 18952 26801 18955
rect 25056 18924 26801 18952
rect 18708 18856 22094 18884
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4617 18819 4675 18825
rect 4617 18816 4629 18819
rect 4212 18788 4629 18816
rect 4212 18776 4218 18788
rect 4617 18785 4629 18788
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 4801 18819 4859 18825
rect 4801 18785 4813 18819
rect 4847 18816 4859 18819
rect 6730 18816 6736 18828
rect 4847 18788 6736 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 6840 18816 6868 18844
rect 6840 18788 9674 18816
rect 3145 18751 3203 18757
rect 3145 18717 3157 18751
rect 3191 18717 3203 18751
rect 3145 18711 3203 18717
rect 3326 18708 3332 18760
rect 3384 18708 3390 18760
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18748 3479 18751
rect 3786 18748 3792 18760
rect 3467 18720 3792 18748
rect 3467 18717 3479 18720
rect 3421 18711 3479 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4304 18720 4537 18748
rect 4304 18708 4310 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4890 18708 4896 18760
rect 4948 18748 4954 18760
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 4948 18720 5549 18748
rect 4948 18708 4954 18720
rect 5537 18717 5549 18720
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18748 5871 18751
rect 6178 18748 6184 18760
rect 5859 18720 6184 18748
rect 5859 18717 5871 18720
rect 5813 18711 5871 18717
rect 2774 18640 2780 18692
rect 2832 18680 2838 18692
rect 4724 18680 4752 18708
rect 2832 18652 4752 18680
rect 5552 18680 5580 18711
rect 6178 18708 6184 18720
rect 6236 18748 6242 18760
rect 6638 18748 6644 18760
rect 6236 18720 6644 18748
rect 6236 18708 6242 18720
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 6840 18757 6868 18788
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 7524 18720 7941 18748
rect 7524 18708 7530 18720
rect 7929 18717 7941 18720
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 5626 18680 5632 18692
rect 5552 18652 5632 18680
rect 2832 18640 2838 18652
rect 5626 18640 5632 18652
rect 5684 18680 5690 18692
rect 6086 18680 6092 18692
rect 5684 18652 6092 18680
rect 5684 18640 5690 18652
rect 6086 18640 6092 18652
rect 6144 18640 6150 18692
rect 7101 18683 7159 18689
rect 7101 18649 7113 18683
rect 7147 18680 7159 18683
rect 7190 18680 7196 18692
rect 7147 18652 7196 18680
rect 7147 18649 7159 18652
rect 7101 18643 7159 18649
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 7944 18680 7972 18711
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 9214 18748 9220 18760
rect 8260 18720 9220 18748
rect 8260 18708 8266 18720
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 9646 18748 9674 18788
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10594 18816 10600 18828
rect 9916 18788 10600 18816
rect 9916 18776 9922 18788
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18816 10747 18819
rect 11054 18816 11060 18828
rect 10735 18788 11060 18816
rect 10735 18785 10747 18788
rect 10689 18779 10747 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11174 18819 11232 18825
rect 11174 18785 11186 18819
rect 11220 18816 11232 18819
rect 11220 18788 11392 18816
rect 11220 18785 11232 18788
rect 11174 18779 11232 18785
rect 10502 18748 10508 18760
rect 9646 18720 10508 18748
rect 10502 18708 10508 18720
rect 10560 18748 10566 18760
rect 11364 18748 11392 18788
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11572 18788 11805 18816
rect 11572 18776 11578 18788
rect 11793 18785 11805 18788
rect 11839 18816 11851 18819
rect 11882 18816 11888 18828
rect 11839 18788 11888 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 18708 18816 18736 18856
rect 23290 18844 23296 18896
rect 23348 18884 23354 18896
rect 25056 18884 25084 18924
rect 26789 18921 26801 18924
rect 26835 18921 26847 18955
rect 26789 18915 26847 18921
rect 23348 18856 25084 18884
rect 23348 18844 23354 18856
rect 12308 18788 14688 18816
rect 12308 18776 12314 18788
rect 10560 18720 11392 18748
rect 10560 18708 10566 18720
rect 8938 18680 8944 18692
rect 7944 18652 8944 18680
rect 8938 18640 8944 18652
rect 8996 18640 9002 18692
rect 9309 18683 9367 18689
rect 9309 18649 9321 18683
rect 9355 18649 9367 18683
rect 9309 18643 9367 18649
rect 9493 18683 9551 18689
rect 9493 18649 9505 18683
rect 9539 18680 9551 18683
rect 10778 18680 10784 18692
rect 9539 18652 10784 18680
rect 9539 18649 9551 18652
rect 9493 18643 9551 18649
rect 2866 18612 2872 18624
rect 2056 18584 2872 18612
rect 2866 18572 2872 18584
rect 2924 18612 2930 18624
rect 5258 18612 5264 18624
rect 2924 18584 5264 18612
rect 2924 18572 2930 18584
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 6178 18612 6184 18624
rect 5776 18584 6184 18612
rect 5776 18572 5782 18584
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7800 18584 8125 18612
rect 7800 18572 7806 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 9324 18612 9352 18643
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 11364 18680 11392 18720
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 13998 18748 14004 18760
rect 11664 18720 14004 18748
rect 11664 18708 11670 18720
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14660 18757 14688 18788
rect 17144 18788 18736 18816
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15378 18748 15384 18760
rect 15335 18720 15384 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 12342 18680 12348 18692
rect 11364 18652 12348 18680
rect 12342 18640 12348 18652
rect 12400 18640 12406 18692
rect 12897 18683 12955 18689
rect 12897 18649 12909 18683
rect 12943 18680 12955 18683
rect 12986 18680 12992 18692
rect 12943 18652 12992 18680
rect 12943 18649 12955 18652
rect 12897 18643 12955 18649
rect 12986 18640 12992 18652
rect 13044 18640 13050 18692
rect 14274 18680 14280 18692
rect 13280 18652 14280 18680
rect 10134 18612 10140 18624
rect 9324 18584 10140 18612
rect 8113 18575 8171 18581
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10744 18584 10977 18612
rect 10744 18572 10750 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 11057 18615 11115 18621
rect 11057 18581 11069 18615
rect 11103 18612 11115 18615
rect 11146 18612 11152 18624
rect 11103 18584 11152 18612
rect 11103 18581 11115 18584
rect 11057 18575 11115 18581
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 12253 18615 12311 18621
rect 12253 18612 12265 18615
rect 11480 18584 12265 18612
rect 11480 18572 11486 18584
rect 12253 18581 12265 18584
rect 12299 18581 12311 18615
rect 12253 18575 12311 18581
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13078 18612 13084 18624
rect 13136 18621 13142 18624
rect 13280 18621 13308 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 14369 18683 14427 18689
rect 14369 18649 14381 18683
rect 14415 18680 14427 18683
rect 14458 18680 14464 18692
rect 14415 18652 14464 18680
rect 14415 18649 14427 18652
rect 14369 18643 14427 18649
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 14568 18680 14596 18711
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 16390 18708 16396 18760
rect 16448 18708 16454 18760
rect 17144 18757 17172 18788
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17862 18748 17868 18760
rect 17543 18720 17868 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18708 18757 18736 18788
rect 18877 18819 18935 18825
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 20714 18816 20720 18828
rect 18923 18788 20720 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 20824 18788 22094 18816
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18104 18720 18521 18748
rect 18104 18708 18110 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19392 18720 19717 18748
rect 19392 18708 19398 18720
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 15194 18680 15200 18692
rect 14568 18652 15200 18680
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 17405 18683 17463 18689
rect 17405 18649 17417 18683
rect 17451 18680 17463 18683
rect 19812 18680 19840 18711
rect 19886 18708 19892 18760
rect 19944 18708 19950 18760
rect 20162 18708 20168 18760
rect 20220 18708 20226 18760
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20824 18748 20852 18788
rect 20404 18720 20852 18748
rect 20404 18708 20410 18720
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21358 18748 21364 18760
rect 20956 18720 21364 18748
rect 20956 18708 20962 18720
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 20254 18680 20260 18692
rect 17451 18652 17954 18680
rect 19812 18652 20260 18680
rect 17451 18649 17463 18652
rect 17405 18643 17463 18649
rect 13136 18615 13155 18621
rect 12860 18584 13084 18612
rect 12860 18572 12866 18584
rect 13078 18572 13084 18584
rect 13143 18581 13155 18615
rect 13136 18575 13155 18581
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18581 13323 18615
rect 13265 18575 13323 18581
rect 13136 18572 13142 18575
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 14829 18615 14887 18621
rect 14829 18612 14841 18615
rect 13688 18584 14841 18612
rect 13688 18572 13694 18584
rect 14829 18581 14841 18584
rect 14875 18581 14887 18615
rect 14829 18575 14887 18581
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 15473 18615 15531 18621
rect 15473 18612 15485 18615
rect 15344 18584 15485 18612
rect 15344 18572 15350 18584
rect 15473 18581 15485 18584
rect 15519 18612 15531 18615
rect 17126 18612 17132 18624
rect 15519 18584 17132 18612
rect 15519 18581 15531 18584
rect 15473 18575 15531 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17678 18572 17684 18624
rect 17736 18572 17742 18624
rect 17926 18612 17954 18652
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 21174 18640 21180 18692
rect 21232 18680 21238 18692
rect 21453 18683 21511 18689
rect 21453 18680 21465 18683
rect 21232 18652 21465 18680
rect 21232 18640 21238 18652
rect 21453 18649 21465 18652
rect 21499 18649 21511 18683
rect 21453 18643 21511 18649
rect 21669 18683 21727 18689
rect 21669 18649 21681 18683
rect 21715 18680 21727 18683
rect 21910 18680 21916 18692
rect 21715 18652 21916 18680
rect 21715 18649 21727 18652
rect 21669 18643 21727 18649
rect 18690 18612 18696 18624
rect 17926 18584 18696 18612
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19426 18572 19432 18624
rect 19484 18572 19490 18624
rect 20073 18615 20131 18621
rect 20073 18581 20085 18615
rect 20119 18612 20131 18615
rect 20806 18612 20812 18624
rect 20119 18584 20812 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 21684 18612 21712 18643
rect 21910 18640 21916 18652
rect 21968 18640 21974 18692
rect 22066 18680 22094 18788
rect 24394 18776 24400 18828
rect 24452 18816 24458 18828
rect 25130 18816 25136 18828
rect 24452 18788 25136 18816
rect 24452 18776 24458 18788
rect 25130 18776 25136 18788
rect 25188 18816 25194 18828
rect 25409 18819 25467 18825
rect 25409 18816 25421 18819
rect 25188 18788 25421 18816
rect 25188 18776 25194 18788
rect 25409 18785 25421 18788
rect 25455 18785 25467 18819
rect 25409 18779 25467 18785
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18748 22339 18751
rect 22830 18748 22836 18760
rect 22327 18720 22836 18748
rect 22327 18717 22339 18720
rect 22281 18711 22339 18717
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 23532 18720 24777 18748
rect 23532 18708 23538 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 22554 18689 22560 18692
rect 22526 18683 22560 18689
rect 22066 18652 22416 18680
rect 21416 18584 21712 18612
rect 21821 18615 21879 18621
rect 21416 18572 21422 18584
rect 21821 18581 21833 18615
rect 21867 18612 21879 18615
rect 22094 18612 22100 18624
rect 21867 18584 22100 18612
rect 21867 18581 21879 18584
rect 21821 18575 21879 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 22388 18612 22416 18652
rect 22526 18649 22538 18683
rect 22526 18643 22560 18649
rect 22554 18640 22560 18643
rect 22612 18640 22618 18692
rect 25654 18683 25712 18689
rect 25654 18680 25666 18683
rect 24780 18652 25666 18680
rect 23566 18612 23572 18624
rect 22388 18584 23572 18612
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 23658 18572 23664 18624
rect 23716 18572 23722 18624
rect 24581 18615 24639 18621
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 24780 18612 24808 18652
rect 25654 18649 25666 18652
rect 25700 18649 25712 18683
rect 25654 18643 25712 18649
rect 24627 18584 24808 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 2130 18368 2136 18420
rect 2188 18368 2194 18420
rect 4522 18368 4528 18420
rect 4580 18368 4586 18420
rect 4982 18408 4988 18420
rect 4724 18380 4988 18408
rect 3053 18343 3111 18349
rect 3053 18309 3065 18343
rect 3099 18340 3111 18343
rect 3694 18340 3700 18352
rect 3099 18312 3700 18340
rect 3099 18309 3111 18312
rect 3053 18303 3111 18309
rect 3694 18300 3700 18312
rect 3752 18300 3758 18352
rect 4540 18340 4568 18368
rect 4724 18349 4752 18380
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5350 18368 5356 18420
rect 5408 18408 5414 18420
rect 5408 18380 5764 18408
rect 5408 18368 5414 18380
rect 4264 18312 4568 18340
rect 4617 18343 4675 18349
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2056 18204 2084 18235
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 2682 18272 2688 18284
rect 2464 18244 2688 18272
rect 2464 18232 2470 18244
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 2866 18281 2872 18284
rect 2833 18275 2872 18281
rect 2833 18241 2845 18275
rect 2833 18235 2872 18241
rect 2866 18232 2872 18235
rect 2924 18232 2930 18284
rect 2958 18232 2964 18284
rect 3016 18232 3022 18284
rect 3191 18275 3249 18281
rect 3191 18241 3203 18275
rect 3237 18272 3249 18275
rect 4264 18272 4292 18312
rect 4617 18309 4629 18343
rect 4663 18309 4675 18343
rect 4617 18303 4675 18309
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18309 4767 18343
rect 4709 18303 4767 18309
rect 3237 18244 4292 18272
rect 3237 18241 3249 18244
rect 3191 18235 3249 18241
rect 4338 18232 4344 18284
rect 4396 18232 4402 18284
rect 4522 18281 4528 18284
rect 4489 18275 4528 18281
rect 4489 18241 4501 18275
rect 4489 18235 4528 18241
rect 4522 18232 4528 18235
rect 4580 18232 4586 18284
rect 4632 18216 4660 18303
rect 4890 18281 4896 18284
rect 4845 18275 4896 18281
rect 4845 18241 4857 18275
rect 4891 18241 4896 18275
rect 4845 18235 4896 18241
rect 4890 18232 4896 18235
rect 4948 18232 4954 18284
rect 5629 18275 5687 18281
rect 5629 18241 5641 18275
rect 5675 18241 5687 18275
rect 5736 18272 5764 18380
rect 7190 18368 7196 18420
rect 7248 18408 7254 18420
rect 8110 18408 8116 18420
rect 7248 18380 8116 18408
rect 7248 18368 7254 18380
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 8628 18380 10517 18408
rect 8628 18368 8634 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 13630 18408 13636 18420
rect 10652 18380 13636 18408
rect 10652 18368 10658 18380
rect 13630 18368 13636 18380
rect 13688 18368 13694 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 16942 18408 16948 18420
rect 14884 18380 16948 18408
rect 14884 18368 14890 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 17034 18368 17040 18420
rect 17092 18408 17098 18420
rect 18233 18411 18291 18417
rect 18233 18408 18245 18411
rect 17092 18380 18245 18408
rect 17092 18368 17098 18380
rect 18233 18377 18245 18380
rect 18279 18377 18291 18411
rect 18233 18371 18291 18377
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 20073 18411 20131 18417
rect 20073 18408 20085 18411
rect 18380 18380 20085 18408
rect 18380 18368 18386 18380
rect 20073 18377 20085 18380
rect 20119 18377 20131 18411
rect 20073 18371 20131 18377
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 23658 18408 23664 18420
rect 20680 18380 23664 18408
rect 20680 18368 20686 18380
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 23937 18411 23995 18417
rect 23937 18377 23949 18411
rect 23983 18377 23995 18411
rect 23937 18371 23995 18377
rect 5813 18343 5871 18349
rect 5813 18309 5825 18343
rect 5859 18340 5871 18343
rect 11974 18340 11980 18352
rect 5859 18312 11980 18340
rect 5859 18309 5871 18312
rect 5813 18303 5871 18309
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 12250 18300 12256 18352
rect 12308 18300 12314 18352
rect 12342 18300 12348 18352
rect 12400 18300 12406 18352
rect 12434 18300 12440 18352
rect 12492 18300 12498 18352
rect 13354 18300 13360 18352
rect 13412 18340 13418 18352
rect 14645 18343 14703 18349
rect 14645 18340 14657 18343
rect 13412 18312 14657 18340
rect 13412 18300 13418 18312
rect 14645 18309 14657 18312
rect 14691 18309 14703 18343
rect 19426 18340 19432 18352
rect 14645 18303 14703 18309
rect 14844 18312 19432 18340
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 5736 18244 5917 18272
rect 5629 18235 5687 18241
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7282 18272 7288 18284
rect 6963 18244 7288 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 3602 18204 3608 18216
rect 2056 18176 3608 18204
rect 3602 18164 3608 18176
rect 3660 18164 3666 18216
rect 4614 18164 4620 18216
rect 4672 18164 4678 18216
rect 5445 18139 5503 18145
rect 5445 18136 5457 18139
rect 2746 18108 5457 18136
rect 1302 18028 1308 18080
rect 1360 18068 1366 18080
rect 2746 18068 2774 18108
rect 5445 18105 5457 18108
rect 5491 18105 5503 18139
rect 5644 18136 5672 18235
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 8110 18232 8116 18284
rect 8168 18232 8174 18284
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 8846 18232 8852 18284
rect 8904 18232 8910 18284
rect 9490 18232 9496 18284
rect 9548 18272 9554 18284
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9548 18244 9597 18272
rect 9548 18232 9554 18244
rect 9585 18241 9597 18244
rect 9631 18272 9643 18275
rect 9766 18272 9772 18284
rect 9631 18244 9772 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10134 18232 10140 18284
rect 10192 18232 10198 18284
rect 10318 18232 10324 18284
rect 10376 18232 10382 18284
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11422 18272 11428 18284
rect 11195 18244 11428 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 13262 18272 13268 18284
rect 12124 18244 13268 18272
rect 12124 18232 12130 18244
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 13538 18272 13544 18284
rect 13372 18244 13544 18272
rect 7098 18164 7104 18216
rect 7156 18164 7162 18216
rect 7300 18204 7328 18232
rect 13372 18216 13400 18244
rect 13538 18232 13544 18244
rect 13596 18272 13602 18284
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 13596 18244 13645 18272
rect 13596 18232 13602 18244
rect 13633 18241 13645 18244
rect 13679 18241 13691 18275
rect 13633 18235 13691 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 14182 18272 14188 18284
rect 14047 18244 14188 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14844 18281 14872 18312
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 20162 18340 20168 18352
rect 19720 18312 20168 18340
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15565 18275 15623 18281
rect 14967 18244 15332 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 7300 18176 9076 18204
rect 5902 18136 5908 18148
rect 5644 18108 5908 18136
rect 5445 18099 5503 18105
rect 5902 18096 5908 18108
rect 5960 18136 5966 18148
rect 6362 18136 6368 18148
rect 5960 18108 6368 18136
rect 5960 18096 5966 18108
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 1360 18040 2774 18068
rect 1360 18028 1366 18040
rect 3142 18028 3148 18080
rect 3200 18068 3206 18080
rect 3329 18071 3387 18077
rect 3329 18068 3341 18071
rect 3200 18040 3341 18068
rect 3200 18028 3206 18040
rect 3329 18037 3341 18040
rect 3375 18037 3387 18071
rect 3329 18031 3387 18037
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 4985 18071 5043 18077
rect 4985 18068 4997 18071
rect 4120 18040 4997 18068
rect 4120 18028 4126 18040
rect 4985 18037 4997 18040
rect 5031 18037 5043 18071
rect 7116 18068 7144 18164
rect 7742 18068 7748 18080
rect 7116 18040 7748 18068
rect 4985 18031 5043 18037
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8846 18068 8852 18080
rect 7892 18040 8852 18068
rect 7892 18028 7898 18040
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9048 18068 9076 18176
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11664 18176 11713 18204
rect 11664 18164 11670 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12894 18204 12900 18216
rect 11931 18176 12900 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13354 18164 13360 18216
rect 13412 18164 13418 18216
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14148 18176 15148 18204
rect 14148 18164 14154 18176
rect 9217 18139 9275 18145
rect 9217 18105 9229 18139
rect 9263 18136 9275 18139
rect 10965 18139 11023 18145
rect 9263 18108 10916 18136
rect 9263 18105 9275 18108
rect 9217 18099 9275 18105
rect 10686 18068 10692 18080
rect 9048 18040 10692 18068
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 10888 18068 10916 18108
rect 10965 18105 10977 18139
rect 11011 18136 11023 18139
rect 15010 18136 15016 18148
rect 11011 18108 15016 18136
rect 11011 18105 11023 18108
rect 10965 18099 11023 18105
rect 15010 18096 15016 18108
rect 15068 18096 15074 18148
rect 15120 18145 15148 18176
rect 15105 18139 15163 18145
rect 15105 18105 15117 18139
rect 15151 18105 15163 18139
rect 15304 18136 15332 18244
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15580 18204 15608 18235
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15712 18244 15761 18272
rect 15712 18232 15718 18244
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 17109 18275 17167 18281
rect 17109 18272 17121 18275
rect 16448 18244 17121 18272
rect 16448 18232 16454 18244
rect 17109 18241 17121 18244
rect 17155 18241 17167 18275
rect 17109 18235 17167 18241
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 18949 18275 19007 18281
rect 18949 18272 18961 18275
rect 17552 18244 18961 18272
rect 17552 18232 17558 18244
rect 18949 18241 18961 18244
rect 18995 18241 19007 18275
rect 18949 18235 19007 18241
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19720 18272 19748 18312
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 20809 18343 20867 18349
rect 20809 18309 20821 18343
rect 20855 18340 20867 18343
rect 21450 18340 21456 18352
rect 20855 18312 21456 18340
rect 20855 18309 20867 18312
rect 20809 18303 20867 18309
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 23952 18340 23980 18371
rect 26234 18368 26240 18420
rect 26292 18368 26298 18420
rect 23400 18312 23888 18340
rect 23952 18312 26464 18340
rect 19392 18244 19748 18272
rect 19392 18232 19398 18244
rect 19794 18232 19800 18284
rect 19852 18272 19858 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 19852 18244 22201 18272
rect 19852 18232 19858 18244
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 22833 18275 22891 18281
rect 22833 18272 22845 18275
rect 22189 18235 22247 18241
rect 22480 18244 22845 18272
rect 15436 18176 15608 18204
rect 15764 18176 16804 18204
rect 15436 18164 15442 18176
rect 15764 18136 15792 18176
rect 16114 18136 16120 18148
rect 15304 18108 15792 18136
rect 15856 18108 16120 18136
rect 15105 18099 15163 18105
rect 13538 18068 13544 18080
rect 10888 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13630 18028 13636 18080
rect 13688 18068 13694 18080
rect 14826 18068 14832 18080
rect 13688 18040 14832 18068
rect 13688 18028 13694 18040
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 14921 18071 14979 18077
rect 14921 18037 14933 18071
rect 14967 18068 14979 18071
rect 15856 18068 15884 18108
rect 16114 18096 16120 18108
rect 16172 18096 16178 18148
rect 14967 18040 15884 18068
rect 15933 18071 15991 18077
rect 14967 18037 14979 18040
rect 14921 18031 14979 18037
rect 15933 18037 15945 18071
rect 15979 18068 15991 18071
rect 16206 18068 16212 18080
rect 15979 18040 16212 18068
rect 15979 18037 15991 18040
rect 15933 18031 15991 18037
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16776 18068 16804 18176
rect 16850 18164 16856 18216
rect 16908 18164 16914 18216
rect 18598 18164 18604 18216
rect 18656 18204 18662 18216
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 18656 18176 18705 18204
rect 18656 18164 18662 18176
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 21269 18207 21327 18213
rect 20128 18176 21220 18204
rect 20128 18164 20134 18176
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21085 18139 21143 18145
rect 21085 18136 21097 18139
rect 20864 18108 21097 18136
rect 20864 18096 20870 18108
rect 21085 18105 21097 18108
rect 21131 18105 21143 18139
rect 21085 18099 21143 18105
rect 19334 18068 19340 18080
rect 16776 18040 19340 18068
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 21192 18068 21220 18176
rect 21269 18173 21281 18207
rect 21315 18204 21327 18207
rect 22480 18204 22508 18244
rect 22833 18241 22845 18244
rect 22879 18241 22891 18275
rect 22833 18235 22891 18241
rect 21315 18176 22508 18204
rect 21315 18173 21327 18176
rect 21269 18167 21327 18173
rect 22005 18139 22063 18145
rect 22005 18105 22017 18139
rect 22051 18136 22063 18139
rect 22462 18136 22468 18148
rect 22051 18108 22468 18136
rect 22051 18105 22063 18108
rect 22005 18099 22063 18105
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 23400 18136 23428 18312
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18272 23535 18275
rect 23750 18272 23756 18284
rect 23523 18244 23756 18272
rect 23523 18241 23535 18244
rect 23477 18235 23535 18241
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 23860 18272 23888 18312
rect 24118 18272 24124 18284
rect 23860 18244 24124 18272
rect 24118 18232 24124 18244
rect 24176 18232 24182 18284
rect 26436 18281 26464 18312
rect 24664 18275 24722 18281
rect 24664 18241 24676 18275
rect 24710 18272 24722 18275
rect 26421 18275 26479 18281
rect 24710 18244 26372 18272
rect 24710 18241 24722 18244
rect 24664 18235 24722 18241
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24394 18204 24400 18216
rect 23716 18176 24400 18204
rect 23716 18164 23722 18176
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 26344 18204 26372 18244
rect 26421 18241 26433 18275
rect 26467 18241 26479 18275
rect 26421 18235 26479 18241
rect 27430 18204 27436 18216
rect 26344 18176 27436 18204
rect 27430 18164 27436 18176
rect 27488 18164 27494 18216
rect 22664 18108 23428 18136
rect 23845 18139 23903 18145
rect 22554 18068 22560 18080
rect 21192 18040 22560 18068
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 22664 18077 22692 18108
rect 23845 18105 23857 18139
rect 23891 18136 23903 18139
rect 23934 18136 23940 18148
rect 23891 18108 23940 18136
rect 23891 18105 23903 18108
rect 23845 18099 23903 18105
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 22649 18071 22707 18077
rect 22649 18037 22661 18071
rect 22695 18037 22707 18071
rect 22649 18031 22707 18037
rect 22738 18028 22744 18080
rect 22796 18068 22802 18080
rect 25038 18068 25044 18080
rect 22796 18040 25044 18068
rect 22796 18028 22802 18040
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 25774 18028 25780 18080
rect 25832 18028 25838 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 1026 17824 1032 17876
rect 1084 17864 1090 17876
rect 2774 17864 2780 17876
rect 1084 17836 2780 17864
rect 1084 17824 1090 17836
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4154 17864 4160 17876
rect 3375 17836 4160 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 5534 17864 5540 17876
rect 4396 17836 5540 17864
rect 4396 17824 4402 17836
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 5626 17824 5632 17876
rect 5684 17824 5690 17876
rect 6454 17824 6460 17876
rect 6512 17824 6518 17876
rect 8294 17864 8300 17876
rect 6564 17836 8300 17864
rect 2685 17799 2743 17805
rect 2685 17765 2697 17799
rect 2731 17796 2743 17799
rect 3970 17796 3976 17808
rect 2731 17768 3976 17796
rect 2731 17765 2743 17768
rect 2685 17759 2743 17765
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 5718 17796 5724 17808
rect 4178 17768 5724 17796
rect 2148 17700 3372 17728
rect 2148 17669 2176 17700
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2133 17623 2191 17629
rect 2501 17663 2559 17669
rect 2501 17629 2513 17663
rect 2547 17660 2559 17663
rect 2590 17660 2596 17672
rect 2547 17632 2596 17660
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 2590 17620 2596 17632
rect 2648 17620 2654 17672
rect 3145 17663 3203 17669
rect 3145 17660 3157 17663
rect 2746 17632 3157 17660
rect 1854 17552 1860 17604
rect 1912 17592 1918 17604
rect 2317 17595 2375 17601
rect 2317 17592 2329 17595
rect 1912 17564 2329 17592
rect 1912 17552 1918 17564
rect 2317 17561 2329 17564
rect 2363 17561 2375 17595
rect 2317 17555 2375 17561
rect 2332 17524 2360 17555
rect 2406 17552 2412 17604
rect 2464 17552 2470 17604
rect 2746 17524 2774 17632
rect 3145 17629 3157 17632
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 3234 17620 3240 17672
rect 3292 17620 3298 17672
rect 2332 17496 2774 17524
rect 3344 17524 3372 17700
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 4178 17728 4206 17768
rect 5718 17756 5724 17768
rect 5776 17796 5782 17808
rect 6564 17796 6592 17836
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 12161 17867 12219 17873
rect 8444 17836 12128 17864
rect 8444 17824 8450 17836
rect 5776 17768 6592 17796
rect 5776 17756 5782 17768
rect 7006 17756 7012 17808
rect 7064 17796 7070 17808
rect 7834 17796 7840 17808
rect 7064 17768 7840 17796
rect 7064 17756 7070 17768
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 9858 17796 9864 17808
rect 8404 17768 9864 17796
rect 3476 17700 4206 17728
rect 4249 17731 4307 17737
rect 3476 17688 3482 17700
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 4338 17728 4344 17740
rect 4295 17700 4344 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 7466 17728 7472 17740
rect 6472 17700 7472 17728
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 3418 17552 3424 17604
rect 3476 17592 3482 17604
rect 3988 17592 4016 17623
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 5166 17660 5172 17672
rect 4948 17632 5172 17660
rect 4948 17620 4954 17632
rect 5166 17620 5172 17632
rect 5224 17660 5230 17672
rect 5445 17663 5503 17669
rect 5445 17660 5457 17663
rect 5224 17632 5457 17660
rect 5224 17620 5230 17632
rect 5445 17629 5457 17632
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 6472 17669 6500 17700
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 8404 17728 8432 17768
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 10229 17799 10287 17805
rect 10229 17765 10241 17799
rect 10275 17796 10287 17799
rect 10502 17796 10508 17808
rect 10275 17768 10508 17796
rect 10275 17765 10287 17768
rect 10229 17759 10287 17765
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 10686 17756 10692 17808
rect 10744 17796 10750 17808
rect 12100 17796 12128 17836
rect 12161 17833 12173 17867
rect 12207 17864 12219 17867
rect 12207 17836 12756 17864
rect 12207 17833 12219 17836
rect 12161 17827 12219 17833
rect 12728 17796 12756 17836
rect 12802 17824 12808 17876
rect 12860 17824 12866 17876
rect 13630 17864 13636 17876
rect 13296 17836 13636 17864
rect 13296 17796 13324 17836
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 13872 17836 14473 17864
rect 13872 17824 13878 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15436 17836 15792 17864
rect 15436 17824 15442 17836
rect 10744 17768 11560 17796
rect 12100 17768 12388 17796
rect 12728 17768 13324 17796
rect 14645 17799 14703 17805
rect 10744 17756 10750 17768
rect 9953 17731 10011 17737
rect 7668 17700 8432 17728
rect 8496 17700 9536 17728
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 5684 17632 6469 17660
rect 5684 17620 5690 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6730 17620 6736 17672
rect 6788 17620 6794 17672
rect 3476 17564 4016 17592
rect 3476 17552 3482 17564
rect 4062 17552 4068 17604
rect 4120 17592 4126 17604
rect 6546 17592 6552 17604
rect 4120 17564 6552 17592
rect 4120 17552 4126 17564
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 7190 17552 7196 17604
rect 7248 17592 7254 17604
rect 7377 17595 7435 17601
rect 7377 17592 7389 17595
rect 7248 17564 7389 17592
rect 7248 17552 7254 17564
rect 7377 17561 7389 17564
rect 7423 17561 7435 17595
rect 7377 17555 7435 17561
rect 7469 17595 7527 17601
rect 7469 17561 7481 17595
rect 7515 17592 7527 17595
rect 7668 17592 7696 17700
rect 8496 17672 8524 17700
rect 7742 17620 7748 17672
rect 7800 17620 7806 17672
rect 7834 17620 7840 17672
rect 7892 17620 7898 17672
rect 8478 17660 8484 17672
rect 7944 17632 8484 17660
rect 7515 17564 7696 17592
rect 7760 17592 7788 17620
rect 7944 17601 7972 17632
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 9508 17669 9536 17700
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 10318 17728 10324 17740
rect 9999 17700 10324 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 11422 17728 11428 17740
rect 10468 17700 11428 17728
rect 10468 17688 10474 17700
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 11532 17737 11560 17768
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17728 11575 17731
rect 11563 17700 11944 17728
rect 11563 17697 11575 17700
rect 11517 17691 11575 17697
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9674 17660 9680 17672
rect 9539 17632 9680 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 7929 17595 7987 17601
rect 7929 17592 7941 17595
rect 7760 17564 7941 17592
rect 7515 17561 7527 17564
rect 7469 17555 7527 17561
rect 7929 17561 7941 17564
rect 7975 17561 7987 17595
rect 7929 17555 7987 17561
rect 8021 17595 8079 17601
rect 8021 17561 8033 17595
rect 8067 17592 8079 17595
rect 8294 17592 8300 17604
rect 8067 17564 8300 17592
rect 8067 17561 8079 17564
rect 8021 17555 8079 17561
rect 8294 17552 8300 17564
rect 8352 17592 8358 17604
rect 9232 17592 9260 17623
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 9858 17620 9864 17672
rect 9916 17620 9922 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 10962 17660 10968 17672
rect 10919 17632 10968 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 9950 17592 9956 17604
rect 8352 17564 9956 17592
rect 8352 17552 8358 17564
rect 9950 17552 9956 17564
rect 10008 17552 10014 17604
rect 10796 17592 10824 17623
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 11054 17620 11060 17672
rect 11112 17660 11118 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11112 17632 11805 17660
rect 11112 17620 11118 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11916 17660 11944 17700
rect 11974 17688 11980 17740
rect 12032 17688 12038 17740
rect 12250 17660 12256 17672
rect 11916 17632 12256 17660
rect 11793 17623 11851 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12360 17660 12388 17768
rect 14645 17765 14657 17799
rect 14691 17796 14703 17799
rect 14691 17768 15608 17796
rect 14691 17765 14703 17768
rect 14645 17759 14703 17765
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 12584 17700 13369 17728
rect 12584 17688 12590 17700
rect 13357 17697 13369 17700
rect 13403 17728 13415 17731
rect 15194 17728 15200 17740
rect 13403 17700 15200 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 15580 17728 15608 17768
rect 15654 17756 15660 17808
rect 15712 17756 15718 17808
rect 15764 17796 15792 17836
rect 16390 17824 16396 17876
rect 16448 17824 16454 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 16500 17836 17233 17864
rect 16500 17796 16528 17836
rect 17221 17833 17233 17836
rect 17267 17864 17279 17867
rect 17770 17864 17776 17876
rect 17267 17836 17776 17864
rect 17267 17833 17279 17836
rect 17221 17827 17279 17833
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 18049 17867 18107 17873
rect 18049 17833 18061 17867
rect 18095 17864 18107 17867
rect 18782 17864 18788 17876
rect 18095 17836 18788 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 19794 17824 19800 17876
rect 19852 17824 19858 17876
rect 20441 17867 20499 17873
rect 20441 17833 20453 17867
rect 20487 17833 20499 17867
rect 20441 17827 20499 17833
rect 21637 17867 21695 17873
rect 21637 17833 21649 17867
rect 21683 17864 21695 17867
rect 21683 17836 23244 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 15764 17768 16528 17796
rect 16758 17756 16764 17808
rect 16816 17796 16822 17808
rect 19978 17796 19984 17808
rect 16816 17768 19984 17796
rect 16816 17756 16822 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 15580 17700 18153 17728
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 18233 17731 18291 17737
rect 18233 17697 18245 17731
rect 18279 17728 18291 17731
rect 20162 17728 20168 17740
rect 18279 17700 20168 17728
rect 18279 17697 18291 17700
rect 18233 17691 18291 17697
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 20456 17728 20484 17827
rect 22554 17756 22560 17808
rect 22612 17796 22618 17808
rect 23014 17796 23020 17808
rect 22612 17768 23020 17796
rect 22612 17756 22618 17768
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 23216 17796 23244 17836
rect 23842 17824 23848 17876
rect 23900 17864 23906 17876
rect 26326 17864 26332 17876
rect 23900 17836 26332 17864
rect 23900 17824 23906 17836
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 26786 17864 26792 17876
rect 26436 17836 26792 17864
rect 24302 17796 24308 17808
rect 23216 17768 24308 17796
rect 24302 17756 24308 17768
rect 24360 17756 24366 17808
rect 23934 17728 23940 17740
rect 20456 17700 23940 17728
rect 23934 17688 23940 17700
rect 23992 17688 23998 17740
rect 26436 17737 26464 17836
rect 26786 17824 26792 17836
rect 26844 17824 26850 17876
rect 27798 17756 27804 17808
rect 27856 17756 27862 17808
rect 26421 17731 26479 17737
rect 26421 17697 26433 17731
rect 26467 17697 26479 17731
rect 26421 17691 26479 17697
rect 12713 17663 12771 17669
rect 12713 17660 12725 17663
rect 12360 17632 12725 17660
rect 12713 17629 12725 17632
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 13320 17632 13553 17660
rect 13320 17620 13326 17632
rect 13541 17629 13553 17632
rect 13587 17629 13599 17663
rect 15010 17660 15016 17672
rect 14537 17635 15016 17660
rect 13541 17623 13599 17629
rect 14507 17632 15016 17635
rect 14507 17629 14565 17632
rect 11146 17592 11152 17604
rect 10796 17564 11152 17592
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 11422 17552 11428 17604
rect 11480 17592 11486 17604
rect 11885 17595 11943 17601
rect 11480 17564 11836 17592
rect 11480 17552 11486 17564
rect 4982 17524 4988 17536
rect 3344 17496 4988 17524
rect 4982 17484 4988 17496
rect 5040 17524 5046 17536
rect 5350 17524 5356 17536
rect 5040 17496 5356 17524
rect 5040 17484 5046 17496
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 6086 17484 6092 17536
rect 6144 17524 6150 17536
rect 6641 17527 6699 17533
rect 6641 17524 6653 17527
rect 6144 17496 6653 17524
rect 6144 17484 6150 17496
rect 6641 17493 6653 17496
rect 6687 17493 6699 17527
rect 6641 17487 6699 17493
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 9858 17524 9864 17536
rect 8904 17496 9864 17524
rect 8904 17484 8910 17496
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 11057 17527 11115 17533
rect 11057 17493 11069 17527
rect 11103 17524 11115 17527
rect 11698 17524 11704 17536
rect 11103 17496 11704 17524
rect 11103 17493 11115 17496
rect 11057 17487 11115 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 11808 17524 11836 17564
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 12342 17592 12348 17604
rect 11931 17564 12348 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 13964 17564 14289 17592
rect 13964 17552 13970 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14507 17595 14519 17629
rect 14553 17595 14565 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15212 17660 15240 17688
rect 15930 17660 15936 17672
rect 15212 17632 15936 17660
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 18322 17620 18328 17672
rect 18380 17620 18386 17672
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 19242 17660 19248 17672
rect 18555 17632 19248 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 14507 17589 14565 17595
rect 15289 17595 15347 17601
rect 14277 17555 14335 17561
rect 15289 17561 15301 17595
rect 15335 17561 15347 17595
rect 15289 17555 15347 17561
rect 12802 17524 12808 17536
rect 11808 17496 12808 17524
rect 12802 17484 12808 17496
rect 12860 17524 12866 17536
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 12860 17496 13737 17524
rect 12860 17484 12866 17496
rect 13725 17493 13737 17496
rect 13771 17493 13783 17527
rect 15304 17524 15332 17555
rect 16022 17552 16028 17604
rect 16080 17592 16086 17604
rect 16209 17595 16267 17601
rect 16209 17592 16221 17595
rect 16080 17564 16221 17592
rect 16080 17552 16086 17564
rect 16209 17561 16221 17564
rect 16255 17592 16267 17595
rect 16298 17592 16304 17604
rect 16255 17564 16304 17592
rect 16255 17561 16267 17564
rect 16209 17555 16267 17561
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 17126 17552 17132 17604
rect 17184 17552 17190 17604
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 17644 17564 18000 17592
rect 17644 17552 17650 17564
rect 15378 17524 15384 17536
rect 15304 17496 15384 17524
rect 13725 17487 13783 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 15654 17484 15660 17536
rect 15712 17524 15718 17536
rect 15749 17527 15807 17533
rect 15749 17524 15761 17527
rect 15712 17496 15761 17524
rect 15712 17484 15718 17496
rect 15749 17493 15761 17496
rect 15795 17493 15807 17527
rect 15749 17487 15807 17493
rect 16390 17484 16396 17536
rect 16448 17533 16454 17536
rect 16448 17527 16467 17533
rect 16455 17493 16467 17527
rect 16448 17487 16467 17493
rect 16448 17484 16454 17487
rect 16574 17484 16580 17536
rect 16632 17484 16638 17536
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17773 17527 17831 17533
rect 17773 17524 17785 17527
rect 16908 17496 17785 17524
rect 16908 17484 16914 17496
rect 17773 17493 17785 17496
rect 17819 17493 17831 17527
rect 17972 17524 18000 17564
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 18524 17592 18552 17623
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19518 17660 19524 17672
rect 19475 17632 19524 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19978 17620 19984 17672
rect 20036 17660 20042 17672
rect 21821 17663 21879 17669
rect 20036 17632 20760 17660
rect 20036 17620 20042 17632
rect 18104 17564 18552 17592
rect 18104 17552 18110 17564
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 18656 17564 19104 17592
rect 18656 17552 18662 17564
rect 18966 17524 18972 17536
rect 17972 17496 18972 17524
rect 17773 17487 17831 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19076 17524 19104 17564
rect 19610 17552 19616 17604
rect 19668 17552 19674 17604
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 20257 17595 20315 17601
rect 20257 17592 20269 17595
rect 20128 17564 20269 17592
rect 20128 17552 20134 17564
rect 20257 17561 20269 17564
rect 20303 17561 20315 17595
rect 20257 17555 20315 17561
rect 19242 17524 19248 17536
rect 19076 17496 19248 17524
rect 19242 17484 19248 17496
rect 19300 17524 19306 17536
rect 20457 17527 20515 17533
rect 20457 17524 20469 17527
rect 19300 17496 20469 17524
rect 19300 17484 19306 17496
rect 20457 17493 20469 17496
rect 20503 17493 20515 17527
rect 20457 17487 20515 17493
rect 20622 17484 20628 17536
rect 20680 17484 20686 17536
rect 20732 17524 20760 17632
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 22462 17660 22468 17672
rect 21867 17632 22468 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 22462 17620 22468 17632
rect 22520 17620 22526 17672
rect 24581 17663 24639 17669
rect 22664 17632 23704 17660
rect 21542 17552 21548 17604
rect 21600 17592 21606 17604
rect 22554 17592 22560 17604
rect 21600 17564 22560 17592
rect 21600 17552 21606 17564
rect 22554 17552 22560 17564
rect 22612 17552 22618 17604
rect 21450 17524 21456 17536
rect 20732 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17524 21514 17536
rect 22664 17524 22692 17632
rect 22741 17595 22799 17601
rect 22741 17561 22753 17595
rect 22787 17592 22799 17595
rect 22787 17564 22968 17592
rect 22787 17561 22799 17564
rect 22741 17555 22799 17561
rect 21508 17496 22692 17524
rect 21508 17484 21514 17496
rect 22830 17484 22836 17536
rect 22888 17484 22894 17536
rect 22940 17524 22968 17564
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 23477 17595 23535 17601
rect 23477 17592 23489 17595
rect 23072 17564 23489 17592
rect 23072 17552 23078 17564
rect 23477 17561 23489 17564
rect 23523 17561 23535 17595
rect 23477 17555 23535 17561
rect 23566 17524 23572 17536
rect 22940 17496 23572 17524
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 23676 17524 23704 17632
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 26436 17660 26464 17691
rect 24627 17632 26464 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 26510 17620 26516 17672
rect 26568 17660 26574 17672
rect 26677 17663 26735 17669
rect 26677 17660 26689 17663
rect 26568 17632 26689 17660
rect 26568 17620 26574 17632
rect 26677 17629 26689 17632
rect 26723 17629 26735 17663
rect 26677 17623 26735 17629
rect 24302 17552 24308 17604
rect 24360 17592 24366 17604
rect 24826 17595 24884 17601
rect 24826 17592 24838 17595
rect 24360 17564 24838 17592
rect 24360 17552 24366 17564
rect 24826 17561 24838 17564
rect 24872 17561 24884 17595
rect 24826 17555 24884 17561
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 23676 17496 25973 17524
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 28350 17524 28356 17536
rect 26200 17496 28356 17524
rect 26200 17484 26206 17496
rect 28350 17484 28356 17496
rect 28408 17484 28414 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 2280 17292 2605 17320
rect 2280 17280 2286 17292
rect 2593 17289 2605 17292
rect 2639 17289 2651 17323
rect 2593 17283 2651 17289
rect 2682 17280 2688 17332
rect 2740 17320 2746 17332
rect 4433 17323 4491 17329
rect 2740 17292 3832 17320
rect 2740 17280 2746 17292
rect 1673 17255 1731 17261
rect 1673 17221 1685 17255
rect 1719 17252 1731 17255
rect 3234 17252 3240 17264
rect 1719 17224 3240 17252
rect 1719 17221 1731 17224
rect 1673 17215 1731 17221
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2038 17184 2044 17196
rect 1811 17156 2044 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 1596 17116 1624 17147
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 2188 17156 2237 17184
rect 2188 17144 2194 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2314 17144 2320 17196
rect 2372 17190 2378 17196
rect 2409 17190 2467 17193
rect 2372 17187 2467 17190
rect 2372 17162 2421 17187
rect 2372 17144 2378 17162
rect 2409 17153 2421 17162
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2498 17144 2504 17196
rect 2556 17184 2562 17196
rect 3804 17193 3832 17292
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 5810 17320 5816 17332
rect 4479 17292 5816 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 5994 17320 6000 17332
rect 5951 17292 6000 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6604 17292 6653 17320
rect 6604 17280 6610 17292
rect 6641 17289 6653 17292
rect 6687 17289 6699 17323
rect 6641 17283 6699 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7432 17292 7849 17320
rect 7432 17280 7438 17292
rect 7837 17289 7849 17292
rect 7883 17320 7895 17323
rect 9214 17320 9220 17332
rect 7883 17292 9220 17320
rect 7883 17289 7895 17292
rect 7837 17283 7895 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10318 17320 10324 17332
rect 9824 17292 10324 17320
rect 9824 17280 9830 17292
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 12066 17320 12072 17332
rect 10919 17292 12072 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12526 17320 12532 17332
rect 12452 17292 12532 17320
rect 7558 17252 7564 17264
rect 3988 17224 7564 17252
rect 3988 17193 4016 17224
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 7653 17255 7711 17261
rect 7653 17221 7665 17255
rect 7699 17252 7711 17255
rect 8021 17255 8079 17261
rect 7699 17224 7880 17252
rect 7699 17221 7711 17224
rect 7653 17215 7711 17221
rect 3789 17187 3847 17193
rect 2556 17156 3740 17184
rect 2556 17144 2562 17156
rect 1946 17116 1952 17128
rect 1596 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2774 17076 2780 17128
rect 2832 17076 2838 17128
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17085 2927 17119
rect 3712 17116 3740 17156
rect 3789 17153 3801 17187
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 3937 17187 4016 17193
rect 3937 17153 3949 17187
rect 3983 17156 4016 17187
rect 4065 17187 4123 17193
rect 3983 17153 3995 17156
rect 3937 17147 3995 17153
rect 4065 17153 4077 17187
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 4080 17116 4108 17147
rect 4154 17144 4160 17196
rect 4212 17144 4218 17196
rect 4295 17187 4353 17193
rect 4295 17153 4307 17187
rect 4341 17184 4353 17187
rect 4706 17184 4712 17196
rect 4341 17156 4712 17184
rect 4341 17153 4353 17156
rect 4295 17147 4353 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4856 17156 4905 17184
rect 4856 17144 4862 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 4430 17116 4436 17128
rect 3712 17088 3980 17116
rect 4080 17088 4436 17116
rect 2869 17079 2927 17085
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 2884 16980 2912 17079
rect 3952 17048 3980 17088
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 5006 17048 5034 17147
rect 5074 17144 5080 17196
rect 5132 17144 5138 17196
rect 5258 17144 5264 17196
rect 5316 17144 5322 17196
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 5810 17184 5816 17196
rect 5644 17156 5816 17184
rect 5092 17116 5120 17144
rect 5644 17116 5672 17156
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 6512 17156 6561 17184
rect 6512 17144 6518 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7745 17187 7803 17193
rect 7745 17184 7757 17187
rect 7340 17156 7757 17184
rect 7340 17144 7346 17156
rect 7745 17153 7757 17156
rect 7791 17153 7803 17187
rect 7852 17184 7880 17224
rect 8021 17221 8033 17255
rect 8067 17252 8079 17255
rect 10962 17252 10968 17264
rect 8067 17224 10968 17252
rect 8067 17221 8079 17224
rect 8021 17215 8079 17221
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 12452 17261 12480 17292
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 12805 17323 12863 17329
rect 12805 17289 12817 17323
rect 12851 17320 12863 17323
rect 13722 17320 13728 17332
rect 12851 17292 13728 17320
rect 12851 17289 12863 17292
rect 12805 17283 12863 17289
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 14921 17323 14979 17329
rect 14921 17289 14933 17323
rect 14967 17320 14979 17323
rect 16298 17320 16304 17332
rect 14967 17292 16304 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16482 17280 16488 17332
rect 16540 17320 16546 17332
rect 19153 17323 19211 17329
rect 19153 17320 19165 17323
rect 16540 17292 19165 17320
rect 16540 17280 16546 17292
rect 19153 17289 19165 17292
rect 19199 17289 19211 17323
rect 19153 17283 19211 17289
rect 19306 17292 20116 17320
rect 12437 17255 12495 17261
rect 12437 17252 12449 17255
rect 11204 17224 12449 17252
rect 11204 17212 11210 17224
rect 12437 17221 12449 17224
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 12653 17255 12711 17261
rect 12653 17221 12665 17255
rect 12699 17252 12711 17255
rect 13170 17252 13176 17264
rect 12699 17224 13176 17252
rect 12699 17221 12711 17224
rect 12653 17215 12711 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 13265 17255 13323 17261
rect 13265 17221 13277 17255
rect 13311 17252 13323 17255
rect 13354 17252 13360 17264
rect 13311 17224 13360 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 13538 17261 13544 17264
rect 13481 17255 13544 17261
rect 13481 17221 13493 17255
rect 13527 17221 13544 17255
rect 13481 17215 13544 17221
rect 13538 17212 13544 17215
rect 13596 17252 13602 17264
rect 13814 17252 13820 17264
rect 13596 17224 13820 17252
rect 13596 17212 13602 17224
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 17129 17255 17187 17261
rect 17129 17252 17141 17255
rect 13964 17224 17141 17252
rect 13964 17212 13970 17224
rect 17129 17221 17141 17224
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 17310 17212 17316 17264
rect 17368 17252 17374 17264
rect 17368 17227 17402 17252
rect 17368 17221 17417 17227
rect 17368 17212 17371 17221
rect 8110 17184 8116 17196
rect 7852 17156 8116 17184
rect 7745 17147 7803 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 8444 17156 8585 17184
rect 8444 17144 8450 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 8938 17184 8944 17196
rect 8803 17156 8944 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 9180 17156 9597 17184
rect 9180 17144 9186 17156
rect 9585 17153 9597 17156
rect 9631 17184 9643 17187
rect 9766 17184 9772 17196
rect 9631 17156 9772 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 10152 17156 10333 17184
rect 5092 17088 5672 17116
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 10042 17116 10048 17128
rect 7055 17088 10048 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 5074 17048 5080 17060
rect 3952 17020 5080 17048
rect 5074 17008 5080 17020
rect 5132 17008 5138 17060
rect 5166 17008 5172 17060
rect 5224 17008 5230 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 5368 17020 6837 17048
rect 1636 16952 2912 16980
rect 1636 16940 1642 16952
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 5368 16980 5396 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 3384 16952 5396 16980
rect 3384 16940 3390 16952
rect 5810 16940 5816 16992
rect 5868 16980 5874 16992
rect 6730 16980 6736 16992
rect 5868 16952 6736 16980
rect 5868 16940 5874 16952
rect 6730 16940 6736 16952
rect 6788 16980 6794 16992
rect 6932 16980 6960 17079
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 7190 17008 7196 17060
rect 7248 17048 7254 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 7248 17020 7481 17048
rect 7248 17008 7254 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 6788 16952 6960 16980
rect 7484 16980 7512 17011
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 8941 17051 8999 17057
rect 8941 17048 8953 17051
rect 7708 17020 8953 17048
rect 7708 17008 7714 17020
rect 8941 17017 8953 17020
rect 8987 17017 8999 17051
rect 8941 17011 8999 17017
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 10152 17048 10180 17156
rect 10321 17153 10333 17156
rect 10367 17153 10379 17187
rect 10321 17147 10379 17153
rect 10980 17116 11008 17212
rect 11054 17144 11060 17196
rect 11112 17144 11118 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11480 17156 11713 17184
rect 11480 17144 11486 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14507 17156 15117 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 12250 17116 12256 17128
rect 10980 17088 12256 17116
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 12986 17076 12992 17128
rect 13044 17116 13050 17128
rect 13262 17116 13268 17128
rect 13044 17088 13268 17116
rect 13044 17076 13050 17088
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 9732 17020 10180 17048
rect 9732 17008 9738 17020
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 13814 17048 13820 17060
rect 10836 17020 12434 17048
rect 10836 17008 10842 17020
rect 8294 16980 8300 16992
rect 7484 16952 8300 16980
rect 6788 16940 6794 16952
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 10192 16952 11897 16980
rect 10192 16940 10198 16952
rect 11885 16949 11897 16952
rect 11931 16980 11943 16983
rect 12066 16980 12072 16992
rect 11931 16952 12072 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12406 16980 12434 17020
rect 12636 17020 13820 17048
rect 12636 16989 12664 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 14108 17048 14136 17147
rect 14292 17116 14320 17147
rect 16206 17144 16212 17196
rect 16264 17144 16270 17196
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17359 17187 17371 17212
rect 17405 17187 17417 17221
rect 18230 17212 18236 17264
rect 18288 17252 18294 17264
rect 18785 17255 18843 17261
rect 18785 17252 18797 17255
rect 18288 17224 18797 17252
rect 18288 17212 18294 17224
rect 18785 17221 18797 17224
rect 18831 17252 18843 17255
rect 19306 17252 19334 17292
rect 20088 17261 20116 17292
rect 20438 17280 20444 17332
rect 20496 17280 20502 17332
rect 21361 17323 21419 17329
rect 21361 17289 21373 17323
rect 21407 17320 21419 17323
rect 22278 17320 22284 17332
rect 21407 17292 22284 17320
rect 21407 17289 21419 17292
rect 21361 17283 21419 17289
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 26142 17320 26148 17332
rect 22480 17292 26148 17320
rect 18831 17224 19334 17252
rect 20073 17255 20131 17261
rect 18831 17221 18843 17224
rect 18785 17215 18843 17221
rect 20073 17221 20085 17255
rect 20119 17221 20131 17255
rect 20073 17215 20131 17221
rect 20165 17255 20223 17261
rect 20165 17221 20177 17255
rect 20211 17252 20223 17255
rect 22370 17252 22376 17264
rect 20211 17224 22376 17252
rect 20211 17221 20223 17224
rect 20165 17215 20223 17221
rect 22370 17212 22376 17224
rect 22428 17212 22434 17264
rect 18690 17193 18696 17196
rect 17359 17184 17417 17187
rect 17092 17181 17417 17184
rect 18509 17187 18567 17193
rect 17092 17156 17402 17181
rect 17092 17144 17098 17156
rect 18509 17153 18521 17187
rect 18555 17153 18567 17187
rect 18509 17147 18567 17153
rect 18657 17187 18696 17193
rect 18657 17153 18669 17187
rect 18657 17147 18696 17153
rect 14642 17116 14648 17128
rect 14292 17088 14648 17116
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 17586 17116 17592 17128
rect 16724 17088 17592 17116
rect 16724 17076 16730 17088
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 15470 17048 15476 17060
rect 14108 17020 15476 17048
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 18524 17048 18552 17147
rect 18690 17144 18696 17147
rect 18748 17144 18754 17196
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18782 17048 18788 17060
rect 17420 17020 18476 17048
rect 18524 17020 18788 17048
rect 12621 16983 12679 16989
rect 12621 16980 12633 16983
rect 12406 16952 12633 16980
rect 12621 16949 12633 16952
rect 12667 16949 12679 16983
rect 12621 16943 12679 16949
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12952 16952 13461 16980
rect 12952 16940 12958 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 13449 16943 13507 16949
rect 13630 16940 13636 16992
rect 13688 16940 13694 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 14734 16980 14740 16992
rect 14424 16952 14740 16980
rect 14424 16940 14430 16952
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 16025 16983 16083 16989
rect 16025 16949 16037 16983
rect 16071 16980 16083 16983
rect 16758 16980 16764 16992
rect 16071 16952 16764 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16980 17371 16983
rect 17420 16980 17448 17020
rect 17359 16952 17448 16980
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 18448 16980 18476 17020
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 18892 17048 18920 17147
rect 18966 17144 18972 17196
rect 19024 17193 19030 17196
rect 19978 17193 19984 17196
rect 19024 17184 19032 17193
rect 19797 17187 19855 17193
rect 19024 17156 19069 17184
rect 19024 17147 19032 17156
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 19945 17187 19984 17193
rect 19945 17153 19957 17187
rect 19945 17147 19984 17153
rect 19024 17144 19030 17147
rect 19812 17116 19840 17147
rect 19978 17144 19984 17147
rect 20036 17144 20042 17196
rect 20303 17187 20361 17193
rect 20303 17153 20315 17187
rect 20349 17184 20361 17187
rect 20714 17184 20720 17196
rect 20349 17156 20720 17184
rect 20349 17153 20361 17156
rect 20303 17147 20361 17153
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 21174 17144 21180 17196
rect 21232 17184 21238 17196
rect 22002 17184 22008 17196
rect 21232 17156 22008 17184
rect 21232 17144 21238 17156
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 20530 17116 20536 17128
rect 19812 17088 20536 17116
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 20901 17119 20959 17125
rect 20901 17085 20913 17119
rect 20947 17116 20959 17119
rect 21910 17116 21916 17128
rect 20947 17088 21916 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 21910 17076 21916 17088
rect 21968 17076 21974 17128
rect 22480 17116 22508 17292
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 26605 17323 26663 17329
rect 26605 17289 26617 17323
rect 26651 17289 26663 17323
rect 26605 17283 26663 17289
rect 22554 17212 22560 17264
rect 22612 17252 22618 17264
rect 26620 17252 26648 17283
rect 22612 17224 26648 17252
rect 22612 17212 22618 17224
rect 23106 17144 23112 17196
rect 23164 17184 23170 17196
rect 23457 17187 23515 17193
rect 23457 17184 23469 17187
rect 23164 17156 23469 17184
rect 23164 17144 23170 17156
rect 23457 17153 23469 17156
rect 23503 17153 23515 17187
rect 23457 17147 23515 17153
rect 25038 17144 25044 17196
rect 25096 17184 25102 17196
rect 25481 17187 25539 17193
rect 25481 17184 25493 17187
rect 25096 17156 25493 17184
rect 25096 17144 25102 17156
rect 25481 17153 25493 17156
rect 25527 17153 25539 17187
rect 25481 17147 25539 17153
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 26292 17156 27353 17184
rect 26292 17144 26298 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 22066 17088 22508 17116
rect 21177 17051 21235 17057
rect 21177 17048 21189 17051
rect 18892 17020 21189 17048
rect 21177 17017 21189 17020
rect 21223 17048 21235 17051
rect 22066 17048 22094 17088
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 23201 17119 23259 17125
rect 23201 17116 23213 17119
rect 22888 17088 23213 17116
rect 22888 17076 22894 17088
rect 23201 17085 23213 17088
rect 23247 17085 23259 17119
rect 23201 17079 23259 17085
rect 25225 17119 25283 17125
rect 25225 17085 25237 17119
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 21223 17020 22094 17048
rect 21223 17017 21235 17020
rect 21177 17011 21235 17017
rect 22370 17008 22376 17060
rect 22428 17008 22434 17060
rect 22462 17008 22468 17060
rect 22520 17008 22526 17060
rect 21082 16980 21088 16992
rect 18448 16952 21088 16980
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 23216 16980 23244 17079
rect 24578 17008 24584 17060
rect 24636 17008 24642 17060
rect 25240 16980 25268 17079
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 27672 17088 27905 17116
rect 27672 17076 27678 17088
rect 27893 17085 27905 17088
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 27798 17008 27804 17060
rect 27856 17048 27862 17060
rect 28169 17051 28227 17057
rect 28169 17048 28181 17051
rect 27856 17020 28181 17048
rect 27856 17008 27862 17020
rect 28169 17017 28181 17020
rect 28215 17017 28227 17051
rect 28169 17011 28227 17017
rect 26786 16980 26792 16992
rect 23216 16952 26792 16980
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27157 16983 27215 16989
rect 27157 16980 27169 16983
rect 27120 16952 27169 16980
rect 27120 16940 27126 16952
rect 27157 16949 27169 16952
rect 27203 16949 27215 16983
rect 27157 16943 27215 16949
rect 27522 16940 27528 16992
rect 27580 16980 27586 16992
rect 28353 16983 28411 16989
rect 28353 16980 28365 16983
rect 27580 16952 28365 16980
rect 27580 16940 27586 16952
rect 28353 16949 28365 16952
rect 28399 16949 28411 16983
rect 28353 16943 28411 16949
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 1762 16736 1768 16788
rect 1820 16736 1826 16788
rect 5169 16779 5227 16785
rect 5169 16745 5181 16779
rect 5215 16776 5227 16779
rect 5350 16776 5356 16788
rect 5215 16748 5356 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5592 16748 5641 16776
rect 5592 16736 5598 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 5629 16739 5687 16745
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7190 16776 7196 16788
rect 7064 16748 7196 16776
rect 7064 16736 7070 16748
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7558 16736 7564 16788
rect 7616 16736 7622 16788
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 12710 16776 12716 16788
rect 10376 16748 12716 16776
rect 10376 16736 10382 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13541 16779 13599 16785
rect 13541 16745 13553 16779
rect 13587 16776 13599 16779
rect 13998 16776 14004 16788
rect 13587 16748 14004 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 15470 16776 15476 16788
rect 14240 16748 15476 16776
rect 14240 16736 14246 16748
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 15930 16736 15936 16788
rect 15988 16776 15994 16788
rect 16942 16776 16948 16788
rect 15988 16748 16948 16776
rect 15988 16736 15994 16748
rect 16942 16736 16948 16748
rect 17000 16776 17006 16788
rect 17770 16776 17776 16788
rect 17000 16748 17776 16776
rect 17000 16736 17006 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 20809 16779 20867 16785
rect 20809 16776 20821 16779
rect 18840 16748 20821 16776
rect 18840 16736 18846 16748
rect 20809 16745 20821 16748
rect 20855 16745 20867 16779
rect 25682 16776 25688 16788
rect 20809 16739 20867 16745
rect 23400 16748 25688 16776
rect 1946 16668 1952 16720
rect 2004 16708 2010 16720
rect 2774 16708 2780 16720
rect 2004 16680 2780 16708
rect 2004 16668 2010 16680
rect 2774 16668 2780 16680
rect 2832 16708 2838 16720
rect 5077 16711 5135 16717
rect 5077 16708 5089 16711
rect 2832 16680 5089 16708
rect 2832 16668 2838 16680
rect 5077 16677 5089 16680
rect 5123 16708 5135 16711
rect 5258 16708 5264 16720
rect 5123 16680 5264 16708
rect 5123 16677 5135 16680
rect 5077 16671 5135 16677
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 8294 16668 8300 16720
rect 8352 16668 8358 16720
rect 11974 16708 11980 16720
rect 9324 16680 11980 16708
rect 6546 16640 6552 16652
rect 5368 16612 6552 16640
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 1949 16575 2007 16581
rect 1949 16572 1961 16575
rect 1636 16544 1961 16572
rect 1636 16532 1642 16544
rect 1949 16541 1961 16544
rect 1995 16541 2007 16575
rect 1949 16535 2007 16541
rect 2222 16532 2228 16584
rect 2280 16532 2286 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3142 16572 3148 16584
rect 3099 16544 3148 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3786 16572 3792 16584
rect 3467 16544 3792 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4249 16575 4307 16581
rect 4111 16544 4200 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 4172 16516 4200 16544
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 5368 16572 5396 16612
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6638 16600 6644 16652
rect 6696 16600 6702 16652
rect 6730 16600 6736 16652
rect 6788 16640 6794 16652
rect 8312 16640 8340 16668
rect 6788 16612 7880 16640
rect 8312 16612 8432 16640
rect 6788 16600 6794 16612
rect 4295 16544 5396 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 5810 16532 5816 16584
rect 5868 16532 5874 16584
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6825 16575 6883 16581
rect 6825 16572 6837 16575
rect 6420 16544 6837 16572
rect 6420 16532 6426 16544
rect 6825 16541 6837 16544
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7650 16572 7656 16584
rect 7147 16544 7656 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7852 16581 7880 16612
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 7926 16532 7932 16584
rect 7984 16572 7990 16584
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 7984 16544 8309 16572
rect 7984 16532 7990 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8404 16572 8432 16612
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9324 16649 9352 16680
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 12986 16708 12992 16720
rect 12216 16680 12992 16708
rect 12216 16668 12222 16680
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 15436 16680 18460 16708
rect 15436 16668 15442 16680
rect 9309 16643 9367 16649
rect 8904 16612 9260 16640
rect 8904 16600 8910 16612
rect 9122 16572 9128 16584
rect 8404 16544 9128 16572
rect 8297 16535 8355 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9232 16572 9260 16612
rect 9309 16609 9321 16643
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10744 16612 10793 16640
rect 10744 16600 10750 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16640 11023 16643
rect 11011 16612 14412 16640
rect 11011 16609 11023 16612
rect 10965 16603 11023 16609
rect 9674 16572 9680 16584
rect 9232 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 11333 16575 11391 16581
rect 9784 16544 10732 16572
rect 2133 16507 2191 16513
rect 2133 16473 2145 16507
rect 2179 16504 2191 16507
rect 2498 16504 2504 16516
rect 2179 16476 2504 16504
rect 2179 16473 2191 16476
rect 2133 16467 2191 16473
rect 2498 16464 2504 16476
rect 2556 16464 2562 16516
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 4154 16504 4160 16516
rect 2648 16476 4160 16504
rect 2648 16464 2654 16476
rect 4154 16464 4160 16476
rect 4212 16504 4218 16516
rect 4212 16476 4660 16504
rect 4212 16464 4218 16476
rect 4246 16396 4252 16448
rect 4304 16396 4310 16448
rect 4632 16436 4660 16476
rect 4706 16464 4712 16516
rect 4764 16464 4770 16516
rect 5997 16507 6055 16513
rect 5997 16473 6009 16507
rect 6043 16504 6055 16507
rect 6043 16476 7512 16504
rect 6043 16473 6055 16476
rect 5997 16467 6055 16473
rect 5166 16436 5172 16448
rect 4632 16408 5172 16436
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 5718 16396 5724 16448
rect 5776 16436 5782 16448
rect 6454 16436 6460 16448
rect 5776 16408 6460 16436
rect 5776 16396 5782 16408
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 7006 16396 7012 16448
rect 7064 16396 7070 16448
rect 7484 16436 7512 16476
rect 7558 16464 7564 16516
rect 7616 16464 7622 16516
rect 7742 16464 7748 16516
rect 7800 16464 7806 16516
rect 9784 16504 9812 16544
rect 8404 16476 9812 16504
rect 9861 16507 9919 16513
rect 8404 16436 8432 16476
rect 9861 16473 9873 16507
rect 9907 16504 9919 16507
rect 9950 16504 9956 16516
rect 9907 16476 9956 16504
rect 9907 16473 9919 16476
rect 9861 16467 9919 16473
rect 9950 16464 9956 16476
rect 10008 16504 10014 16516
rect 10226 16504 10232 16516
rect 10008 16476 10232 16504
rect 10008 16464 10014 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10704 16504 10732 16544
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 11379 16544 12081 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 12069 16541 12081 16544
rect 12115 16572 12127 16575
rect 12342 16572 12348 16584
rect 12115 16544 12348 16572
rect 12115 16541 12127 16544
rect 12069 16535 12127 16541
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 12492 16544 12633 16572
rect 12492 16532 12498 16544
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 13136 16544 14289 16572
rect 13136 16532 13142 16544
rect 14277 16541 14289 16544
rect 14323 16541 14335 16575
rect 14384 16572 14412 16612
rect 16040 16612 16903 16640
rect 16040 16572 16068 16612
rect 14384 16544 16068 16572
rect 14277 16535 14335 16541
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 16390 16532 16396 16584
rect 16448 16532 16454 16584
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16572 16543 16575
rect 16666 16572 16672 16584
rect 16531 16544 16672 16572
rect 16531 16541 16543 16544
rect 16485 16535 16543 16541
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16875 16572 16903 16612
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 17000 16612 17141 16640
rect 17000 16600 17006 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17497 16643 17555 16649
rect 17129 16603 17187 16609
rect 17236 16612 17448 16640
rect 17236 16572 17264 16612
rect 16875 16544 17264 16572
rect 17310 16532 17316 16584
rect 17368 16532 17374 16584
rect 17420 16572 17448 16612
rect 17497 16609 17509 16643
rect 17543 16640 17555 16643
rect 17586 16640 17592 16652
rect 17543 16612 17592 16640
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17828 16612 17969 16640
rect 17828 16600 17834 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 18046 16600 18052 16652
rect 18104 16640 18110 16652
rect 18325 16643 18383 16649
rect 18325 16640 18337 16643
rect 18104 16612 18337 16640
rect 18104 16600 18110 16612
rect 18325 16609 18337 16612
rect 18371 16609 18383 16643
rect 18432 16640 18460 16680
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19797 16711 19855 16717
rect 19797 16708 19809 16711
rect 19024 16680 19809 16708
rect 19024 16668 19030 16680
rect 19797 16677 19809 16680
rect 19843 16708 19855 16711
rect 20714 16708 20720 16720
rect 19843 16680 20720 16708
rect 19843 16677 19855 16680
rect 19797 16671 19855 16677
rect 20714 16668 20720 16680
rect 20772 16668 20778 16720
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 23400 16708 23428 16748
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 26786 16776 26792 16788
rect 26620 16748 26792 16776
rect 22336 16680 23428 16708
rect 23569 16711 23627 16717
rect 22336 16668 22342 16680
rect 23569 16677 23581 16711
rect 23615 16708 23627 16711
rect 23842 16708 23848 16720
rect 23615 16680 23848 16708
rect 23615 16677 23627 16680
rect 23569 16671 23627 16677
rect 18432 16612 19196 16640
rect 18325 16603 18383 16609
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 17420 16544 18153 16572
rect 18141 16541 18153 16544
rect 18187 16572 18199 16575
rect 18690 16572 18696 16584
rect 18187 16544 18696 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 11054 16504 11060 16516
rect 10704 16476 11060 16504
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 11422 16464 11428 16516
rect 11480 16464 11486 16516
rect 11514 16464 11520 16516
rect 11572 16464 11578 16516
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12253 16507 12311 16513
rect 12253 16504 12265 16507
rect 12216 16476 12265 16504
rect 12216 16464 12222 16476
rect 12253 16473 12265 16476
rect 12299 16473 12311 16507
rect 12253 16467 12311 16473
rect 12805 16507 12863 16513
rect 12805 16473 12817 16507
rect 12851 16473 12863 16507
rect 12805 16467 12863 16473
rect 7484 16408 8432 16436
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16436 8539 16439
rect 9398 16436 9404 16448
rect 8527 16408 9404 16436
rect 8527 16405 8539 16408
rect 8481 16399 8539 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 9769 16439 9827 16445
rect 9769 16405 9781 16439
rect 9815 16436 9827 16439
rect 10042 16436 10048 16448
rect 9815 16408 10048 16436
rect 9815 16405 9827 16408
rect 9769 16399 9827 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 12820 16436 12848 16467
rect 13354 16464 13360 16516
rect 13412 16464 13418 16516
rect 14522 16507 14580 16513
rect 14522 16504 14534 16507
rect 13464 16476 14534 16504
rect 10744 16408 12848 16436
rect 10744 16396 10750 16408
rect 12986 16396 12992 16448
rect 13044 16436 13050 16448
rect 13464 16436 13492 16476
rect 14522 16473 14534 16476
rect 14568 16473 14580 16507
rect 14522 16467 14580 16473
rect 16301 16507 16359 16513
rect 16301 16473 16313 16507
rect 16347 16504 16359 16507
rect 17862 16504 17868 16516
rect 16347 16476 17868 16504
rect 16347 16473 16359 16476
rect 16301 16467 16359 16473
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 19168 16504 19196 16612
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19429 16643 19487 16649
rect 19300 16612 19380 16640
rect 19300 16600 19306 16612
rect 19352 16572 19380 16612
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19886 16640 19892 16652
rect 19475 16612 19892 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19886 16600 19892 16612
rect 19944 16600 19950 16652
rect 21174 16640 21180 16652
rect 20732 16612 21180 16640
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 19352 16544 19625 16572
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 20732 16504 20760 16612
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21453 16643 21511 16649
rect 21453 16609 21465 16643
rect 21499 16640 21511 16643
rect 23584 16640 23612 16671
rect 23842 16668 23848 16680
rect 23900 16668 23906 16720
rect 26145 16711 26203 16717
rect 26145 16677 26157 16711
rect 26191 16677 26203 16711
rect 26145 16671 26203 16677
rect 21499 16612 23612 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 24765 16643 24823 16649
rect 24765 16640 24777 16643
rect 24636 16612 24777 16640
rect 24636 16600 24642 16612
rect 24765 16609 24777 16612
rect 24811 16609 24823 16643
rect 24765 16603 24823 16609
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20956 16544 21005 16572
rect 20956 16532 20962 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16572 21143 16575
rect 23382 16572 23388 16584
rect 21131 16544 23388 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 23382 16532 23388 16544
rect 23440 16572 23446 16584
rect 26160 16572 26188 16671
rect 26620 16649 26648 16748
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 26605 16643 26663 16649
rect 26605 16609 26617 16643
rect 26651 16609 26663 16643
rect 26605 16603 26663 16609
rect 23440 16544 26188 16572
rect 23440 16532 23446 16544
rect 19168 16476 20760 16504
rect 21174 16464 21180 16516
rect 21232 16464 21238 16516
rect 21295 16507 21353 16513
rect 21295 16473 21307 16507
rect 21341 16473 21353 16507
rect 21295 16467 21353 16473
rect 13044 16408 13492 16436
rect 13044 16396 13050 16408
rect 13538 16396 13544 16448
rect 13596 16445 13602 16448
rect 13596 16439 13615 16445
rect 13603 16405 13615 16439
rect 13596 16399 13615 16405
rect 13596 16396 13602 16399
rect 13722 16396 13728 16448
rect 13780 16396 13786 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 15657 16439 15715 16445
rect 15657 16436 15669 16439
rect 13872 16408 15669 16436
rect 13872 16396 13878 16408
rect 15657 16405 15669 16408
rect 15703 16405 15715 16439
rect 15657 16399 15715 16405
rect 16666 16396 16672 16448
rect 16724 16396 16730 16448
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 20346 16436 20352 16448
rect 17000 16408 20352 16436
rect 17000 16396 17006 16408
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 20990 16436 20996 16448
rect 20496 16408 20996 16436
rect 20496 16396 20502 16408
rect 20990 16396 20996 16408
rect 21048 16436 21054 16448
rect 21310 16436 21338 16467
rect 21634 16464 21640 16516
rect 21692 16504 21698 16516
rect 21910 16504 21916 16516
rect 21692 16476 21916 16504
rect 21692 16464 21698 16476
rect 21910 16464 21916 16476
rect 21968 16464 21974 16516
rect 22002 16464 22008 16516
rect 22060 16504 22066 16516
rect 23201 16507 23259 16513
rect 23201 16504 23213 16507
rect 22060 16476 23213 16504
rect 22060 16464 22066 16476
rect 23201 16473 23213 16476
rect 23247 16504 23259 16507
rect 23290 16504 23296 16516
rect 23247 16476 23296 16504
rect 23247 16473 23259 16476
rect 23201 16467 23259 16473
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 24854 16464 24860 16516
rect 24912 16504 24918 16516
rect 25010 16507 25068 16513
rect 25010 16504 25022 16507
rect 24912 16476 25022 16504
rect 24912 16464 24918 16476
rect 25010 16473 25022 16476
rect 25056 16473 25068 16507
rect 25010 16467 25068 16473
rect 26050 16464 26056 16516
rect 26108 16504 26114 16516
rect 26850 16507 26908 16513
rect 26850 16504 26862 16507
rect 26108 16476 26862 16504
rect 26108 16464 26114 16476
rect 26850 16473 26862 16476
rect 26896 16473 26908 16507
rect 26850 16467 26908 16473
rect 21048 16408 21338 16436
rect 22373 16439 22431 16445
rect 21048 16396 21054 16408
rect 22373 16405 22385 16439
rect 22419 16436 22431 16439
rect 23474 16436 23480 16448
rect 22419 16408 23480 16436
rect 22419 16405 22431 16408
rect 22373 16399 22431 16405
rect 23474 16396 23480 16408
rect 23532 16396 23538 16448
rect 23661 16439 23719 16445
rect 23661 16405 23673 16439
rect 23707 16436 23719 16439
rect 24026 16436 24032 16448
rect 23707 16408 24032 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 24026 16396 24032 16408
rect 24084 16396 24090 16448
rect 24118 16396 24124 16448
rect 24176 16436 24182 16448
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 24176 16408 27997 16436
rect 24176 16396 24182 16408
rect 27985 16405 27997 16408
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 1857 16235 1915 16241
rect 1857 16201 1869 16235
rect 1903 16232 1915 16235
rect 3786 16232 3792 16244
rect 1903 16204 3792 16232
rect 1903 16201 1915 16204
rect 1857 16195 1915 16201
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 3878 16192 3884 16244
rect 3936 16192 3942 16244
rect 5997 16235 6055 16241
rect 5997 16201 6009 16235
rect 6043 16232 6055 16235
rect 7006 16232 7012 16244
rect 6043 16204 7012 16232
rect 6043 16201 6055 16204
rect 5997 16195 6055 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 8846 16192 8852 16244
rect 8904 16192 8910 16244
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 10226 16232 10232 16244
rect 8987 16204 10232 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 10410 16192 10416 16244
rect 10468 16192 10474 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 10928 16204 10977 16232
rect 10928 16192 10934 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11974 16232 11980 16244
rect 11112 16204 11980 16232
rect 11112 16192 11118 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 14642 16232 14648 16244
rect 12768 16204 14648 16232
rect 12768 16192 12774 16204
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 15565 16235 15623 16241
rect 15565 16232 15577 16235
rect 14976 16204 15577 16232
rect 14976 16192 14982 16204
rect 15565 16201 15577 16204
rect 15611 16201 15623 16235
rect 18049 16235 18107 16241
rect 15565 16195 15623 16201
rect 15948 16204 17540 16232
rect 4985 16167 5043 16173
rect 4985 16133 4997 16167
rect 5031 16164 5043 16167
rect 5350 16164 5356 16176
rect 5031 16136 5356 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 5350 16124 5356 16136
rect 5408 16124 5414 16176
rect 6270 16164 6276 16176
rect 5828 16136 6276 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1762 16096 1768 16108
rect 1719 16068 1768 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 2498 16096 2504 16108
rect 1995 16068 2504 16096
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2590 16056 2596 16108
rect 2648 16056 2654 16108
rect 4062 16056 4068 16108
rect 4120 16096 4126 16108
rect 4706 16096 4712 16108
rect 4120 16068 4712 16096
rect 4120 16056 4126 16068
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4764 16068 4813 16096
rect 4764 16056 4770 16068
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5258 16096 5264 16108
rect 5123 16068 5264 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5828 16105 5856 16136
rect 6270 16124 6276 16136
rect 6328 16124 6334 16176
rect 6454 16124 6460 16176
rect 6512 16164 6518 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 6512 16136 6561 16164
rect 6512 16124 6518 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 6749 16167 6807 16173
rect 6749 16164 6761 16167
rect 6549 16127 6607 16133
rect 6748 16133 6761 16164
rect 6795 16164 6807 16167
rect 8386 16164 8392 16176
rect 6795 16136 8392 16164
rect 6795 16133 6807 16136
rect 6748 16127 6807 16133
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5994 16056 6000 16108
rect 6052 16096 6058 16108
rect 6288 16096 6316 16124
rect 6748 16096 6776 16127
rect 8386 16124 8392 16136
rect 8444 16124 8450 16176
rect 8956 16136 13216 16164
rect 6052 16068 6132 16096
rect 6288 16068 6776 16096
rect 6052 16056 6058 16068
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 2188 16000 6040 16028
rect 2188 15988 2194 16000
rect 6012 15972 6040 16000
rect 5994 15920 6000 15972
rect 6052 15920 6058 15972
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 3050 15892 3056 15904
rect 1719 15864 3056 15892
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 4801 15895 4859 15901
rect 4801 15861 4813 15895
rect 4847 15892 4859 15895
rect 5534 15892 5540 15904
rect 4847 15864 5540 15892
rect 4847 15861 4859 15864
rect 4801 15855 4859 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 6104 15892 6132 16068
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7282 16096 7288 16108
rect 7156 16068 7288 16096
rect 7156 16056 7162 16068
rect 7282 16056 7288 16068
rect 7340 16096 7346 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7340 16068 7389 16096
rect 7340 16056 7346 16068
rect 7377 16065 7389 16068
rect 7423 16096 7435 16099
rect 7423 16068 7788 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 7558 15988 7564 16040
rect 7616 15988 7622 16040
rect 7760 16028 7788 16068
rect 8294 16056 8300 16108
rect 8352 16056 8358 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8956 16096 8984 16136
rect 13188 16108 13216 16136
rect 13262 16124 13268 16176
rect 13320 16164 13326 16176
rect 13541 16167 13599 16173
rect 13541 16164 13553 16167
rect 13320 16136 13553 16164
rect 13320 16124 13326 16136
rect 13541 16133 13553 16136
rect 13587 16133 13599 16167
rect 13541 16127 13599 16133
rect 13771 16133 13829 16139
rect 13771 16130 13783 16133
rect 8527 16068 8984 16096
rect 9033 16099 9091 16105
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9122 16096 9128 16108
rect 9079 16068 9128 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9122 16056 9128 16068
rect 9180 16096 9186 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9180 16068 9965 16096
rect 9180 16056 9186 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10502 16096 10508 16108
rect 10275 16068 10508 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 10928 16068 11161 16096
rect 10928 16056 10934 16068
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11296 16068 11713 16096
rect 11296 16056 11302 16068
rect 11701 16065 11713 16068
rect 11747 16096 11759 16099
rect 12526 16096 12532 16108
rect 11747 16068 12532 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 10042 16028 10048 16040
rect 7760 16000 10048 16028
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10686 16028 10692 16040
rect 10183 16000 10692 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 12636 16028 12664 16059
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12894 16056 12900 16108
rect 12952 16056 12958 16108
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 12802 16028 12808 16040
rect 12636 16000 12808 16028
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 13004 16028 13032 16059
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13761 16099 13783 16130
rect 13817 16099 13829 16133
rect 14458 16124 14464 16176
rect 14516 16164 14522 16176
rect 15948 16164 15976 16204
rect 17405 16167 17463 16173
rect 17405 16164 17417 16167
rect 14516 16136 15976 16164
rect 16040 16136 17417 16164
rect 14516 16124 14522 16136
rect 13761 16096 13829 16099
rect 15194 16096 15200 16108
rect 13228 16068 15200 16096
rect 13228 16056 13234 16068
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15562 16056 15568 16108
rect 15620 16056 15626 16108
rect 15746 16056 15752 16108
rect 15804 16056 15810 16108
rect 16040 16105 16068 16136
rect 17405 16133 17417 16136
rect 17451 16133 17463 16167
rect 17512 16164 17540 16204
rect 18049 16201 18061 16235
rect 18095 16232 18107 16235
rect 19058 16232 19064 16244
rect 18095 16204 19064 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 19334 16192 19340 16244
rect 19392 16192 19398 16244
rect 20533 16235 20591 16241
rect 20533 16232 20545 16235
rect 19444 16204 20545 16232
rect 19444 16164 19472 16204
rect 20533 16201 20545 16204
rect 20579 16201 20591 16235
rect 20533 16195 20591 16201
rect 21177 16235 21235 16241
rect 21177 16201 21189 16235
rect 21223 16232 21235 16235
rect 22278 16232 22284 16244
rect 21223 16204 22284 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 23753 16235 23811 16241
rect 23753 16201 23765 16235
rect 23799 16232 23811 16235
rect 26234 16232 26240 16244
rect 23799 16204 26240 16232
rect 23799 16201 23811 16204
rect 23753 16195 23811 16201
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 27341 16235 27399 16241
rect 27341 16201 27353 16235
rect 27387 16201 27399 16235
rect 27341 16195 27399 16201
rect 17512 16136 19472 16164
rect 19935 16167 19993 16173
rect 17405 16127 17463 16133
rect 19935 16133 19947 16167
rect 19981 16164 19993 16167
rect 22370 16164 22376 16176
rect 19981 16136 22376 16164
rect 19981 16133 19993 16136
rect 19935 16127 19993 16133
rect 22370 16124 22376 16136
rect 22428 16164 22434 16176
rect 22428 16136 22784 16164
rect 22428 16124 22434 16136
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16206 16056 16212 16108
rect 16264 16056 16270 16108
rect 17494 16056 17500 16108
rect 17552 16096 17558 16108
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 17552 16068 17785 16096
rect 17552 16056 17558 16068
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17920 16068 18153 16096
rect 17920 16056 17926 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 18656 16068 18705 16096
rect 18656 16056 18662 16068
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16096 18935 16099
rect 19426 16096 19432 16108
rect 18923 16068 19432 16096
rect 18923 16065 18935 16068
rect 18877 16059 18935 16065
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 20073 16099 20131 16105
rect 20073 16096 20085 16099
rect 19536 16068 20085 16096
rect 17678 16028 17684 16040
rect 13004 16000 17684 16028
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 19536 16028 19564 16068
rect 20073 16065 20085 16068
rect 20119 16096 20131 16099
rect 20438 16096 20444 16108
rect 20119 16068 20444 16096
rect 20119 16065 20131 16068
rect 20073 16059 20131 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20772 16068 21281 16096
rect 20772 16056 20778 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 22646 16096 22652 16108
rect 21269 16059 21327 16065
rect 21468 16068 22652 16096
rect 19306 16000 19564 16028
rect 19797 16031 19855 16037
rect 8202 15960 8208 15972
rect 6748 15932 8208 15960
rect 6748 15901 6776 15932
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 8938 15960 8944 15972
rect 8260 15932 8944 15960
rect 8260 15920 8266 15932
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13262 15960 13268 15972
rect 12676 15932 13268 15960
rect 12676 15920 12682 15932
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 17218 15920 17224 15972
rect 17276 15960 17282 15972
rect 19306 15960 19334 16000
rect 19797 15997 19809 16031
rect 19843 16028 19855 16031
rect 20622 16028 20628 16040
rect 19843 16000 20628 16028
rect 19843 15997 19855 16000
rect 19797 15991 19855 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 16028 20867 16031
rect 21468 16028 21496 16068
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 22756 16096 22784 16136
rect 23290 16124 23296 16176
rect 23348 16124 23354 16176
rect 24480 16167 24538 16173
rect 24480 16133 24492 16167
rect 24526 16164 24538 16167
rect 27356 16164 27384 16195
rect 27430 16192 27436 16244
rect 27488 16232 27494 16244
rect 27985 16235 28043 16241
rect 27985 16232 27997 16235
rect 27488 16204 27997 16232
rect 27488 16192 27494 16204
rect 27985 16201 27997 16204
rect 28031 16201 28043 16235
rect 27985 16195 28043 16201
rect 24526 16136 27384 16164
rect 24526 16133 24538 16136
rect 24480 16127 24538 16133
rect 25590 16096 25596 16108
rect 22756 16068 25596 16096
rect 25590 16056 25596 16068
rect 25648 16056 25654 16108
rect 27522 16056 27528 16108
rect 27580 16056 27586 16108
rect 28166 16056 28172 16108
rect 28224 16056 28230 16108
rect 20855 16000 21496 16028
rect 22005 16031 22063 16037
rect 20855 15997 20867 16000
rect 20809 15991 20867 15997
rect 22005 15997 22017 16031
rect 22051 16028 22063 16031
rect 22554 16028 22560 16040
rect 22051 16000 22560 16028
rect 22051 15997 22063 16000
rect 22005 15991 22063 15997
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 24026 15988 24032 16040
rect 24084 16028 24090 16040
rect 24213 16031 24271 16037
rect 24213 16028 24225 16031
rect 24084 16000 24225 16028
rect 24084 15988 24090 16000
rect 24213 15997 24225 16000
rect 24259 15997 24271 16031
rect 24213 15991 24271 15997
rect 17276 15932 19334 15960
rect 17276 15920 17282 15932
rect 19426 15920 19432 15972
rect 19484 15960 19490 15972
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 19484 15932 19717 15960
rect 19484 15920 19490 15932
rect 19705 15929 19717 15932
rect 19751 15929 19763 15963
rect 19705 15923 19763 15929
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 22373 15963 22431 15969
rect 22373 15960 22385 15963
rect 20404 15932 22385 15960
rect 20404 15920 20410 15932
rect 22373 15929 22385 15932
rect 22419 15960 22431 15963
rect 23566 15960 23572 15972
rect 22419 15932 23572 15960
rect 22419 15929 22431 15932
rect 22373 15923 22431 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 23658 15920 23664 15972
rect 23716 15960 23722 15972
rect 24118 15960 24124 15972
rect 23716 15932 24124 15960
rect 23716 15920 23722 15932
rect 24118 15920 24124 15932
rect 24176 15920 24182 15972
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 5684 15864 6745 15892
rect 5684 15852 5690 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 6733 15855 6791 15861
rect 6914 15852 6920 15904
rect 6972 15852 6978 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 9490 15892 9496 15904
rect 8352 15864 9496 15892
rect 8352 15852 8358 15864
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15892 10287 15895
rect 10318 15892 10324 15904
rect 10275 15864 10324 15892
rect 10275 15861 10287 15864
rect 10229 15855 10287 15861
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11885 15895 11943 15901
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 12066 15892 12072 15904
rect 11931 15864 12072 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12434 15852 12440 15904
rect 12492 15852 12498 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13596 15864 13737 15892
rect 13596 15852 13602 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 13909 15895 13967 15901
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 14642 15892 14648 15904
rect 13955 15864 14648 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 17678 15852 17684 15904
rect 17736 15852 17742 15904
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17828 15864 17877 15892
rect 17828 15852 17834 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 20438 15892 20444 15904
rect 19659 15864 20444 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 20993 15895 21051 15901
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 21818 15892 21824 15904
rect 21039 15864 21824 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 22465 15895 22523 15901
rect 22465 15861 22477 15895
rect 22511 15892 22523 15895
rect 23290 15892 23296 15904
rect 22511 15864 23296 15892
rect 22511 15861 22523 15864
rect 22465 15855 22523 15861
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 25593 15895 25651 15901
rect 25593 15861 25605 15895
rect 25639 15892 25651 15895
rect 27706 15892 27712 15904
rect 25639 15864 27712 15892
rect 25639 15861 25651 15864
rect 25593 15855 25651 15861
rect 27706 15852 27712 15864
rect 27764 15852 27770 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1210 15648 1216 15700
rect 1268 15688 1274 15700
rect 2130 15688 2136 15700
rect 1268 15660 2136 15688
rect 1268 15648 1274 15660
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2222 15648 2228 15700
rect 2280 15688 2286 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2280 15660 2513 15688
rect 2280 15648 2286 15660
rect 2501 15657 2513 15660
rect 2547 15688 2559 15691
rect 4062 15688 4068 15700
rect 2547 15660 4068 15688
rect 2547 15657 2559 15660
rect 2501 15651 2559 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 5077 15691 5135 15697
rect 5077 15657 5089 15691
rect 5123 15688 5135 15691
rect 6086 15688 6092 15700
rect 5123 15660 6092 15688
rect 5123 15657 5135 15660
rect 5077 15651 5135 15657
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 14918 15688 14924 15700
rect 8536 15660 14924 15688
rect 8536 15648 8542 15660
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 17037 15691 17095 15697
rect 16080 15660 16903 15688
rect 16080 15648 16086 15660
rect 3234 15580 3240 15632
rect 3292 15620 3298 15632
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 3292 15592 4353 15620
rect 3292 15580 3298 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 4798 15580 4804 15632
rect 4856 15620 4862 15632
rect 5629 15623 5687 15629
rect 5629 15620 5641 15623
rect 4856 15592 5641 15620
rect 4856 15580 4862 15592
rect 5629 15589 5641 15592
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 8113 15623 8171 15629
rect 8113 15620 8125 15623
rect 7432 15592 8125 15620
rect 7432 15580 7438 15592
rect 8113 15589 8125 15592
rect 8159 15589 8171 15623
rect 8113 15583 8171 15589
rect 8294 15580 8300 15632
rect 8352 15580 8358 15632
rect 14458 15580 14464 15632
rect 14516 15620 14522 15632
rect 14553 15623 14611 15629
rect 14553 15620 14565 15623
rect 14516 15592 14565 15620
rect 14516 15580 14522 15592
rect 14553 15589 14565 15592
rect 14599 15589 14611 15623
rect 14553 15583 14611 15589
rect 14645 15623 14703 15629
rect 14645 15589 14657 15623
rect 14691 15620 14703 15623
rect 16482 15620 16488 15632
rect 14691 15592 16488 15620
rect 14691 15589 14703 15592
rect 14645 15583 14703 15589
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 16875 15620 16903 15660
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 17494 15688 17500 15700
rect 17083 15660 17500 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 17494 15648 17500 15660
rect 17552 15688 17558 15700
rect 17862 15688 17868 15700
rect 17552 15660 17868 15688
rect 17552 15648 17558 15660
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18601 15691 18659 15697
rect 18601 15657 18613 15691
rect 18647 15688 18659 15691
rect 20346 15688 20352 15700
rect 18647 15660 20352 15688
rect 18647 15657 18659 15660
rect 18601 15651 18659 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20441 15691 20499 15697
rect 20441 15657 20453 15691
rect 20487 15688 20499 15691
rect 20487 15660 21128 15688
rect 20487 15657 20499 15660
rect 20441 15651 20499 15657
rect 16875 15592 16988 15620
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 3510 15552 3516 15564
rect 2832 15524 3516 15552
rect 2832 15512 2838 15524
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15552 4307 15555
rect 4295 15524 5580 15552
rect 4295 15521 4307 15524
rect 4249 15515 4307 15521
rect 5552 15496 5580 15524
rect 5718 15512 5724 15564
rect 5776 15552 5782 15564
rect 6825 15555 6883 15561
rect 5776 15524 5948 15552
rect 5776 15512 5782 15524
rect 474 15444 480 15496
rect 532 15484 538 15496
rect 1673 15487 1731 15493
rect 1673 15484 1685 15487
rect 532 15456 1685 15484
rect 532 15444 538 15456
rect 1673 15453 1685 15456
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 1903 15456 2636 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 2608 15416 2636 15456
rect 2682 15444 2688 15496
rect 2740 15444 2746 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4430 15444 4436 15496
rect 4488 15444 4494 15496
rect 4982 15444 4988 15496
rect 5040 15493 5046 15496
rect 5040 15484 5049 15493
rect 5169 15487 5227 15493
rect 5040 15456 5085 15484
rect 5040 15447 5049 15456
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5258 15484 5264 15496
rect 5215 15456 5264 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5040 15444 5046 15447
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 5920 15493 5948 15524
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 8312 15552 8340 15580
rect 6871 15524 8340 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 9950 15512 9956 15564
rect 10008 15512 10014 15564
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 10962 15552 10968 15564
rect 10468 15524 10968 15552
rect 10468 15512 10474 15524
rect 10962 15512 10968 15524
rect 11020 15552 11026 15564
rect 11020 15524 11284 15552
rect 11020 15512 11026 15524
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5592 15456 5825 15484
rect 5592 15444 5598 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 5994 15444 6000 15496
rect 6052 15484 6058 15496
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 6052 15456 6101 15484
rect 6052 15444 6058 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15453 6239 15487
rect 6181 15447 6239 15453
rect 7101 15487 7159 15493
rect 7101 15453 7113 15487
rect 7147 15484 7159 15487
rect 8294 15484 8300 15496
rect 7147 15456 8300 15484
rect 7147 15453 7159 15456
rect 7101 15447 7159 15453
rect 2774 15416 2780 15428
rect 2608 15388 2780 15416
rect 2774 15376 2780 15388
rect 2832 15376 2838 15428
rect 2961 15419 3019 15425
rect 2961 15385 2973 15419
rect 3007 15416 3019 15419
rect 3234 15416 3240 15428
rect 3007 15388 3240 15416
rect 3007 15385 3019 15388
rect 2961 15379 3019 15385
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 4798 15376 4804 15428
rect 4856 15416 4862 15428
rect 6196 15416 6224 15447
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8570 15484 8576 15496
rect 8435 15456 8576 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9732 15456 9781 15484
rect 9732 15444 9738 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 11146 15444 11152 15496
rect 11204 15444 11210 15496
rect 11256 15493 11284 15524
rect 11882 15512 11888 15564
rect 11940 15512 11946 15564
rect 14182 15512 14188 15564
rect 14240 15552 14246 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 14240 15524 14289 15552
rect 14240 15512 14246 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 14366 15512 14372 15564
rect 14424 15552 14430 15564
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 14424 15524 14749 15552
rect 14424 15512 14430 15524
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 14844 15524 15792 15552
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 13078 15484 13084 15496
rect 11471 15456 13084 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 14844 15484 14872 15524
rect 13412 15456 14872 15484
rect 15013 15487 15071 15493
rect 13412 15444 13418 15456
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 4856 15388 6224 15416
rect 8113 15419 8171 15425
rect 4856 15376 4862 15388
rect 5828 15360 5856 15388
rect 8113 15385 8125 15419
rect 8159 15385 8171 15419
rect 8113 15379 8171 15385
rect 2869 15351 2927 15357
rect 2869 15317 2881 15351
rect 2915 15348 2927 15351
rect 3050 15348 3056 15360
rect 2915 15320 3056 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 3050 15308 3056 15320
rect 3108 15348 3114 15360
rect 3878 15348 3884 15360
rect 3108 15320 3884 15348
rect 3108 15308 3114 15320
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 3970 15308 3976 15360
rect 4028 15308 4034 15360
rect 5810 15308 5816 15360
rect 5868 15308 5874 15360
rect 6454 15308 6460 15360
rect 6512 15348 6518 15360
rect 8128 15348 8156 15379
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 12141 15419 12199 15425
rect 12141 15416 12153 15419
rect 9640 15388 11376 15416
rect 9640 15376 9646 15388
rect 6512 15320 8156 15348
rect 6512 15308 6518 15320
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 8297 15351 8355 15357
rect 8297 15348 8309 15351
rect 8260 15320 8309 15348
rect 8260 15308 8266 15320
rect 8297 15317 8309 15320
rect 8343 15317 8355 15351
rect 8297 15311 8355 15317
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 8996 15320 9413 15348
rect 8996 15308 9002 15320
rect 9401 15317 9413 15320
rect 9447 15317 9459 15351
rect 9401 15311 9459 15317
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 11348 15348 11376 15388
rect 12084 15388 12153 15416
rect 12084 15348 12112 15388
rect 12141 15385 12153 15388
rect 12187 15385 12199 15419
rect 12141 15379 12199 15385
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 15028 15416 15056 15447
rect 15654 15444 15660 15496
rect 15712 15444 15718 15496
rect 15764 15484 15792 15524
rect 16298 15512 16304 15564
rect 16356 15552 16362 15564
rect 16758 15552 16764 15564
rect 16356 15524 16764 15552
rect 16356 15512 16362 15524
rect 16758 15512 16764 15524
rect 16816 15552 16822 15564
rect 16816 15524 16896 15552
rect 16816 15512 16822 15524
rect 16868 15493 16896 15524
rect 16669 15487 16727 15493
rect 16669 15484 16681 15487
rect 15764 15456 16681 15484
rect 16669 15453 16681 15456
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15453 16911 15487
rect 16960 15484 16988 15592
rect 17678 15580 17684 15632
rect 17736 15620 17742 15632
rect 18785 15623 18843 15629
rect 18785 15620 18797 15623
rect 17736 15592 18797 15620
rect 17736 15580 17742 15592
rect 18785 15589 18797 15592
rect 18831 15589 18843 15623
rect 18785 15583 18843 15589
rect 20162 15580 20168 15632
rect 20220 15620 20226 15632
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20220 15592 20637 15620
rect 20220 15580 20226 15592
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 17218 15512 17224 15564
rect 17276 15552 17282 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17276 15524 17877 15552
rect 17276 15512 17282 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 18414 15512 18420 15564
rect 18472 15552 18478 15564
rect 20070 15552 20076 15564
rect 18472 15524 20076 15552
rect 18472 15512 18478 15524
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 16960 15456 17509 15484
rect 16853 15447 16911 15453
rect 17497 15453 17509 15456
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 17678 15444 17684 15496
rect 17736 15444 17742 15496
rect 18647 15453 18705 15459
rect 18322 15416 18328 15428
rect 12860 15388 15056 15416
rect 15488 15388 18328 15416
rect 12860 15376 12866 15388
rect 11348 15320 12112 15348
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13265 15351 13323 15357
rect 13265 15348 13277 15351
rect 12768 15320 13277 15348
rect 12768 15308 12774 15320
rect 13265 15317 13277 15320
rect 13311 15317 13323 15351
rect 13265 15311 13323 15317
rect 14921 15351 14979 15357
rect 14921 15317 14933 15351
rect 14967 15348 14979 15351
rect 15286 15348 15292 15360
rect 14967 15320 15292 15348
rect 14967 15317 14979 15320
rect 14921 15311 14979 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 15488 15357 15516 15388
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 18414 15376 18420 15428
rect 18472 15376 18478 15428
rect 18647 15419 18659 15453
rect 18693 15428 18705 15453
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19024 15456 19441 15484
rect 19024 15444 19030 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 18693 15419 18696 15428
rect 18647 15413 18696 15419
rect 18672 15388 18696 15413
rect 18690 15376 18696 15388
rect 18748 15376 18754 15428
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 18840 15388 19625 15416
rect 18840 15376 18846 15388
rect 19613 15385 19625 15388
rect 19659 15416 19671 15419
rect 19996 15416 20024 15524
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 21100 15552 21128 15660
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 21358 15688 21364 15700
rect 21232 15660 21364 15688
rect 21232 15648 21238 15660
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21637 15691 21695 15697
rect 21637 15657 21649 15691
rect 21683 15688 21695 15691
rect 23201 15691 23259 15697
rect 21683 15660 22094 15688
rect 21683 15657 21695 15660
rect 21637 15651 21695 15657
rect 21818 15580 21824 15632
rect 21876 15580 21882 15632
rect 22066 15620 22094 15660
rect 23201 15657 23213 15691
rect 23247 15688 23259 15691
rect 24946 15688 24952 15700
rect 23247 15660 24952 15688
rect 23247 15657 23259 15660
rect 23201 15651 23259 15657
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 25590 15648 25596 15700
rect 25648 15688 25654 15700
rect 28169 15691 28227 15697
rect 28169 15688 28181 15691
rect 25648 15660 28181 15688
rect 25648 15648 25654 15660
rect 28169 15657 28181 15660
rect 28215 15657 28227 15691
rect 28169 15651 28227 15657
rect 23109 15623 23167 15629
rect 23109 15620 23121 15623
rect 22066 15592 23121 15620
rect 23109 15589 23121 15592
rect 23155 15589 23167 15623
rect 23109 15583 23167 15589
rect 22738 15552 22744 15564
rect 21100 15524 22744 15552
rect 22738 15512 22744 15524
rect 22796 15512 22802 15564
rect 23124 15552 23152 15583
rect 25958 15580 25964 15632
rect 26016 15580 26022 15632
rect 23124 15524 24716 15552
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 21542 15484 21548 15496
rect 20220 15456 21548 15484
rect 20220 15444 20226 15456
rect 20487 15453 20545 15456
rect 20257 15419 20315 15425
rect 20257 15416 20269 15419
rect 19659 15388 19932 15416
rect 19996 15388 20269 15416
rect 19659 15385 19671 15388
rect 19613 15379 19671 15385
rect 15473 15351 15531 15357
rect 15473 15317 15485 15351
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 15562 15308 15568 15360
rect 15620 15348 15626 15360
rect 16850 15348 16856 15360
rect 15620 15320 16856 15348
rect 15620 15308 15626 15320
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 18432 15348 18460 15376
rect 17368 15320 18460 15348
rect 17368 15308 17374 15320
rect 19794 15308 19800 15360
rect 19852 15308 19858 15360
rect 19904 15348 19932 15388
rect 20257 15385 20269 15388
rect 20303 15385 20315 15419
rect 20487 15419 20499 15453
rect 20533 15419 20545 15453
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21692 15456 22094 15484
rect 21692 15444 21698 15456
rect 20487 15413 20545 15419
rect 20257 15379 20315 15385
rect 21082 15376 21088 15428
rect 21140 15416 21146 15428
rect 21453 15419 21511 15425
rect 21453 15416 21465 15419
rect 21140 15388 21465 15416
rect 21140 15376 21146 15388
rect 21453 15385 21465 15388
rect 21499 15385 21511 15419
rect 22066 15416 22094 15456
rect 24026 15444 24032 15496
rect 24084 15484 24090 15496
rect 24578 15484 24584 15496
rect 24084 15456 24584 15484
rect 24084 15444 24090 15456
rect 24578 15444 24584 15456
rect 24636 15444 24642 15496
rect 24688 15484 24716 15524
rect 25774 15484 25780 15496
rect 24688 15456 25780 15484
rect 25774 15444 25780 15456
rect 25832 15444 25838 15496
rect 26418 15444 26424 15496
rect 26476 15484 26482 15496
rect 27062 15493 27068 15496
rect 26789 15487 26847 15493
rect 26789 15484 26801 15487
rect 26476 15456 26801 15484
rect 26476 15444 26482 15456
rect 26789 15453 26801 15456
rect 26835 15453 26847 15487
rect 27056 15484 27068 15493
rect 27023 15456 27068 15484
rect 26789 15447 26847 15453
rect 27056 15447 27068 15456
rect 27062 15444 27068 15447
rect 27120 15444 27126 15496
rect 22741 15419 22799 15425
rect 22741 15416 22753 15419
rect 22066 15388 22753 15416
rect 21453 15379 21511 15385
rect 22741 15385 22753 15388
rect 22787 15385 22799 15419
rect 22741 15379 22799 15385
rect 21174 15348 21180 15360
rect 19904 15320 21180 15348
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 21653 15351 21711 15357
rect 21653 15348 21665 15351
rect 21600 15320 21665 15348
rect 21600 15308 21606 15320
rect 21653 15317 21665 15320
rect 21699 15317 21711 15351
rect 22756 15348 22784 15379
rect 23198 15376 23204 15428
rect 23256 15416 23262 15428
rect 23753 15419 23811 15425
rect 23753 15416 23765 15419
rect 23256 15388 23765 15416
rect 23256 15376 23262 15388
rect 23753 15385 23765 15388
rect 23799 15385 23811 15419
rect 23753 15379 23811 15385
rect 24848 15419 24906 15425
rect 24848 15385 24860 15419
rect 24894 15416 24906 15419
rect 28074 15416 28080 15428
rect 24894 15388 28080 15416
rect 24894 15385 24906 15388
rect 24848 15379 24906 15385
rect 28074 15376 28080 15388
rect 28132 15376 28138 15428
rect 23474 15348 23480 15360
rect 22756 15320 23480 15348
rect 21653 15311 21711 15317
rect 23474 15308 23480 15320
rect 23532 15348 23538 15360
rect 23845 15351 23903 15357
rect 23845 15348 23857 15351
rect 23532 15320 23857 15348
rect 23532 15308 23538 15320
rect 23845 15317 23857 15320
rect 23891 15348 23903 15351
rect 27522 15348 27528 15360
rect 23891 15320 27528 15348
rect 23891 15317 23903 15320
rect 23845 15311 23903 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 1765 15147 1823 15153
rect 1765 15113 1777 15147
rect 1811 15144 1823 15147
rect 1854 15144 1860 15156
rect 1811 15116 1860 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 5626 15144 5632 15156
rect 3568 15116 5632 15144
rect 3568 15104 3574 15116
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 6730 15144 6736 15156
rect 6472 15116 6736 15144
rect 1670 15036 1676 15088
rect 1728 15076 1734 15088
rect 6472 15076 6500 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 7248 15116 7389 15144
rect 7248 15104 7254 15116
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 7558 15104 7564 15156
rect 7616 15104 7622 15156
rect 8202 15104 8208 15156
rect 8260 15104 8266 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8904 15116 8953 15144
rect 8904 15104 8910 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 8941 15107 8999 15113
rect 9030 15104 9036 15156
rect 9088 15144 9094 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9088 15116 9321 15144
rect 9088 15104 9094 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 12434 15144 12440 15156
rect 10735 15116 12440 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 12434 15104 12440 15116
rect 12492 15104 12498 15156
rect 12529 15147 12587 15153
rect 12529 15113 12541 15147
rect 12575 15144 12587 15147
rect 12986 15144 12992 15156
rect 12575 15116 12992 15144
rect 12575 15113 12587 15116
rect 12529 15107 12587 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 13136 15116 14228 15144
rect 13136 15104 13142 15116
rect 10778 15076 10784 15088
rect 1728 15048 6500 15076
rect 6564 15048 10784 15076
rect 1728 15036 1734 15048
rect 1946 14968 1952 15020
rect 2004 14968 2010 15020
rect 2038 14968 2044 15020
rect 2096 14968 2102 15020
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2056 14872 2084 14968
rect 2240 14940 2268 14971
rect 2314 14968 2320 15020
rect 2372 14968 2378 15020
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 4396 14980 5549 15008
rect 4396 14968 4402 14980
rect 5537 14977 5549 14980
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 3326 14940 3332 14952
rect 2240 14912 3332 14940
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 4430 14940 4436 14952
rect 3844 14912 4436 14940
rect 3844 14900 3850 14912
rect 4430 14900 4436 14912
rect 4488 14940 4494 14952
rect 5718 14940 5724 14952
rect 4488 14912 5724 14940
rect 4488 14900 4494 14912
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 2682 14872 2688 14884
rect 2056 14844 2688 14872
rect 2682 14832 2688 14844
rect 2740 14872 2746 14884
rect 5350 14872 5356 14884
rect 2740 14844 5356 14872
rect 2740 14832 2746 14844
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 6564 14872 6592 15048
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 11701 15079 11759 15085
rect 11701 15045 11713 15079
rect 11747 15076 11759 15079
rect 11917 15079 11975 15085
rect 11747 15048 11836 15076
rect 11747 15045 11759 15048
rect 11701 15039 11759 15045
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 6788 14980 6914 15008
rect 6788 14968 6794 14980
rect 5644 14844 6592 14872
rect 6886 14872 6914 14980
rect 8294 14968 8300 15020
rect 8352 14968 8358 15020
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 8444 14980 8493 15008
rect 8444 14968 8450 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 10137 15011 10195 15017
rect 10137 15008 10149 15011
rect 9824 14980 10149 15008
rect 9824 14968 9830 14980
rect 10137 14977 10149 14980
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 10284 14980 10425 15008
rect 10284 14968 10290 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 11808 15008 11836 15048
rect 11917 15045 11929 15079
rect 11963 15076 11975 15079
rect 12250 15076 12256 15088
rect 11963 15048 12256 15076
rect 11963 15045 11975 15048
rect 11917 15039 11975 15045
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 13814 15076 13820 15088
rect 12728 15048 13820 15076
rect 12618 15008 12624 15020
rect 11808 14980 12624 15008
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12728 15017 12756 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 13412 14980 13461 15008
rect 13412 14968 13418 14980
rect 13449 14977 13461 14980
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 13596 14980 13737 15008
rect 13596 14968 13602 14980
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13998 14968 14004 15020
rect 14056 14968 14062 15020
rect 14200 15017 14228 15116
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15010 15144 15016 15156
rect 14792 15116 15016 15144
rect 14792 15104 14798 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 16022 15104 16028 15156
rect 16080 15104 16086 15156
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17862 15144 17868 15156
rect 17543 15116 17868 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18049 15147 18107 15153
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 20714 15144 20720 15156
rect 18095 15116 20720 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 22005 15147 22063 15153
rect 22005 15144 22017 15147
rect 20916 15116 22017 15144
rect 16850 15036 16856 15088
rect 16908 15076 16914 15088
rect 17034 15076 17040 15088
rect 16908 15048 17040 15076
rect 16908 15036 16914 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 19794 15076 19800 15088
rect 18248 15048 19800 15076
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 14792 14980 15117 15008
rect 14792 14968 14798 14980
rect 15105 14977 15117 14980
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 8628 14912 9413 14940
rect 8628 14900 8634 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14909 15347 14943
rect 15396 14940 15424 14971
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 15804 14980 16221 15008
rect 15804 14968 15810 14980
rect 16209 14977 16221 14980
rect 16255 14977 16267 15011
rect 16209 14971 16267 14977
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 17129 15011 17187 15017
rect 17129 15008 17141 15011
rect 16632 14980 17141 15008
rect 16632 14968 16638 14980
rect 17129 14977 17141 14980
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 15008 17647 15011
rect 18046 15008 18052 15020
rect 17635 14980 18052 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 18248 15017 18276 15048
rect 19794 15036 19800 15048
rect 19852 15036 19858 15088
rect 19886 15036 19892 15088
rect 19944 15076 19950 15088
rect 20916 15076 20944 15116
rect 22005 15113 22017 15116
rect 22051 15113 22063 15147
rect 22005 15107 22063 15113
rect 23109 15147 23167 15153
rect 23109 15113 23121 15147
rect 23155 15144 23167 15147
rect 24854 15144 24860 15156
rect 23155 15116 24860 15144
rect 23155 15113 23167 15116
rect 23109 15107 23167 15113
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 28077 15147 28135 15153
rect 28077 15113 28089 15147
rect 28123 15144 28135 15147
rect 28166 15144 28172 15156
rect 28123 15116 28172 15144
rect 28123 15113 28135 15116
rect 28077 15107 28135 15113
rect 28166 15104 28172 15116
rect 28224 15104 28230 15156
rect 19944 15048 20944 15076
rect 20993 15079 21051 15085
rect 19944 15036 19950 15048
rect 20993 15045 21005 15079
rect 21039 15076 21051 15079
rect 21634 15076 21640 15088
rect 21039 15048 21640 15076
rect 21039 15045 21051 15048
rect 20993 15039 21051 15045
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 22281 15079 22339 15085
rect 22281 15045 22293 15079
rect 22327 15076 22339 15079
rect 25866 15076 25872 15088
rect 22327 15048 25872 15076
rect 22327 15045 22339 15048
rect 22281 15039 22339 15045
rect 25866 15036 25872 15048
rect 25924 15076 25930 15088
rect 27798 15076 27804 15088
rect 25924 15048 27804 15076
rect 25924 15036 25930 15048
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18949 15011 19007 15017
rect 18949 15008 18961 15011
rect 18380 14980 18961 15008
rect 18380 14968 18386 14980
rect 18949 14977 18961 14980
rect 18995 14977 19007 15011
rect 18949 14971 19007 14977
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20588 14980 20637 15008
rect 20588 14968 20594 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 14977 20959 15011
rect 21111 15011 21169 15017
rect 21111 15008 21123 15011
rect 20901 14971 20959 14977
rect 21008 14980 21123 15008
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 15396 14912 16865 14940
rect 15289 14903 15347 14909
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 7009 14875 7067 14881
rect 7009 14872 7021 14875
rect 6886 14844 7021 14872
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 2648 14776 4169 14804
rect 2648 14764 2654 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 5644 14813 5672 14844
rect 7009 14841 7021 14844
rect 7055 14872 7067 14875
rect 9214 14872 9220 14884
rect 7055 14844 9220 14872
rect 7055 14841 7067 14844
rect 7009 14835 7067 14841
rect 9214 14832 9220 14844
rect 9272 14872 9278 14884
rect 9508 14872 9536 14903
rect 9272 14844 9536 14872
rect 9272 14832 9278 14844
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 11149 14875 11207 14881
rect 11149 14872 11161 14875
rect 9732 14844 11161 14872
rect 9732 14832 9738 14844
rect 11149 14841 11161 14844
rect 11195 14841 11207 14875
rect 11149 14835 11207 14841
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 12069 14875 12127 14881
rect 11756 14844 12020 14872
rect 11756 14832 11762 14844
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 4304 14776 5641 14804
rect 4304 14764 4310 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 5629 14767 5687 14773
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 5776 14776 7389 14804
rect 5776 14764 5782 14776
rect 7377 14773 7389 14776
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 8018 14764 8024 14816
rect 8076 14764 8082 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 10594 14804 10600 14816
rect 8904 14776 10600 14804
rect 8904 14764 8910 14776
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11848 14776 11897 14804
rect 11848 14764 11854 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 11992 14804 12020 14844
rect 12069 14841 12081 14875
rect 12115 14872 12127 14875
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 12115 14844 13829 14872
rect 12115 14841 12127 14844
rect 12069 14835 12127 14841
rect 13817 14841 13829 14844
rect 13863 14841 13875 14875
rect 13817 14835 13875 14841
rect 13906 14832 13912 14884
rect 13964 14832 13970 14884
rect 14550 14832 14556 14884
rect 14608 14872 14614 14884
rect 15102 14872 15108 14884
rect 14608 14844 15108 14872
rect 14608 14832 14614 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15304 14872 15332 14903
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 18138 14940 18144 14952
rect 17092 14912 18144 14940
rect 17092 14900 17098 14912
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 16114 14872 16120 14884
rect 15304 14844 16120 14872
rect 16114 14832 16120 14844
rect 16172 14832 16178 14884
rect 17313 14875 17371 14881
rect 17313 14872 17325 14875
rect 16224 14844 17325 14872
rect 12250 14804 12256 14816
rect 11992 14776 12256 14804
rect 11885 14767 11943 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 14332 14776 15209 14804
rect 14332 14764 14338 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15197 14767 15255 14773
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 15565 14807 15623 14813
rect 15565 14804 15577 14807
rect 15344 14776 15577 14804
rect 15344 14764 15350 14776
rect 15565 14773 15577 14776
rect 15611 14773 15623 14807
rect 15565 14767 15623 14773
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16224 14804 16252 14844
rect 17313 14841 17325 14844
rect 17359 14841 17371 14875
rect 17313 14835 17371 14841
rect 15988 14776 16252 14804
rect 18708 14804 18736 14903
rect 19978 14900 19984 14952
rect 20036 14940 20042 14952
rect 20824 14940 20852 14971
rect 20036 14912 20852 14940
rect 20036 14900 20042 14912
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 20916 14872 20944 14971
rect 21008 14952 21036 14980
rect 21111 14977 21123 14980
rect 21157 14977 21169 15011
rect 21111 14971 21169 14977
rect 21542 14968 21548 15020
rect 21600 15008 21606 15020
rect 22190 15011 22248 15017
rect 22190 15008 22202 15011
rect 21600 14980 22202 15008
rect 21600 14968 21606 14980
rect 22190 14977 22202 14980
rect 22236 14977 22248 15011
rect 22190 14971 22248 14977
rect 22370 14968 22376 15020
rect 22428 14968 22434 15020
rect 22462 14968 22468 15020
rect 22520 15017 22526 15020
rect 22520 15011 22549 15017
rect 22537 14977 22549 15011
rect 22520 14971 22549 14977
rect 22520 14968 22526 14971
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 24193 15011 24251 15017
rect 24193 15008 24205 15011
rect 23532 14980 24205 15008
rect 23532 14968 23538 14980
rect 24193 14977 24205 14980
rect 24239 14977 24251 15011
rect 24193 14971 24251 14977
rect 20990 14900 20996 14952
rect 21048 14900 21054 14952
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14940 21327 14943
rect 22649 14943 22707 14949
rect 21315 14912 22600 14940
rect 21315 14909 21327 14912
rect 21269 14903 21327 14909
rect 22572 14872 22600 14912
rect 22649 14909 22661 14943
rect 22695 14940 22707 14943
rect 22695 14912 23888 14940
rect 22695 14909 22707 14912
rect 22649 14903 22707 14909
rect 23658 14872 23664 14884
rect 20404 14844 20760 14872
rect 20916 14844 22094 14872
rect 22572 14844 23664 14872
rect 20404 14832 20410 14844
rect 19794 14804 19800 14816
rect 18708 14776 19800 14804
rect 15988 14764 15994 14776
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 20070 14764 20076 14816
rect 20128 14764 20134 14816
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 20622 14804 20628 14816
rect 20312 14776 20628 14804
rect 20312 14764 20318 14776
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 20732 14804 20760 14844
rect 21266 14804 21272 14816
rect 20732 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 22066 14804 22094 14844
rect 23658 14832 23664 14844
rect 23716 14832 23722 14884
rect 23750 14804 23756 14816
rect 22066 14776 23756 14804
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 23860 14804 23888 14912
rect 23934 14900 23940 14952
rect 23992 14900 23998 14952
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27580 14912 27629 14940
rect 27580 14900 27586 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 25958 14832 25964 14884
rect 26016 14872 26022 14884
rect 27893 14875 27951 14881
rect 27893 14872 27905 14875
rect 26016 14844 27905 14872
rect 26016 14832 26022 14844
rect 27893 14841 27905 14844
rect 27939 14841 27951 14875
rect 27893 14835 27951 14841
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 23860 14776 25329 14804
rect 25317 14773 25329 14776
rect 25363 14804 25375 14807
rect 27430 14804 27436 14816
rect 25363 14776 27436 14804
rect 25363 14773 25375 14776
rect 25317 14767 25375 14773
rect 27430 14764 27436 14776
rect 27488 14764 27494 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14600 1731 14603
rect 1946 14600 1952 14612
rect 1719 14572 1952 14600
rect 1719 14569 1731 14572
rect 1673 14563 1731 14569
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14569 3295 14603
rect 3237 14563 3295 14569
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 4154 14600 4160 14612
rect 3467 14572 4160 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 1964 14464 1992 14560
rect 3252 14532 3280 14563
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4985 14603 5043 14609
rect 4985 14569 4997 14603
rect 5031 14600 5043 14603
rect 5258 14600 5264 14612
rect 5031 14572 5264 14600
rect 5031 14569 5043 14572
rect 4985 14563 5043 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 8018 14600 8024 14612
rect 6420 14572 8024 14600
rect 6420 14560 6426 14572
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 8662 14600 8668 14612
rect 8527 14572 8668 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 9490 14560 9496 14612
rect 9548 14560 9554 14612
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 12710 14600 12716 14612
rect 11379 14572 12716 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14600 13323 14603
rect 13722 14600 13728 14612
rect 13311 14572 13728 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 13872 14572 14749 14600
rect 13872 14560 13878 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 15746 14600 15752 14612
rect 15703 14572 15752 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 17313 14603 17371 14609
rect 17313 14600 17325 14603
rect 16264 14572 17325 14600
rect 16264 14560 16270 14572
rect 17313 14569 17325 14572
rect 17359 14569 17371 14603
rect 17313 14563 17371 14569
rect 17589 14603 17647 14609
rect 17589 14569 17601 14603
rect 17635 14600 17647 14603
rect 17954 14600 17960 14612
rect 17635 14572 17960 14600
rect 17635 14569 17647 14572
rect 17589 14563 17647 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 20346 14600 20352 14612
rect 18739 14572 20352 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 20441 14603 20499 14609
rect 20441 14569 20453 14603
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 4062 14532 4068 14544
rect 3252 14504 4068 14532
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 7742 14532 7748 14544
rect 4724 14504 7748 14532
rect 1964 14436 3280 14464
rect 1854 14356 1860 14408
rect 1912 14356 1918 14408
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 3252 14396 3280 14436
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4028 14436 4476 14464
rect 4028 14424 4034 14436
rect 3252 14371 3296 14396
rect 3252 14368 3341 14371
rect 3268 14365 3341 14368
rect 2682 14288 2688 14340
rect 2740 14328 2746 14340
rect 3053 14331 3111 14337
rect 3268 14334 3295 14365
rect 3053 14328 3065 14331
rect 2740 14300 3065 14328
rect 2740 14288 2746 14300
rect 3053 14297 3065 14300
rect 3099 14297 3111 14331
rect 3283 14331 3295 14334
rect 3329 14331 3341 14365
rect 4154 14356 4160 14408
rect 4212 14356 4218 14408
rect 4448 14405 4476 14436
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 3283 14325 3341 14331
rect 4264 14328 4292 14359
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 4724 14328 4752 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 11790 14532 11796 14544
rect 7892 14504 9076 14532
rect 7892 14492 7898 14504
rect 9048 14476 9076 14504
rect 10336 14504 11796 14532
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 5132 14436 5457 14464
rect 5132 14424 5138 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 6972 14436 8432 14464
rect 6972 14424 6978 14436
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4856 14368 5181 14396
rect 4856 14356 4862 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5718 14396 5724 14408
rect 5399 14368 5724 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 4264 14300 4752 14328
rect 3053 14291 3111 14297
rect 4890 14288 4896 14340
rect 4948 14328 4954 14340
rect 5276 14328 5304 14359
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6362 14356 6368 14408
rect 6420 14356 6426 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7098 14396 7104 14408
rect 6687 14368 7104 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7248 14368 7573 14396
rect 7248 14356 7254 14368
rect 7561 14365 7573 14368
rect 7607 14396 7619 14399
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7607 14368 8309 14396
rect 7607 14365 7619 14368
rect 7561 14359 7619 14365
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8404 14396 8432 14436
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 9088 14436 9137 14464
rect 9088 14424 9094 14436
rect 9125 14433 9137 14436
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8404 14368 9321 14396
rect 8297 14359 8355 14365
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10226 14396 10232 14408
rect 10183 14368 10232 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10336 14405 10364 14504
rect 11790 14492 11796 14504
rect 11848 14492 11854 14544
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 12032 14504 12081 14532
rect 12032 14492 12038 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12308 14504 13584 14532
rect 12308 14492 12314 14504
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11238 14464 11244 14476
rect 10928 14436 11244 14464
rect 10928 14424 10934 14436
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 11514 14424 11520 14476
rect 11572 14464 11578 14476
rect 12894 14464 12900 14476
rect 11572 14436 12900 14464
rect 11572 14424 11578 14436
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 11624 14405 12020 14406
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14365 10379 14399
rect 11624 14399 12035 14405
rect 11624 14396 11989 14399
rect 10321 14359 10379 14365
rect 11532 14378 11989 14396
rect 11532 14368 11652 14378
rect 4948 14300 5304 14328
rect 4948 14288 4954 14300
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 10870 14328 10876 14340
rect 6512 14300 10876 14328
rect 6512 14288 6518 14300
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 11146 14288 11152 14340
rect 11204 14288 11210 14340
rect 11330 14288 11336 14340
rect 11388 14337 11394 14340
rect 11388 14331 11407 14337
rect 11395 14297 11407 14331
rect 11532 14328 11560 14368
rect 11977 14365 11989 14378
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12250 14396 12256 14408
rect 12207 14368 12256 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 13078 14356 13084 14408
rect 13136 14356 13142 14408
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 11388 14291 11407 14297
rect 11440 14300 11560 14328
rect 13188 14328 13216 14359
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13556 14405 13584 14504
rect 13906 14492 13912 14544
rect 13964 14532 13970 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 13964 14504 14565 14532
rect 13964 14492 13970 14504
rect 14553 14501 14565 14504
rect 14599 14501 14611 14535
rect 14553 14495 14611 14501
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 16022 14532 16028 14544
rect 15611 14504 16028 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 16022 14492 16028 14504
rect 16080 14532 16086 14544
rect 16080 14504 17320 14532
rect 16080 14492 16086 14504
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 14700 14436 16497 14464
rect 14700 14424 14706 14436
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 17034 14464 17040 14476
rect 16485 14427 16543 14433
rect 16684 14436 17040 14464
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13320 14368 13369 14396
rect 13320 14356 13326 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14365 13599 14399
rect 14550 14396 14556 14408
rect 13541 14359 13599 14365
rect 14200 14368 14556 14396
rect 14200 14328 14228 14368
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 15160 14368 16344 14396
rect 15160 14356 15166 14368
rect 13188 14300 14228 14328
rect 15197 14331 15255 14337
rect 11388 14288 11394 14291
rect 2038 14220 2044 14272
rect 2096 14220 2102 14272
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 3973 14263 4031 14269
rect 3973 14260 3985 14263
rect 3016 14232 3985 14260
rect 3016 14220 3022 14232
rect 3973 14229 3985 14232
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5224 14232 6193 14260
rect 5224 14220 5230 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 7006 14260 7012 14272
rect 6595 14232 7012 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 8754 14260 8760 14272
rect 7791 14232 8760 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 8754 14220 8760 14232
rect 8812 14260 8818 14272
rect 9122 14260 9128 14272
rect 8812 14232 9128 14260
rect 8812 14220 8818 14232
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9490 14260 9496 14272
rect 9272 14232 9496 14260
rect 9272 14220 9278 14232
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11440 14260 11468 14300
rect 15197 14297 15209 14331
rect 15243 14328 15255 14331
rect 15378 14328 15384 14340
rect 15243 14300 15384 14328
rect 15243 14297 15255 14300
rect 15197 14291 15255 14297
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 16316 14328 16344 14368
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 16574 14356 16580 14408
rect 16632 14356 16638 14408
rect 16684 14405 16712 14436
rect 17034 14424 17040 14436
rect 17092 14424 17098 14476
rect 17292 14464 17320 14504
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 18877 14535 18935 14541
rect 18877 14532 18889 14535
rect 18104 14504 18889 14532
rect 18104 14492 18110 14504
rect 18877 14501 18889 14504
rect 18923 14501 18935 14535
rect 20456 14532 20484 14563
rect 20622 14560 20628 14612
rect 20680 14560 20686 14612
rect 21453 14603 21511 14609
rect 21453 14569 21465 14603
rect 21499 14600 21511 14603
rect 25958 14600 25964 14612
rect 21499 14572 25964 14600
rect 21499 14569 21511 14572
rect 21453 14563 21511 14569
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 27617 14603 27675 14609
rect 27617 14600 27629 14603
rect 26068 14572 27629 14600
rect 22557 14535 22615 14541
rect 20456 14504 22094 14532
rect 18877 14495 18935 14501
rect 20070 14464 20076 14476
rect 17292 14436 20076 14464
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14396 16911 14399
rect 17126 14396 17132 14408
rect 16899 14368 17132 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14365 17739 14399
rect 17681 14359 17739 14365
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 17696 14328 17724 14359
rect 16316 14300 17724 14328
rect 10836 14232 11468 14260
rect 11517 14263 11575 14269
rect 10836 14220 10842 14232
rect 11517 14229 11529 14263
rect 11563 14260 11575 14263
rect 11974 14260 11980 14272
rect 11563 14232 11980 14260
rect 11563 14229 11575 14232
rect 11517 14223 11575 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12805 14263 12863 14269
rect 12805 14229 12817 14263
rect 12851 14260 12863 14263
rect 14182 14260 14188 14272
rect 12851 14232 14188 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 17788 14260 17816 14359
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18966 14396 18972 14408
rect 18095 14368 18972 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18966 14356 18972 14368
rect 19024 14396 19030 14408
rect 19610 14396 19616 14408
rect 19024 14368 19616 14396
rect 19024 14356 19030 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 21542 14396 21548 14408
rect 20487 14365 20545 14371
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18509 14331 18567 14337
rect 18509 14328 18521 14331
rect 18012 14300 18521 14328
rect 18012 14288 18018 14300
rect 18509 14297 18521 14300
rect 18555 14297 18567 14331
rect 18509 14291 18567 14297
rect 18725 14331 18783 14337
rect 18725 14297 18737 14331
rect 18771 14328 18783 14331
rect 19058 14328 19064 14340
rect 18771 14300 19064 14328
rect 18771 14297 18783 14300
rect 18725 14291 18783 14297
rect 19058 14288 19064 14300
rect 19116 14288 19122 14340
rect 20257 14331 20315 14337
rect 20257 14297 20269 14331
rect 20303 14297 20315 14331
rect 20487 14331 20499 14365
rect 20533 14331 20545 14365
rect 21484 14365 21548 14396
rect 20487 14328 20545 14331
rect 20714 14328 20720 14340
rect 20487 14325 20720 14328
rect 20502 14300 20720 14325
rect 20257 14291 20315 14297
rect 14516 14232 17816 14260
rect 14516 14220 14522 14232
rect 19150 14220 19156 14272
rect 19208 14260 19214 14272
rect 20162 14260 20168 14272
rect 19208 14232 20168 14260
rect 19208 14220 19214 14232
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20272 14260 20300 14291
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 21269 14331 21327 14337
rect 21484 14334 21511 14365
rect 21269 14297 21281 14331
rect 21315 14297 21327 14331
rect 21499 14331 21511 14334
rect 21545 14356 21548 14365
rect 21600 14356 21606 14408
rect 22066 14396 22094 14504
rect 22557 14501 22569 14535
rect 22603 14532 22615 14535
rect 22830 14532 22836 14544
rect 22603 14504 22836 14532
rect 22603 14501 22615 14504
rect 22557 14495 22615 14501
rect 22830 14492 22836 14504
rect 22888 14492 22894 14544
rect 23382 14492 23388 14544
rect 23440 14492 23446 14544
rect 23566 14492 23572 14544
rect 23624 14532 23630 14544
rect 26068 14532 26096 14572
rect 27617 14569 27629 14572
rect 27663 14569 27675 14603
rect 27617 14563 27675 14569
rect 23624 14504 26096 14532
rect 23624 14492 23630 14504
rect 22649 14467 22707 14473
rect 22649 14433 22661 14467
rect 22695 14464 22707 14467
rect 22695 14436 24808 14464
rect 22695 14433 22707 14436
rect 22649 14427 22707 14433
rect 22922 14396 22928 14408
rect 22066 14368 22928 14396
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 24780 14405 24808 14436
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 25409 14399 25467 14405
rect 25409 14396 25421 14399
rect 25004 14368 25421 14396
rect 25004 14356 25010 14368
rect 25409 14365 25421 14368
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 26237 14399 26295 14405
rect 26237 14365 26249 14399
rect 26283 14396 26295 14399
rect 26326 14396 26332 14408
rect 26283 14368 26332 14396
rect 26283 14365 26295 14368
rect 26237 14359 26295 14365
rect 26326 14356 26332 14368
rect 26384 14356 26390 14408
rect 21545 14331 21557 14356
rect 21499 14325 21557 14331
rect 22189 14331 22247 14337
rect 21269 14291 21327 14297
rect 22189 14297 22201 14331
rect 22235 14328 22247 14331
rect 22554 14328 22560 14340
rect 22235 14300 22560 14328
rect 22235 14297 22247 14300
rect 22189 14291 22247 14297
rect 20806 14260 20812 14272
rect 20272 14232 20812 14260
rect 20806 14220 20812 14232
rect 20864 14260 20870 14272
rect 21284 14260 21312 14291
rect 22554 14288 22560 14300
rect 22612 14328 22618 14340
rect 23106 14328 23112 14340
rect 22612 14300 23112 14328
rect 22612 14288 22618 14300
rect 23106 14288 23112 14300
rect 23164 14288 23170 14340
rect 26482 14331 26540 14337
rect 26482 14328 26494 14331
rect 24596 14300 26494 14328
rect 20864 14232 21312 14260
rect 21637 14263 21695 14269
rect 20864 14220 20870 14232
rect 21637 14229 21649 14263
rect 21683 14260 21695 14263
rect 22278 14260 22284 14272
rect 21683 14232 22284 14260
rect 21683 14229 21695 14232
rect 21637 14223 21695 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 23566 14220 23572 14272
rect 23624 14220 23630 14272
rect 23750 14220 23756 14272
rect 23808 14260 23814 14272
rect 24486 14260 24492 14272
rect 23808 14232 24492 14260
rect 23808 14220 23814 14232
rect 24486 14220 24492 14232
rect 24544 14220 24550 14272
rect 24596 14269 24624 14300
rect 26482 14297 26494 14300
rect 26528 14297 26540 14331
rect 26482 14291 26540 14297
rect 24581 14263 24639 14269
rect 24581 14229 24593 14263
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 25225 14263 25283 14269
rect 25225 14229 25237 14263
rect 25271 14260 25283 14263
rect 26694 14260 26700 14272
rect 25271 14232 26700 14260
rect 25271 14229 25283 14232
rect 25225 14223 25283 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 1578 14016 1584 14068
rect 1636 14016 1642 14068
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 2372 14028 5641 14056
rect 2372 14016 2378 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6512 14028 6561 14056
rect 6512 14016 6518 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 7834 14056 7840 14068
rect 6549 14019 6607 14025
rect 7024 14028 7840 14056
rect 1964 13960 3556 13988
rect 1964 13929 1992 13960
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2498 13920 2504 13932
rect 2271 13892 2504 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 1780 13852 1808 13883
rect 2498 13880 2504 13892
rect 2556 13920 2562 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2556 13892 3249 13920
rect 2556 13880 2562 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 2041 13855 2099 13861
rect 1780 13824 1992 13852
rect 1857 13787 1915 13793
rect 1857 13753 1869 13787
rect 1903 13753 1915 13787
rect 1964 13784 1992 13824
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 2774 13852 2780 13864
rect 2087 13824 2780 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 2774 13812 2780 13824
rect 2832 13852 2838 13864
rect 3528 13861 3556 13960
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4120 13960 5580 13988
rect 4120 13948 4126 13960
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 3878 13920 3884 13932
rect 3835 13892 3884 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 4890 13920 4896 13932
rect 4847 13892 4896 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 2832 13824 3433 13852
rect 2832 13812 2838 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3970 13852 3976 13864
rect 3559 13824 3976 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 4246 13812 4252 13864
rect 4304 13852 4310 13864
rect 4816 13852 4844 13883
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 4304 13824 4844 13852
rect 5000 13852 5028 13883
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5552 13929 5580 13960
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5132 13892 5273 13920
rect 5132 13880 5138 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7024 13920 7052 14028
rect 7834 14016 7840 14028
rect 7892 14056 7898 14068
rect 8202 14056 8208 14068
rect 7892 14028 8208 14056
rect 7892 14016 7898 14028
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 9272 14028 9321 14056
rect 9272 14016 9278 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 10134 14056 10140 14068
rect 9309 14019 9367 14025
rect 9876 14028 10140 14056
rect 7558 13988 7564 14000
rect 7208 13960 7564 13988
rect 7208 13954 7236 13960
rect 7098 13929 7236 13954
rect 7558 13948 7564 13960
rect 7616 13948 7622 14000
rect 9490 13988 9496 14000
rect 8496 13960 9496 13988
rect 6871 13892 7052 13920
rect 7083 13926 7236 13929
rect 7083 13923 7141 13926
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7083 13889 7095 13923
rect 7129 13889 7141 13923
rect 7083 13883 7141 13889
rect 5718 13852 5724 13864
rect 5000 13824 5724 13852
rect 4304 13812 4310 13824
rect 3050 13784 3056 13796
rect 1964 13756 3056 13784
rect 1857 13747 1915 13753
rect 1872 13716 1900 13747
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3326 13744 3332 13796
rect 3384 13744 3390 13796
rect 4890 13744 4896 13796
rect 4948 13784 4954 13796
rect 5000 13784 5028 13824
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6748 13852 6776 13883
rect 7926 13880 7932 13932
rect 7984 13880 7990 13932
rect 8202 13880 8208 13932
rect 8260 13880 8266 13932
rect 8496 13929 8524 13960
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 9876 13997 9904 14028
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 11790 14056 11796 14068
rect 10284 14028 11796 14056
rect 10284 14016 10290 14028
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 11940 14028 12839 14056
rect 11940 14016 11946 14028
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 10045 13991 10103 13997
rect 10045 13957 10057 13991
rect 10091 13988 10103 13991
rect 12710 13988 12716 14000
rect 10091 13960 12716 13988
rect 10091 13957 10103 13960
rect 10045 13951 10103 13957
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 12811 13988 12839 14028
rect 13538 14016 13544 14068
rect 13596 14016 13602 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 13872 14028 14289 14056
rect 13872 14016 13878 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 15488 14028 15792 14056
rect 15488 13997 15516 14028
rect 15473 13991 15531 13997
rect 12811 13960 14688 13988
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 8665 13924 8723 13929
rect 8754 13924 8760 13932
rect 8665 13923 8760 13924
rect 8665 13889 8677 13923
rect 8711 13896 8760 13923
rect 8711 13889 8723 13896
rect 8665 13883 8723 13889
rect 8754 13880 8760 13896
rect 8812 13880 8818 13932
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9582 13920 9588 13932
rect 9447 13892 9588 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 7944 13852 7972 13880
rect 6748 13824 7972 13852
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8076 13824 8401 13852
rect 8076 13812 8082 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 9232 13852 9260 13883
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10744 13892 10793 13920
rect 10744 13880 10750 13892
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11957 13923 12015 13929
rect 11957 13920 11969 13923
rect 11204 13892 11969 13920
rect 11204 13880 11210 13892
rect 11957 13889 11969 13892
rect 12003 13889 12015 13923
rect 11957 13883 12015 13889
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 12894 13920 12900 13932
rect 12400 13892 12900 13920
rect 12400 13880 12406 13892
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 14182 13880 14188 13932
rect 14240 13880 14246 13932
rect 14660 13929 14688 13960
rect 15473 13957 15485 13991
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 15654 13948 15660 14000
rect 15712 13997 15718 14000
rect 15712 13991 15731 13997
rect 15719 13957 15731 13991
rect 15764 13988 15792 14028
rect 15838 14016 15844 14068
rect 15896 14016 15902 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 18601 14059 18659 14065
rect 18601 14056 18613 14059
rect 16632 14028 18613 14056
rect 16632 14016 16638 14028
rect 18601 14025 18613 14028
rect 18647 14025 18659 14059
rect 18601 14019 18659 14025
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 19116 14028 20545 14056
rect 19116 14016 19122 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 22186 14056 22192 14068
rect 21315 14028 22192 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23566 14056 23572 14068
rect 22388 14028 23572 14056
rect 17310 13988 17316 14000
rect 15764 13960 17316 13988
rect 15712 13951 15731 13957
rect 15712 13948 15718 13951
rect 17310 13948 17316 13960
rect 17368 13988 17374 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 17368 13960 17417 13988
rect 17368 13948 17374 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17605 13991 17663 13997
rect 17605 13988 17617 13991
rect 17405 13951 17463 13957
rect 17512 13960 17617 13988
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15562 13920 15568 13932
rect 14967 13892 15568 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 9766 13852 9772 13864
rect 9232 13824 9772 13852
rect 8389 13815 8447 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13852 10287 13855
rect 10870 13852 10876 13864
rect 10275 13824 10876 13852
rect 10275 13821 10287 13824
rect 10229 13815 10287 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11698 13812 11704 13864
rect 11756 13812 11762 13864
rect 4948 13756 5028 13784
rect 4948 13744 4954 13756
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 7006 13784 7012 13796
rect 6696 13756 7012 13784
rect 6696 13744 6702 13756
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 10410 13744 10416 13796
rect 10468 13784 10474 13796
rect 11057 13787 11115 13793
rect 11057 13784 11069 13787
rect 10468 13756 11069 13784
rect 10468 13744 10474 13756
rect 11057 13753 11069 13756
rect 11103 13784 11115 13787
rect 11514 13784 11520 13796
rect 11103 13756 11520 13784
rect 11103 13753 11115 13756
rect 11057 13747 11115 13753
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 14476 13784 14504 13883
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15688 13920 15716 13948
rect 16022 13920 16028 13932
rect 15688 13892 16028 13920
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 16850 13880 16856 13932
rect 16908 13920 16914 13932
rect 17512 13920 17540 13960
rect 17605 13957 17617 13960
rect 17651 13957 17663 13991
rect 17605 13951 17663 13957
rect 17954 13948 17960 14000
rect 18012 13988 18018 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 18012 13960 18245 13988
rect 18012 13948 18018 13960
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 18690 13988 18696 14000
rect 18478 13963 18696 13988
rect 18233 13951 18291 13957
rect 18463 13960 18696 13963
rect 18463 13957 18521 13960
rect 18322 13920 18328 13932
rect 16908 13892 18328 13920
rect 16908 13880 16914 13892
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18463 13923 18475 13957
rect 18509 13923 18521 13957
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 19429 13991 19487 13997
rect 19429 13957 19441 13991
rect 19475 13988 19487 13991
rect 20162 13988 20168 14000
rect 19475 13960 20168 13988
rect 19475 13957 19487 13960
rect 19429 13951 19487 13957
rect 20162 13948 20168 13960
rect 20220 13948 20226 14000
rect 20257 13991 20315 13997
rect 20257 13957 20269 13991
rect 20303 13988 20315 13991
rect 22388 13988 22416 14028
rect 23566 14016 23572 14028
rect 23624 14016 23630 14068
rect 24029 14059 24087 14065
rect 24029 14025 24041 14059
rect 24075 14056 24087 14059
rect 24210 14056 24216 14068
rect 24075 14028 24216 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 24486 14016 24492 14068
rect 24544 14056 24550 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 24544 14028 26617 14056
rect 24544 14016 24550 14028
rect 26605 14025 26617 14028
rect 26651 14025 26663 14059
rect 26605 14019 26663 14025
rect 28074 14016 28080 14068
rect 28132 14016 28138 14068
rect 20303 13960 21312 13988
rect 20303 13957 20315 13960
rect 20257 13951 20315 13957
rect 21284 13932 21312 13960
rect 21468 13960 22416 13988
rect 18463 13917 18521 13923
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 19208 13892 19257 13920
rect 19208 13880 19214 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 19886 13880 19892 13932
rect 19944 13880 19950 13932
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 20354 13923 20412 13929
rect 20354 13920 20366 13923
rect 20180 13892 20366 13920
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15746 13852 15752 13864
rect 15528 13824 15752 13852
rect 15528 13812 15534 13824
rect 15746 13812 15752 13824
rect 15804 13852 15810 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 15804 13824 19073 13852
rect 15804 13812 15810 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 20180 13852 20208 13892
rect 20354 13889 20366 13892
rect 20400 13920 20412 13923
rect 20530 13920 20536 13932
rect 20400 13892 20536 13920
rect 20400 13889 20412 13892
rect 20354 13883 20412 13889
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 21266 13880 21272 13932
rect 21324 13880 21330 13932
rect 21468 13929 21496 13960
rect 22462 13948 22468 14000
rect 22520 13997 22526 14000
rect 25498 13997 25504 14000
rect 22520 13991 22549 13997
rect 22537 13957 22549 13991
rect 25492 13988 25504 13997
rect 25459 13960 25504 13988
rect 22520 13951 22549 13957
rect 25492 13951 25504 13960
rect 22520 13948 22526 13951
rect 25498 13948 25504 13951
rect 25556 13948 25562 14000
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 21542 13880 21548 13932
rect 21600 13920 21606 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21600 13892 22201 13920
rect 21600 13880 21606 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 22374 13923 22432 13929
rect 22374 13889 22386 13923
rect 22420 13889 22432 13923
rect 22374 13883 22432 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22695 13892 24164 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 19668 13824 20208 13852
rect 19668 13812 19674 13824
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 20680 13824 22017 13852
rect 20680 13812 20686 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22296 13852 22324 13883
rect 22152 13824 22324 13852
rect 22152 13812 22158 13824
rect 14240 13756 14504 13784
rect 14240 13744 14246 13756
rect 16942 13744 16948 13796
rect 17000 13784 17006 13796
rect 17494 13784 17500 13796
rect 17000 13756 17500 13784
rect 17000 13744 17006 13756
rect 17494 13744 17500 13756
rect 17552 13744 17558 13796
rect 18432 13756 21496 13784
rect 3605 13719 3663 13725
rect 3605 13716 3617 13719
rect 1872 13688 3617 13716
rect 3605 13685 3617 13688
rect 3651 13716 3663 13719
rect 4982 13716 4988 13728
rect 3651 13688 4988 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5442 13716 5448 13728
rect 5316 13688 5448 13716
rect 5316 13676 5322 13688
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 6454 13676 6460 13728
rect 6512 13716 6518 13728
rect 9306 13716 9312 13728
rect 6512 13688 9312 13716
rect 6512 13676 6518 13688
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 12066 13716 12072 13728
rect 11020 13688 12072 13716
rect 11020 13676 11026 13688
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 13081 13719 13139 13725
rect 13081 13716 13093 13719
rect 12676 13688 13093 13716
rect 12676 13676 12682 13688
rect 13081 13685 13093 13688
rect 13127 13716 13139 13719
rect 13262 13716 13268 13728
rect 13127 13688 13268 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 15286 13716 15292 13728
rect 13780 13688 15292 13716
rect 13780 13676 13786 13688
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15654 13676 15660 13728
rect 15712 13676 15718 13728
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17589 13719 17647 13725
rect 17589 13716 17601 13719
rect 17184 13688 17601 13716
rect 17184 13676 17190 13688
rect 17589 13685 17601 13688
rect 17635 13685 17647 13719
rect 17589 13679 17647 13685
rect 17770 13676 17776 13728
rect 17828 13676 17834 13728
rect 18432 13725 18460 13756
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 19610 13716 19616 13728
rect 18564 13688 19616 13716
rect 18564 13676 18570 13688
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 21468 13716 21496 13756
rect 21634 13744 21640 13796
rect 21692 13784 21698 13796
rect 22388 13784 22416 13883
rect 23106 13812 23112 13864
rect 23164 13812 23170 13864
rect 24136 13852 24164 13892
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 28258 13880 28264 13932
rect 28316 13880 28322 13932
rect 24946 13852 24952 13864
rect 24136 13824 24952 13852
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25188 13824 25237 13852
rect 25188 13812 25194 13824
rect 25225 13821 25237 13824
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 27154 13812 27160 13864
rect 27212 13812 27218 13864
rect 22830 13784 22836 13796
rect 21692 13756 22416 13784
rect 22572 13756 22836 13784
rect 21692 13744 21698 13756
rect 22572 13728 22600 13756
rect 22830 13744 22836 13756
rect 22888 13744 22894 13796
rect 23385 13787 23443 13793
rect 23385 13753 23397 13787
rect 23431 13784 23443 13787
rect 23431 13756 23704 13784
rect 23431 13753 23443 13756
rect 23385 13747 23443 13753
rect 22554 13716 22560 13728
rect 21468 13688 22560 13716
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 23400 13716 23428 13747
rect 22796 13688 23428 13716
rect 22796 13676 22802 13688
rect 23566 13676 23572 13728
rect 23624 13676 23630 13728
rect 23676 13716 23704 13756
rect 27430 13744 27436 13796
rect 27488 13744 27494 13796
rect 25038 13716 25044 13728
rect 23676 13688 25044 13716
rect 25038 13676 25044 13688
rect 25096 13676 25102 13728
rect 27614 13676 27620 13728
rect 27672 13676 27678 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2096 13484 2774 13512
rect 2096 13472 2102 13484
rect 2746 13444 2774 13484
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 5258 13512 5264 13524
rect 3200 13484 5264 13512
rect 3200 13472 3206 13484
rect 5258 13472 5264 13484
rect 5316 13512 5322 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 5316 13484 5457 13512
rect 5316 13472 5322 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 9125 13515 9183 13521
rect 5868 13484 9076 13512
rect 5868 13472 5874 13484
rect 3053 13447 3111 13453
rect 3053 13444 3065 13447
rect 2746 13416 3065 13444
rect 3053 13413 3065 13416
rect 3099 13444 3111 13447
rect 4706 13444 4712 13456
rect 3099 13416 4712 13444
rect 3099 13413 3111 13416
rect 3053 13407 3111 13413
rect 4706 13404 4712 13416
rect 4764 13444 4770 13456
rect 4890 13444 4896 13456
rect 4764 13416 4896 13444
rect 4764 13404 4770 13416
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13413 5687 13447
rect 5629 13407 5687 13413
rect 5166 13376 5172 13388
rect 2746 13348 5172 13376
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 1940 13311 1998 13317
rect 1940 13277 1952 13311
rect 1986 13308 1998 13311
rect 2746 13308 2774 13348
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 5644 13376 5672 13407
rect 6546 13404 6552 13456
rect 6604 13444 6610 13456
rect 8481 13447 8539 13453
rect 8481 13444 8493 13447
rect 6604 13416 8493 13444
rect 6604 13404 6610 13416
rect 8481 13413 8493 13416
rect 8527 13413 8539 13447
rect 9048 13444 9076 13484
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9858 13512 9864 13524
rect 9171 13484 9864 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 11146 13512 11152 13524
rect 10183 13484 11152 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 11330 13472 11336 13524
rect 11388 13512 11394 13524
rect 11388 13484 12434 13512
rect 11388 13472 11394 13484
rect 9490 13444 9496 13456
rect 9048 13416 9496 13444
rect 8481 13407 8539 13413
rect 9490 13404 9496 13416
rect 9548 13404 9554 13456
rect 9582 13404 9588 13456
rect 9640 13404 9646 13456
rect 11057 13447 11115 13453
rect 11057 13413 11069 13447
rect 11103 13444 11115 13447
rect 12158 13444 12164 13456
rect 11103 13416 12164 13444
rect 11103 13413 11115 13416
rect 11057 13407 11115 13413
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 12406 13444 12434 13484
rect 13354 13472 13360 13524
rect 13412 13472 13418 13524
rect 14553 13515 14611 13521
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 17402 13512 17408 13524
rect 14599 13484 17408 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 21269 13515 21327 13521
rect 17512 13484 20944 13512
rect 13814 13444 13820 13456
rect 12406 13416 13820 13444
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 17512 13444 17540 13484
rect 16724 13416 17540 13444
rect 16724 13404 16730 13416
rect 17770 13404 17776 13456
rect 17828 13404 17834 13456
rect 5500 13348 5672 13376
rect 5500 13336 5506 13348
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 6972 13348 7604 13376
rect 6972 13336 6978 13348
rect 1986 13280 2774 13308
rect 1986 13277 1998 13280
rect 1940 13271 1998 13277
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 4120 13280 4261 13308
rect 4120 13268 4126 13280
rect 4249 13277 4261 13280
rect 4295 13277 4307 13311
rect 4614 13308 4620 13320
rect 4249 13271 4307 13277
rect 4356 13280 4620 13308
rect 3602 13200 3608 13252
rect 3660 13240 3666 13252
rect 4356 13240 4384 13280
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4948 13280 5089 13308
rect 4948 13268 4954 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 5684 13280 6653 13308
rect 5684 13268 5690 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6641 13271 6699 13277
rect 6932 13280 7113 13308
rect 3660 13212 4384 13240
rect 4448 13212 6224 13240
rect 3660 13200 3666 13212
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4448 13181 4476 13212
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4212 13144 4445 13172
rect 4212 13132 4218 13144
rect 4433 13141 4445 13144
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5442 13172 5448 13184
rect 4672 13144 5448 13172
rect 4672 13132 4678 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6196 13172 6224 13212
rect 6270 13200 6276 13252
rect 6328 13200 6334 13252
rect 6454 13200 6460 13252
rect 6512 13200 6518 13252
rect 6362 13172 6368 13184
rect 6196 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13172 6426 13184
rect 6932 13172 6960 13280
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7576 13317 7604 13348
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 10134 13376 10140 13388
rect 7892 13348 10140 13376
rect 7892 13336 7898 13348
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10962 13376 10968 13388
rect 10827 13348 10968 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 12989 13379 13047 13385
rect 12989 13376 13001 13379
rect 11204 13348 13001 13376
rect 11204 13336 11210 13348
rect 12989 13345 13001 13348
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 19334 13376 19340 13388
rect 17292 13348 19340 13376
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7650 13308 7656 13320
rect 7607 13280 7656 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8478 13308 8484 13320
rect 8251 13280 8484 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 6420 13144 6960 13172
rect 6420 13132 6426 13144
rect 7282 13132 7288 13184
rect 7340 13132 7346 13184
rect 8036 13172 8064 13271
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 8662 13308 8668 13320
rect 8619 13280 8668 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 9416 13240 9444 13271
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9548 13280 9689 13308
rect 9548 13268 9554 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10502 13308 10508 13320
rect 10367 13280 10508 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 12342 13308 12348 13320
rect 10888 13280 12348 13308
rect 10888 13240 10916 13280
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12492 13280 13093 13308
rect 12492 13268 12498 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 13504 13280 14565 13308
rect 13504 13268 13510 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 11330 13240 11336 13252
rect 9416 13212 10916 13240
rect 10980 13212 11336 13240
rect 8754 13172 8760 13184
rect 8036 13144 8760 13172
rect 8754 13132 8760 13144
rect 8812 13172 8818 13184
rect 10980 13172 11008 13212
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 11701 13243 11759 13249
rect 11701 13209 11713 13243
rect 11747 13240 11759 13243
rect 11790 13240 11796 13252
rect 11747 13212 11796 13240
rect 11747 13209 11759 13212
rect 11701 13203 11759 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 11885 13243 11943 13249
rect 11885 13209 11897 13243
rect 11931 13240 11943 13243
rect 13998 13240 14004 13252
rect 11931 13212 14004 13240
rect 11931 13209 11943 13212
rect 11885 13203 11943 13209
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14277 13243 14335 13249
rect 14277 13209 14289 13243
rect 14323 13240 14335 13243
rect 15470 13240 15476 13252
rect 14323 13212 15476 13240
rect 14323 13209 14335 13212
rect 14277 13203 14335 13209
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 8812 13144 11008 13172
rect 8812 13132 8818 13144
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 11204 13144 11253 13172
rect 11204 13132 11210 13144
rect 11241 13141 11253 13144
rect 11287 13141 11299 13175
rect 11241 13135 11299 13141
rect 11422 13132 11428 13184
rect 11480 13172 11486 13184
rect 12069 13175 12127 13181
rect 12069 13172 12081 13175
rect 11480 13144 12081 13172
rect 11480 13132 11486 13144
rect 12069 13141 12081 13144
rect 12115 13141 12127 13175
rect 12069 13135 12127 13141
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 13354 13172 13360 13184
rect 12400 13144 13360 13172
rect 12400 13132 12406 13144
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 13504 13144 14749 13172
rect 13504 13132 13510 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 15948 13172 15976 13271
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 17292 13317 17320 13348
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 20622 13376 20628 13388
rect 19996 13348 20628 13376
rect 17277 13311 17335 13317
rect 17277 13277 17289 13311
rect 17323 13277 17335 13311
rect 17277 13271 17335 13277
rect 17591 13268 17597 13320
rect 17649 13268 17655 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18417 13311 18475 13317
rect 18417 13308 18429 13311
rect 18012 13280 18429 13308
rect 18012 13268 18018 13280
rect 18417 13277 18429 13280
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 18782 13308 18788 13320
rect 18647 13280 18788 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 19996 13317 20024 13348
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 20916 13376 20944 13484
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 21542 13512 21548 13524
rect 21315 13484 21548 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23934 13512 23940 13524
rect 23164 13484 23940 13512
rect 23164 13472 23170 13484
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24029 13515 24087 13521
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24210 13512 24216 13524
rect 24075 13484 24216 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 24854 13512 24860 13524
rect 24320 13484 24860 13512
rect 20990 13404 20996 13456
rect 21048 13444 21054 13456
rect 21453 13447 21511 13453
rect 21453 13444 21465 13447
rect 21048 13416 21465 13444
rect 21048 13404 21054 13416
rect 21453 13413 21465 13416
rect 21499 13413 21511 13447
rect 21453 13407 21511 13413
rect 22738 13404 22744 13456
rect 22796 13404 22802 13456
rect 23845 13447 23903 13453
rect 23845 13413 23857 13447
rect 23891 13444 23903 13447
rect 24320 13444 24348 13484
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 24946 13472 24952 13524
rect 25004 13512 25010 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25004 13484 25973 13512
rect 25004 13472 25010 13484
rect 25961 13481 25973 13484
rect 26007 13512 26019 13515
rect 26142 13512 26148 13524
rect 26007 13484 26148 13512
rect 26007 13481 26019 13484
rect 25961 13475 26019 13481
rect 26142 13472 26148 13484
rect 26200 13472 26206 13524
rect 27154 13512 27160 13524
rect 26252 13484 27160 13512
rect 23891 13416 24348 13444
rect 23891 13413 23903 13416
rect 23845 13407 23903 13413
rect 23860 13376 23888 13407
rect 20916 13348 23888 13376
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 23992 13348 24716 13376
rect 23992 13336 23998 13348
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20074 13311 20132 13317
rect 20074 13277 20086 13311
rect 20120 13277 20132 13311
rect 20074 13271 20132 13277
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 17000 13212 17417 13240
rect 17000 13200 17006 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 19242 13240 19248 13252
rect 17543 13212 19248 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 19242 13200 19248 13212
rect 19300 13200 19306 13252
rect 19886 13200 19892 13252
rect 19944 13240 19950 13252
rect 20088 13240 20116 13271
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 20530 13317 20536 13320
rect 20487 13311 20536 13317
rect 20487 13277 20499 13311
rect 20533 13277 20536 13311
rect 20487 13271 20536 13277
rect 20530 13268 20536 13271
rect 20588 13268 20594 13320
rect 22738 13268 22744 13320
rect 22796 13308 22802 13320
rect 22796 13280 23980 13308
rect 22796 13268 22802 13280
rect 19944 13212 20116 13240
rect 20349 13243 20407 13249
rect 19944 13200 19950 13212
rect 20349 13209 20361 13243
rect 20395 13240 20407 13243
rect 20990 13240 20996 13252
rect 20395 13212 20996 13240
rect 20395 13209 20407 13212
rect 20349 13203 20407 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 21082 13200 21088 13252
rect 21140 13200 21146 13252
rect 22373 13243 22431 13249
rect 22373 13209 22385 13243
rect 22419 13240 22431 13243
rect 23106 13240 23112 13252
rect 22419 13212 23112 13240
rect 22419 13209 22431 13212
rect 22373 13203 22431 13209
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 23569 13243 23627 13249
rect 23569 13209 23581 13243
rect 23615 13240 23627 13243
rect 23842 13240 23848 13252
rect 23615 13212 23848 13240
rect 23615 13209 23627 13212
rect 23569 13203 23627 13209
rect 23842 13200 23848 13212
rect 23900 13200 23906 13252
rect 23952 13240 23980 13280
rect 24026 13268 24032 13320
rect 24084 13308 24090 13320
rect 24578 13308 24584 13320
rect 24084 13280 24584 13308
rect 24084 13268 24090 13280
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 24688 13308 24716 13348
rect 26252 13308 26280 13484
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 24688 13280 26280 13308
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 26694 13317 26700 13320
rect 26688 13308 26700 13317
rect 26655 13280 26700 13308
rect 26688 13271 26700 13280
rect 26694 13268 26700 13271
rect 26752 13268 26758 13320
rect 24848 13243 24906 13249
rect 23952 13212 24799 13240
rect 16022 13172 16028 13184
rect 15948 13144 16028 13172
rect 14737 13135 14795 13141
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16206 13132 16212 13184
rect 16264 13132 16270 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 18230 13172 18236 13184
rect 16816 13144 18236 13172
rect 16816 13132 16822 13144
rect 18230 13132 18236 13144
rect 18288 13172 18294 13184
rect 18785 13175 18843 13181
rect 18785 13172 18797 13175
rect 18288 13144 18797 13172
rect 18288 13132 18294 13144
rect 18785 13141 18797 13144
rect 18831 13141 18843 13175
rect 18785 13135 18843 13141
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 19576 13144 20637 13172
rect 19576 13132 19582 13144
rect 20625 13141 20637 13144
rect 20671 13141 20683 13175
rect 20625 13135 20683 13141
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21285 13175 21343 13181
rect 21285 13172 21297 13175
rect 20772 13144 21297 13172
rect 20772 13132 20778 13144
rect 21285 13141 21297 13144
rect 21331 13141 21343 13175
rect 21285 13135 21343 13141
rect 22833 13175 22891 13181
rect 22833 13141 22845 13175
rect 22879 13172 22891 13175
rect 24670 13172 24676 13184
rect 22879 13144 24676 13172
rect 22879 13141 22891 13144
rect 22833 13135 22891 13141
rect 24670 13132 24676 13144
rect 24728 13132 24734 13184
rect 24771 13172 24799 13212
rect 24848 13209 24860 13243
rect 24894 13240 24906 13243
rect 28074 13240 28080 13252
rect 24894 13212 28080 13240
rect 24894 13209 24906 13212
rect 24848 13203 24906 13209
rect 28074 13200 28080 13212
rect 28132 13200 28138 13252
rect 27801 13175 27859 13181
rect 27801 13172 27813 13175
rect 24771 13144 27813 13172
rect 27801 13141 27813 13144
rect 27847 13141 27859 13175
rect 27801 13135 27859 13141
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 1912 12940 2145 12968
rect 1912 12928 1918 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 3418 12928 3424 12980
rect 3476 12977 3482 12980
rect 3476 12971 3495 12977
rect 3483 12937 3495 12971
rect 3476 12931 3495 12937
rect 3605 12971 3663 12977
rect 3605 12937 3617 12971
rect 3651 12968 3663 12971
rect 4338 12968 4344 12980
rect 3651 12940 4344 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 3476 12928 3482 12931
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5350 12968 5356 12980
rect 5215 12940 5356 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5776 12940 5917 12968
rect 5776 12928 5782 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 7466 12928 7472 12980
rect 7524 12928 7530 12980
rect 8478 12928 8484 12980
rect 8536 12928 8542 12980
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 10318 12968 10324 12980
rect 8996 12940 10324 12968
rect 8996 12928 9002 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10778 12968 10784 12980
rect 10612 12940 10784 12968
rect 2682 12900 2688 12912
rect 2516 12872 2688 12900
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 2516 12841 2544 12872
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 3237 12903 3295 12909
rect 3237 12869 3249 12903
rect 3283 12869 3295 12903
rect 3452 12900 3480 12928
rect 4890 12900 4896 12912
rect 3452 12872 4896 12900
rect 3237 12863 3295 12869
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 2372 12804 2421 12832
rect 2372 12792 2378 12804
rect 2409 12801 2421 12804
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3050 12832 3056 12844
rect 2823 12804 3056 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2608 12764 2636 12795
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3252 12832 3280 12863
rect 4890 12860 4896 12872
rect 4948 12860 4954 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 8386 12900 8392 12912
rect 6328 12872 8392 12900
rect 6328 12860 6334 12872
rect 8386 12860 8392 12872
rect 8444 12900 8450 12912
rect 10612 12909 10640 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11146 12968 11152 12980
rect 11020 12940 11152 12968
rect 11020 12928 11026 12940
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 12069 12971 12127 12977
rect 11664 12940 12020 12968
rect 11664 12928 11670 12940
rect 10597 12903 10655 12909
rect 8444 12872 9076 12900
rect 8444 12860 8450 12872
rect 3602 12832 3608 12844
rect 3252 12804 3608 12832
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4798 12832 4804 12844
rect 4479 12804 4804 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4798 12792 4804 12804
rect 4856 12832 4862 12844
rect 4856 12804 4936 12832
rect 4856 12792 4862 12804
rect 2958 12764 2964 12776
rect 2608 12736 2964 12764
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3292 12736 4200 12764
rect 3292 12724 3298 12736
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 4172 12696 4200 12736
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4525 12767 4583 12773
rect 4525 12764 4537 12767
rect 4304 12736 4537 12764
rect 4304 12724 4310 12736
rect 4525 12733 4537 12736
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 4706 12724 4712 12776
rect 4764 12724 4770 12776
rect 4908 12764 4936 12804
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6822 12832 6828 12844
rect 6604 12804 6828 12832
rect 6604 12792 6610 12804
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 8754 12832 8760 12844
rect 8619 12804 8760 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 5350 12764 5356 12776
rect 4908 12736 5356 12764
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12764 7527 12767
rect 7558 12764 7564 12776
rect 7515 12736 7564 12764
rect 7515 12733 7527 12736
rect 7469 12727 7527 12733
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 8312 12764 8340 12795
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9048 12841 9076 12872
rect 10597 12869 10609 12903
rect 10643 12869 10655 12903
rect 11747 12903 11805 12909
rect 11747 12900 11759 12903
rect 10597 12863 10655 12869
rect 11624 12872 11759 12900
rect 11624 12844 11652 12872
rect 11747 12869 11759 12872
rect 11793 12869 11805 12903
rect 11747 12863 11805 12869
rect 11901 12903 11959 12909
rect 11901 12869 11913 12903
rect 11947 12869 11959 12903
rect 11992 12900 12020 12940
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 13814 12968 13820 12980
rect 12115 12940 13820 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 13998 12968 14004 12980
rect 13955 12940 14004 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14792 12940 15025 12968
rect 14792 12928 14798 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 16540 12940 18337 12968
rect 16540 12928 16546 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 18874 12928 18880 12980
rect 18932 12928 18938 12980
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 19208 12940 19334 12968
rect 19208 12928 19214 12940
rect 12894 12900 12900 12912
rect 11992 12872 12572 12900
rect 11901 12863 11959 12869
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11146 12832 11152 12844
rect 10827 12804 11152 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11606 12792 11612 12844
rect 11664 12792 11670 12844
rect 8662 12764 8668 12776
rect 8312 12736 8668 12764
rect 8662 12724 8668 12736
rect 8720 12764 8726 12776
rect 9858 12764 9864 12776
rect 8720 12736 9864 12764
rect 8720 12724 8726 12736
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 11422 12764 11428 12776
rect 10100 12736 11428 12764
rect 10100 12724 10106 12736
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11916 12764 11944 12863
rect 12544 12841 12572 12872
rect 12636 12872 12900 12900
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12636 12764 12664 12872
rect 12894 12860 12900 12872
rect 12952 12900 12958 12912
rect 14366 12900 14372 12912
rect 12952 12872 14372 12900
rect 12952 12860 12958 12872
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 17129 12903 17187 12909
rect 16356 12872 16989 12900
rect 16356 12860 16362 12872
rect 12802 12841 12808 12844
rect 12796 12795 12808 12841
rect 12802 12792 12808 12795
rect 12860 12792 12866 12844
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14274 12832 14280 12844
rect 13872 12804 14280 12832
rect 13872 12792 13878 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14734 12832 14740 12844
rect 14599 12804 14740 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15160 12804 15485 12832
rect 15160 12792 15166 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 15562 12792 15568 12844
rect 15620 12792 15626 12844
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 16206 12832 16212 12844
rect 15795 12804 16212 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16961 12841 16989 12872
rect 17129 12869 17141 12903
rect 17175 12900 17187 12903
rect 17494 12900 17500 12912
rect 17175 12872 17500 12900
rect 17175 12869 17187 12872
rect 17129 12863 17187 12869
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 17586 12860 17592 12912
rect 17644 12860 17650 12912
rect 17954 12860 17960 12912
rect 18012 12860 18018 12912
rect 18138 12860 18144 12912
rect 18196 12909 18202 12912
rect 18196 12903 18215 12909
rect 18203 12869 18215 12903
rect 19306 12900 19334 12940
rect 19702 12928 19708 12980
rect 19760 12968 19766 12980
rect 19889 12971 19947 12977
rect 19889 12968 19901 12971
rect 19760 12940 19901 12968
rect 19760 12928 19766 12940
rect 19889 12937 19901 12940
rect 19935 12937 19947 12971
rect 19889 12931 19947 12937
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 20714 12968 20720 12980
rect 20128 12940 20720 12968
rect 20128 12928 20134 12940
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 22649 12971 22707 12977
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 24026 12968 24032 12980
rect 22695 12940 24032 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 27982 12968 27988 12980
rect 24136 12940 27988 12968
rect 20806 12900 20812 12912
rect 19306 12872 20812 12900
rect 18196 12863 18215 12869
rect 18196 12860 18202 12863
rect 20806 12860 20812 12872
rect 20864 12860 20870 12912
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 21499 12872 22416 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 16860 12835 16918 12841
rect 16860 12832 16872 12835
rect 16776 12804 16872 12832
rect 11916 12736 12664 12764
rect 5810 12696 5816 12708
rect 3200 12668 3464 12696
rect 4172 12668 5816 12696
rect 3200 12656 3206 12668
rect 3436 12637 3464 12668
rect 5810 12656 5816 12668
rect 5868 12656 5874 12708
rect 5902 12656 5908 12708
rect 5960 12696 5966 12708
rect 6454 12696 6460 12708
rect 5960 12668 6460 12696
rect 5960 12656 5966 12668
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 8260 12668 10149 12696
rect 8260 12656 8266 12668
rect 10137 12665 10149 12668
rect 10183 12665 10195 12699
rect 10137 12659 10195 12665
rect 12176 12640 12204 12736
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 13688 12736 15393 12764
rect 13688 12724 13694 12736
rect 15381 12733 15393 12736
rect 15427 12733 15439 12767
rect 16776 12764 16804 12804
rect 16860 12801 16872 12804
rect 16906 12801 16918 12835
rect 16860 12795 16918 12801
rect 16946 12835 17004 12841
rect 16946 12801 16958 12835
rect 16992 12801 17004 12835
rect 16946 12795 17004 12801
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 17092 12804 17233 12832
rect 17092 12792 17098 12804
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17359 12835 17417 12841
rect 17359 12801 17371 12835
rect 17405 12832 17417 12835
rect 17604 12832 17632 12860
rect 17405 12804 17632 12832
rect 17405 12801 17417 12804
rect 17359 12795 17417 12801
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 19245 12835 19303 12841
rect 19245 12832 19257 12835
rect 17736 12804 19257 12832
rect 17736 12792 17742 12804
rect 19245 12801 19257 12804
rect 19291 12832 19303 12835
rect 19291 12804 20040 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 17586 12764 17592 12776
rect 16776 12736 17592 12764
rect 15381 12727 15439 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 18782 12764 18788 12776
rect 18064 12736 18788 12764
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12696 14427 12699
rect 14415 12668 17816 12696
rect 14415 12665 14427 12668
rect 14369 12659 14427 12665
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12597 3479 12631
rect 3421 12591 3479 12597
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 6362 12628 6368 12640
rect 4120 12600 6368 12628
rect 4120 12588 4126 12600
rect 6362 12588 6368 12600
rect 6420 12628 6426 12640
rect 6730 12628 6736 12640
rect 6420 12600 6736 12628
rect 6420 12588 6426 12600
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7892 12600 8125 12628
rect 7892 12588 7898 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 8846 12628 8852 12640
rect 8444 12600 8852 12628
rect 8444 12588 8450 12600
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 9088 12600 9137 12628
rect 9088 12588 9094 12600
rect 9125 12597 9137 12600
rect 9171 12597 9183 12631
rect 9125 12591 9183 12597
rect 9950 12588 9956 12640
rect 10008 12588 10014 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10284 12600 10977 12628
rect 10284 12588 10290 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11112 12600 11897 12628
rect 11112 12588 11118 12600
rect 11885 12597 11897 12600
rect 11931 12597 11943 12631
rect 11885 12591 11943 12597
rect 12158 12588 12164 12640
rect 12216 12588 12222 12640
rect 15286 12588 15292 12640
rect 15344 12588 15350 12640
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 15804 12600 17509 12628
rect 15804 12588 15810 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 17788 12628 17816 12668
rect 18064 12628 18092 12736
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19058 12724 19064 12776
rect 19116 12724 19122 12776
rect 19150 12724 19156 12776
rect 19208 12724 19214 12776
rect 19334 12724 19340 12776
rect 19392 12724 19398 12776
rect 20012 12764 20040 12804
rect 20070 12792 20076 12844
rect 20128 12792 20134 12844
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20622 12832 20628 12844
rect 20211 12804 20628 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 20732 12804 21281 12832
rect 20254 12764 20260 12776
rect 20012 12736 20260 12764
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12733 20407 12767
rect 20732 12764 20760 12804
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 22278 12792 22284 12844
rect 22336 12792 22342 12844
rect 22388 12832 22416 12872
rect 22554 12860 22560 12912
rect 22612 12900 22618 12912
rect 24136 12900 24164 12940
rect 27982 12928 27988 12940
rect 28040 12928 28046 12980
rect 28074 12928 28080 12980
rect 28132 12928 28138 12980
rect 22612 12872 24164 12900
rect 24305 12903 24363 12909
rect 22612 12860 22618 12872
rect 24305 12869 24317 12903
rect 24351 12900 24363 12903
rect 24578 12900 24584 12912
rect 24351 12872 24584 12900
rect 24351 12869 24363 12872
rect 24305 12863 24363 12869
rect 24578 12860 24584 12872
rect 24636 12900 24642 12912
rect 26418 12900 26424 12912
rect 24636 12872 26424 12900
rect 24636 12860 24642 12872
rect 22462 12832 22468 12844
rect 22388 12804 22468 12832
rect 22462 12792 22468 12804
rect 22520 12832 22526 12844
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 22520 12804 22753 12832
rect 22520 12792 22526 12804
rect 22741 12801 22753 12804
rect 22787 12801 22799 12835
rect 22741 12795 22799 12801
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 23658 12792 23664 12844
rect 23716 12832 23722 12844
rect 25240 12841 25268 12872
rect 26418 12860 26424 12872
rect 26476 12860 26482 12912
rect 27154 12860 27160 12912
rect 27212 12860 27218 12912
rect 24121 12835 24179 12841
rect 24121 12832 24133 12835
rect 23716 12804 24133 12832
rect 23716 12792 23722 12804
rect 24121 12801 24133 12804
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 25314 12792 25320 12844
rect 25372 12832 25378 12844
rect 25481 12835 25539 12841
rect 25481 12832 25493 12835
rect 25372 12804 25493 12832
rect 25372 12792 25378 12804
rect 25481 12801 25493 12804
rect 25527 12801 25539 12835
rect 25481 12795 25539 12801
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 28261 12835 28319 12841
rect 28261 12832 28273 12835
rect 27672 12804 28273 12832
rect 27672 12792 27678 12804
rect 28261 12801 28273 12804
rect 28307 12801 28319 12835
rect 28261 12795 28319 12801
rect 20349 12727 20407 12733
rect 20548 12736 20760 12764
rect 19978 12696 19984 12708
rect 18156 12668 19984 12696
rect 18156 12637 18184 12668
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 20162 12656 20168 12708
rect 20220 12696 20226 12708
rect 20364 12696 20392 12727
rect 20220 12668 20392 12696
rect 20220 12656 20226 12668
rect 17788 12600 18092 12628
rect 18141 12631 18199 12637
rect 17497 12591 17555 12597
rect 18141 12597 18153 12631
rect 18187 12597 18199 12631
rect 18141 12591 18199 12597
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 19150 12628 19156 12640
rect 18656 12600 19156 12628
rect 18656 12588 18662 12600
rect 19150 12588 19156 12600
rect 19208 12628 19214 12640
rect 20548 12628 20576 12736
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21085 12767 21143 12773
rect 21085 12764 21097 12767
rect 20956 12736 21097 12764
rect 20956 12724 20962 12736
rect 21085 12733 21097 12736
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 23385 12699 23443 12705
rect 23385 12665 23397 12699
rect 23431 12696 23443 12699
rect 23474 12696 23480 12708
rect 23431 12668 23480 12696
rect 23431 12665 23443 12668
rect 23385 12659 23443 12665
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 26234 12656 26240 12708
rect 26292 12696 26298 12708
rect 27433 12699 27491 12705
rect 27433 12696 27445 12699
rect 26292 12668 27445 12696
rect 26292 12656 26298 12668
rect 27433 12665 27445 12668
rect 27479 12665 27491 12699
rect 27433 12659 27491 12665
rect 19208 12600 20576 12628
rect 19208 12588 19214 12600
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 20772 12600 22017 12628
rect 20772 12588 20778 12600
rect 22005 12597 22017 12600
rect 22051 12597 22063 12631
rect 22005 12591 22063 12597
rect 22370 12588 22376 12640
rect 22428 12588 22434 12640
rect 22462 12588 22468 12640
rect 22520 12588 22526 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 26605 12631 26663 12637
rect 26605 12628 26617 12631
rect 23348 12600 26617 12628
rect 23348 12588 23354 12600
rect 26605 12597 26617 12600
rect 26651 12597 26663 12631
rect 26605 12591 26663 12597
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27617 12631 27675 12637
rect 27617 12628 27629 12631
rect 26752 12600 27629 12628
rect 26752 12588 26758 12600
rect 27617 12597 27629 12600
rect 27663 12597 27675 12631
rect 27617 12591 27675 12597
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 4246 12424 4252 12436
rect 2363 12396 4252 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 5074 12424 5080 12436
rect 4479 12396 5080 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 3329 12359 3387 12365
rect 3329 12356 3341 12359
rect 2424 12328 3341 12356
rect 2424 12300 2452 12328
rect 3329 12325 3341 12328
rect 3375 12325 3387 12359
rect 3329 12319 3387 12325
rect 2406 12288 2412 12300
rect 1964 12260 2412 12288
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 1780 12084 1808 12183
rect 1964 12164 1992 12260
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3878 12288 3884 12300
rect 3200 12260 3884 12288
rect 3200 12248 3206 12260
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 3936 12260 4660 12288
rect 3936 12248 3942 12260
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 4632 12229 4660 12260
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5736 12288 5764 12387
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6546 12424 6552 12436
rect 6144 12396 6552 12424
rect 6144 12384 6150 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7024 12396 7941 12424
rect 4764 12260 5764 12288
rect 5828 12328 6316 12356
rect 4764 12248 4770 12260
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 1946 12112 1952 12164
rect 2004 12112 2010 12164
rect 2041 12155 2099 12161
rect 2041 12121 2053 12155
rect 2087 12152 2099 12155
rect 2222 12152 2228 12164
rect 2087 12124 2228 12152
rect 2087 12121 2099 12124
rect 2041 12115 2099 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 3252 12152 3280 12183
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5074 12220 5080 12232
rect 4939 12192 5080 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5828 12220 5856 12328
rect 5460 12192 5856 12220
rect 5460 12152 5488 12192
rect 3252 12124 5488 12152
rect 5537 12155 5595 12161
rect 5537 12121 5549 12155
rect 5583 12121 5595 12155
rect 5537 12115 5595 12121
rect 3234 12084 3240 12096
rect 1780 12056 3240 12084
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 5552 12084 5580 12115
rect 4396 12056 5580 12084
rect 5747 12087 5805 12093
rect 4396 12044 4402 12056
rect 5747 12053 5759 12087
rect 5793 12084 5805 12087
rect 5902 12084 5908 12096
rect 5793 12056 5908 12084
rect 5793 12053 5805 12056
rect 5747 12047 5805 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6288 12084 6316 12328
rect 6454 12288 6460 12300
rect 6380 12260 6460 12288
rect 6380 12229 6408 12260
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 6822 12288 6828 12300
rect 6564 12260 6828 12288
rect 6564 12229 6592 12260
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7024 12229 7052 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10192 12396 10701 12424
rect 10192 12384 10198 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11204 12396 12480 12424
rect 11204 12384 11210 12396
rect 7282 12316 7288 12368
rect 7340 12316 7346 12368
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 8110 12356 8116 12368
rect 7708 12328 8116 12356
rect 7708 12316 7714 12328
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8202 12316 8208 12368
rect 8260 12316 8266 12368
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12356 8355 12359
rect 8386 12356 8392 12368
rect 8343 12328 8392 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 11054 12356 11060 12368
rect 10376 12328 11060 12356
rect 10376 12316 10382 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 12342 12316 12348 12368
rect 12400 12316 12406 12368
rect 12452 12356 12480 12396
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12860 12396 13001 12424
rect 12860 12384 12866 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14516 12396 14933 12424
rect 14516 12384 14522 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 14921 12387 14979 12393
rect 15028 12396 15945 12424
rect 14182 12356 14188 12368
rect 12452 12328 14188 12356
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 15028 12356 15056 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 15933 12387 15991 12393
rect 16666 12384 16672 12436
rect 16724 12384 16730 12436
rect 16850 12384 16856 12436
rect 16908 12384 16914 12436
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 18138 12424 18144 12436
rect 17788 12396 18144 12424
rect 14292 12328 15056 12356
rect 9214 12288 9220 12300
rect 8128 12260 9220 12288
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6696 12192 7021 12220
rect 6696 12180 6702 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7834 12220 7840 12232
rect 7340 12192 7840 12220
rect 7340 12180 7346 12192
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8128 12229 8156 12260
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 10042 12288 10048 12300
rect 9324 12260 10048 12288
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8570 12180 8576 12232
rect 8628 12180 8634 12232
rect 9324 12229 9352 12260
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 10428 12260 10609 12288
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10226 12220 10232 12232
rect 9907 12192 10232 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10428 12164 10456 12260
rect 10597 12257 10609 12260
rect 10643 12257 10655 12291
rect 10597 12251 10655 12257
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 14292 12232 14320 12328
rect 15102 12316 15108 12368
rect 15160 12316 15166 12368
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 16448 12328 17693 12356
rect 16448 12316 16454 12328
rect 17681 12325 17693 12328
rect 17727 12325 17739 12359
rect 17681 12319 17739 12325
rect 17788 12288 17816 12396
rect 18138 12384 18144 12396
rect 18196 12424 18202 12436
rect 18322 12424 18328 12436
rect 18196 12396 18328 12424
rect 18196 12384 18202 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 18506 12424 18512 12436
rect 18463 12396 18512 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 18601 12427 18659 12433
rect 18601 12393 18613 12427
rect 18647 12424 18659 12427
rect 19426 12424 19432 12436
rect 18647 12396 19432 12424
rect 18647 12393 18659 12396
rect 18601 12387 18659 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 19702 12424 19708 12436
rect 19659 12396 19708 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 22094 12424 22100 12436
rect 19944 12396 22100 12424
rect 19944 12384 19950 12396
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 23842 12424 23848 12436
rect 23532 12396 23848 12424
rect 23532 12384 23538 12396
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 25038 12384 25044 12436
rect 25096 12424 25102 12436
rect 28353 12427 28411 12433
rect 28353 12424 28365 12427
rect 25096 12396 28365 12424
rect 25096 12384 25102 12396
rect 28353 12393 28365 12396
rect 28399 12393 28411 12427
rect 28353 12387 28411 12393
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 19978 12356 19984 12368
rect 18288 12328 19984 12356
rect 18288 12316 18294 12328
rect 19978 12316 19984 12328
rect 20036 12356 20042 12368
rect 20898 12356 20904 12368
rect 20036 12328 20904 12356
rect 20036 12316 20042 12328
rect 20898 12316 20904 12328
rect 20956 12316 20962 12368
rect 21542 12316 21548 12368
rect 21600 12356 21606 12368
rect 21729 12359 21787 12365
rect 21729 12356 21741 12359
rect 21600 12328 21741 12356
rect 21600 12316 21606 12328
rect 21729 12325 21741 12328
rect 21775 12325 21787 12359
rect 21729 12319 21787 12325
rect 22741 12359 22799 12365
rect 22741 12325 22753 12359
rect 22787 12356 22799 12359
rect 22922 12356 22928 12368
rect 22787 12328 22928 12356
rect 22787 12325 22799 12328
rect 22741 12319 22799 12325
rect 22922 12316 22928 12328
rect 22980 12356 22986 12368
rect 23382 12356 23388 12368
rect 22980 12328 23388 12356
rect 22980 12316 22986 12328
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 23661 12359 23719 12365
rect 23661 12325 23673 12359
rect 23707 12356 23719 12359
rect 23750 12356 23756 12368
rect 23707 12328 23756 12356
rect 23707 12325 23719 12328
rect 23661 12319 23719 12325
rect 23750 12316 23756 12328
rect 23808 12316 23814 12368
rect 15120 12260 16528 12288
rect 15120 12232 15148 12260
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10686 12222 10692 12232
rect 10612 12220 10692 12222
rect 10551 12194 10692 12220
rect 10551 12192 10640 12194
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10686 12180 10692 12194
rect 10744 12180 10750 12232
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 10928 12192 11437 12220
rect 10928 12180 10934 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 11425 12183 11483 12189
rect 11532 12192 13185 12220
rect 6457 12155 6515 12161
rect 6457 12121 6469 12155
rect 6503 12152 6515 12155
rect 8294 12152 8300 12164
rect 6503 12124 8300 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 8294 12112 8300 12124
rect 8352 12112 8358 12164
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 10045 12155 10103 12161
rect 10045 12152 10057 12155
rect 9640 12124 10057 12152
rect 9640 12112 9646 12124
rect 10045 12121 10057 12124
rect 10091 12152 10103 12155
rect 10410 12152 10416 12164
rect 10091 12124 10416 12152
rect 10091 12121 10103 12124
rect 10045 12115 10103 12121
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 11532 12152 11560 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14424 12195 14996 12220
rect 14424 12192 15025 12195
rect 14424 12180 14430 12192
rect 14967 12189 15025 12192
rect 10836 12124 11560 12152
rect 10836 12112 10842 12124
rect 12066 12112 12072 12164
rect 12124 12152 12130 12164
rect 13446 12152 13452 12164
rect 12124 12124 13452 12152
rect 12124 12112 12130 12124
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 14737 12155 14795 12161
rect 14737 12121 14749 12155
rect 14783 12152 14795 12155
rect 14826 12152 14832 12164
rect 14783 12124 14832 12152
rect 14783 12121 14795 12124
rect 14737 12115 14795 12121
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 14967 12155 14979 12189
rect 15013 12155 15025 12189
rect 15102 12180 15108 12232
rect 15160 12180 15166 12232
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15712 12192 15761 12220
rect 15712 12180 15718 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 14967 12149 15025 12155
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15672 12152 15700 12180
rect 16500 12164 16528 12260
rect 16776 12260 17816 12288
rect 15252 12124 15700 12152
rect 15252 12112 15258 12124
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 16690 12155 16748 12161
rect 16690 12121 16702 12155
rect 16736 12152 16748 12155
rect 16776 12152 16804 12260
rect 18322 12248 18328 12300
rect 18380 12288 18386 12300
rect 20070 12288 20076 12300
rect 18380 12260 20076 12288
rect 18380 12248 18386 12260
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 21450 12288 21456 12300
rect 20824 12260 21456 12288
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 20714 12220 20720 12232
rect 16908 12192 20720 12220
rect 16908 12180 16914 12192
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 20824 12229 20852 12260
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 21913 12291 21971 12297
rect 21913 12257 21925 12291
rect 21959 12288 21971 12291
rect 23566 12288 23572 12300
rect 21959 12260 23572 12288
rect 21959 12257 21971 12260
rect 21913 12251 21971 12257
rect 23566 12248 23572 12260
rect 23624 12248 23630 12300
rect 26326 12288 26332 12300
rect 23768 12260 26332 12288
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12220 21051 12223
rect 22278 12220 22284 12232
rect 21039 12192 22284 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 23474 12220 23480 12232
rect 22388 12192 23480 12220
rect 16736 12124 16804 12152
rect 16736 12121 16748 12124
rect 16690 12115 16748 12121
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17313 12155 17371 12161
rect 17313 12152 17325 12155
rect 17000 12124 17325 12152
rect 17000 12112 17006 12124
rect 17313 12121 17325 12124
rect 17359 12152 17371 12155
rect 17954 12152 17960 12164
rect 17359 12124 17960 12152
rect 17359 12121 17371 12124
rect 17313 12115 17371 12121
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 18230 12112 18236 12164
rect 18288 12112 18294 12164
rect 19058 12152 19064 12164
rect 18356 12124 19064 12152
rect 8938 12084 8944 12096
rect 6288 12056 8944 12084
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9122 12044 9128 12096
rect 9180 12044 9186 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10870 12084 10876 12096
rect 9916 12056 10876 12084
rect 9916 12044 9922 12056
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12529 12087 12587 12093
rect 12529 12084 12541 12087
rect 11848 12056 12541 12084
rect 11848 12044 11854 12056
rect 12529 12053 12541 12056
rect 12575 12053 12587 12087
rect 12529 12047 12587 12053
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 15838 12084 15844 12096
rect 13136 12056 15844 12084
rect 13136 12044 13142 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17513 12087 17571 12093
rect 17513 12084 17525 12087
rect 16632 12056 17525 12084
rect 16632 12044 16638 12056
rect 17513 12053 17525 12056
rect 17559 12084 17571 12087
rect 18138 12084 18144 12096
rect 17559 12056 18144 12084
rect 17559 12053 17571 12056
rect 17513 12047 17571 12053
rect 18138 12044 18144 12056
rect 18196 12084 18202 12096
rect 18356 12084 18384 12124
rect 19058 12112 19064 12124
rect 19116 12152 19122 12164
rect 19116 12124 19334 12152
rect 19116 12112 19122 12124
rect 18196 12056 18384 12084
rect 18433 12087 18491 12093
rect 18196 12044 18202 12056
rect 18433 12053 18445 12087
rect 18479 12084 18491 12087
rect 18690 12084 18696 12096
rect 18479 12056 18696 12084
rect 18479 12053 18491 12056
rect 18433 12047 18491 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 19306 12084 19334 12124
rect 19426 12112 19432 12164
rect 19484 12152 19490 12164
rect 19978 12152 19984 12164
rect 19484 12124 19984 12152
rect 19484 12112 19490 12124
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20625 12155 20683 12161
rect 20625 12121 20637 12155
rect 20671 12152 20683 12155
rect 20898 12152 20904 12164
rect 20671 12124 20904 12152
rect 20671 12121 20683 12124
rect 20625 12115 20683 12121
rect 20898 12112 20904 12124
rect 20956 12112 20962 12164
rect 21358 12112 21364 12164
rect 21416 12152 21422 12164
rect 22388 12161 22416 12192
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 21453 12155 21511 12161
rect 21453 12152 21465 12155
rect 21416 12124 21465 12152
rect 21416 12112 21422 12124
rect 21453 12121 21465 12124
rect 21499 12152 21511 12155
rect 22373 12155 22431 12161
rect 22373 12152 22385 12155
rect 21499 12124 22385 12152
rect 21499 12121 21511 12124
rect 21453 12115 21511 12121
rect 22373 12121 22385 12124
rect 22419 12121 22431 12155
rect 22373 12115 22431 12121
rect 22462 12112 22468 12164
rect 22520 12152 22526 12164
rect 23014 12152 23020 12164
rect 22520 12124 23020 12152
rect 22520 12112 22526 12124
rect 23014 12112 23020 12124
rect 23072 12152 23078 12164
rect 23293 12155 23351 12161
rect 23293 12152 23305 12155
rect 23072 12124 23305 12152
rect 23072 12112 23078 12124
rect 23293 12121 23305 12124
rect 23339 12121 23351 12155
rect 23293 12115 23351 12121
rect 19629 12087 19687 12093
rect 19629 12084 19641 12087
rect 19306 12056 19641 12084
rect 19629 12053 19641 12056
rect 19675 12053 19687 12087
rect 19629 12047 19687 12053
rect 19794 12044 19800 12096
rect 19852 12044 19858 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20530 12084 20536 12096
rect 20220 12056 20536 12084
rect 20220 12044 20226 12056
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12084 22891 12087
rect 23198 12084 23204 12096
rect 22879 12056 23204 12084
rect 22879 12053 22891 12056
rect 22833 12047 22891 12053
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 23768 12093 23796 12260
rect 26326 12248 26332 12260
rect 26384 12248 26390 12300
rect 26418 12248 26424 12300
rect 26476 12288 26482 12300
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 26476 12260 26985 12288
rect 26476 12248 26482 12260
rect 26973 12257 26985 12260
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24728 12192 24777 12220
rect 24728 12180 24734 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 27218 12155 27276 12161
rect 27218 12152 27230 12155
rect 24596 12124 27230 12152
rect 24596 12093 24624 12124
rect 27218 12121 27230 12124
rect 27264 12121 27276 12155
rect 27218 12115 27276 12121
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12053 23811 12087
rect 23753 12047 23811 12053
rect 24581 12087 24639 12093
rect 24581 12053 24593 12087
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 382 11840 388 11892
rect 440 11880 446 11892
rect 934 11880 940 11892
rect 440 11852 940 11880
rect 440 11840 446 11852
rect 934 11840 940 11852
rect 992 11840 998 11892
rect 2958 11840 2964 11892
rect 3016 11840 3022 11892
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3510 11880 3516 11892
rect 3108 11852 3516 11880
rect 3108 11840 3114 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3789 11883 3847 11889
rect 3789 11849 3801 11883
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 1762 11772 1768 11824
rect 1820 11772 1826 11824
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 3804 11812 3832 11843
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 3936 11852 4629 11880
rect 3936 11840 3942 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5537 11883 5595 11889
rect 4764 11852 5488 11880
rect 4764 11840 4770 11852
rect 2188 11784 3832 11812
rect 2188 11772 2194 11784
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 5460 11812 5488 11852
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 8662 11880 8668 11892
rect 5583 11852 8668 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9674 11880 9680 11892
rect 8772 11852 9680 11880
rect 4212 11784 5396 11812
rect 5460 11784 5580 11812
rect 4212 11772 4218 11784
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1118 11744 1124 11756
rect 992 11716 1124 11744
rect 992 11704 998 11716
rect 1118 11704 1124 11716
rect 1176 11704 1182 11756
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2406 11744 2412 11756
rect 1995 11716 2412 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 658 11636 664 11688
rect 716 11676 722 11688
rect 1210 11676 1216 11688
rect 716 11648 1216 11676
rect 716 11636 722 11648
rect 1210 11636 1216 11648
rect 1268 11636 1274 11688
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2608 11676 2636 11707
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3568 11716 3709 11744
rect 3568 11704 3574 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11744 4675 11747
rect 4706 11744 4712 11756
rect 4663 11716 4712 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 2096 11648 2636 11676
rect 2096 11636 2102 11648
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3896 11676 3924 11707
rect 3016 11648 3924 11676
rect 3988 11676 4016 11707
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 5368 11753 5396 11784
rect 5552 11756 5580 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8113 11815 8171 11821
rect 8113 11812 8125 11815
rect 7708 11784 8125 11812
rect 7708 11772 7714 11784
rect 8113 11781 8125 11784
rect 8159 11781 8171 11815
rect 8113 11775 8171 11781
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 8772 11812 8800 11852
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 12066 11880 12072 11892
rect 10060 11852 12072 11880
rect 10060 11812 10088 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 12308 11852 13093 11880
rect 12308 11840 12314 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 13633 11883 13691 11889
rect 13633 11849 13645 11883
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 8536 11784 8800 11812
rect 9048 11784 10088 11812
rect 8536 11772 8542 11784
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 5534 11704 5540 11756
rect 5592 11704 5598 11756
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6512 11716 6653 11744
rect 6512 11704 6518 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6880 11716 6929 11744
rect 6880 11704 6886 11716
rect 6917 11713 6929 11716
rect 6963 11744 6975 11747
rect 7282 11744 7288 11756
rect 6963 11716 7288 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7742 11704 7748 11756
rect 7800 11704 7806 11756
rect 8938 11704 8944 11756
rect 8996 11704 9002 11756
rect 9048 11753 9076 11784
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 10060 11753 10088 11784
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11957 11815 12015 11821
rect 11957 11812 11969 11815
rect 11296 11784 11969 11812
rect 11296 11772 11302 11784
rect 11957 11781 11969 11784
rect 12003 11781 12015 11815
rect 13648 11812 13676 11843
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15528 11852 15577 11880
rect 15528 11840 15534 11852
rect 15565 11849 15577 11852
rect 15611 11849 15623 11883
rect 15565 11843 15623 11849
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 16540 11852 17172 11880
rect 16540 11840 16546 11852
rect 14090 11812 14096 11824
rect 11957 11775 12015 11781
rect 12084 11784 13676 11812
rect 13832 11784 14096 11812
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9692 11716 9781 11744
rect 4062 11676 4068 11688
rect 3988 11648 4068 11676
rect 3016 11636 3022 11648
rect 4062 11636 4068 11648
rect 4120 11676 4126 11688
rect 5184 11676 5212 11704
rect 4120 11648 5212 11676
rect 6733 11679 6791 11685
rect 4120 11636 4126 11648
rect 6733 11645 6745 11679
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 1118 11568 1124 11620
rect 1176 11608 1182 11620
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 1176 11580 5181 11608
rect 1176 11568 1182 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5169 11571 5227 11577
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 6748 11608 6776 11639
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7929 11679 7987 11685
rect 7064 11648 7880 11676
rect 7064 11636 7070 11648
rect 7852 11620 7880 11648
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 8956 11676 8984 11704
rect 9692 11676 9720 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10410 11744 10416 11756
rect 10367 11716 10416 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 8956 11648 9720 11676
rect 7929 11639 7987 11645
rect 6696 11580 6776 11608
rect 6932 11580 7696 11608
rect 6696 11568 6702 11580
rect 1210 11500 1216 11552
rect 1268 11540 1274 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 1268 11512 2145 11540
rect 1268 11500 1274 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2133 11503 2191 11509
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3602 11540 3608 11552
rect 2924 11512 3608 11540
rect 2924 11500 2930 11512
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 6546 11540 6552 11552
rect 3752 11512 6552 11540
rect 3752 11500 3758 11512
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 6932 11549 6960 11580
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11509 6975 11543
rect 6917 11503 6975 11509
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7466 11540 7472 11552
rect 7147 11512 7472 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7668 11540 7696 11580
rect 7834 11568 7840 11620
rect 7892 11568 7898 11620
rect 7944 11608 7972 11639
rect 10134 11636 10140 11688
rect 10192 11636 10198 11688
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10520 11676 10548 11707
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11664 11716 11713 11744
rect 11664 11704 11670 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 12084 11744 12112 11784
rect 11701 11707 11759 11713
rect 11808 11716 12112 11744
rect 11808 11676 11836 11716
rect 13630 11704 13636 11756
rect 13688 11704 13694 11756
rect 13832 11753 13860 11784
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 14366 11812 14372 11824
rect 14240 11784 14372 11812
rect 14240 11772 14246 11784
rect 14366 11772 14372 11784
rect 14424 11812 14430 11824
rect 15105 11815 15163 11821
rect 15105 11812 15117 11815
rect 14424 11784 15117 11812
rect 14424 11772 14430 11784
rect 15105 11781 15117 11784
rect 15151 11812 15163 11815
rect 15378 11812 15384 11824
rect 15151 11784 15384 11812
rect 15151 11781 15163 11784
rect 15105 11775 15163 11781
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 17144 11821 17172 11852
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18690 11880 18696 11892
rect 18012 11852 18696 11880
rect 18012 11840 18018 11852
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 18877 11883 18935 11889
rect 18877 11849 18889 11883
rect 18923 11880 18935 11883
rect 18966 11880 18972 11892
rect 18923 11852 18972 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 20254 11880 20260 11892
rect 19475 11852 20260 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 20346 11840 20352 11892
rect 20404 11880 20410 11892
rect 21634 11880 21640 11892
rect 20404 11852 21640 11880
rect 20404 11840 20410 11852
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25041 11883 25099 11889
rect 25041 11880 25053 11883
rect 24912 11852 25053 11880
rect 24912 11840 24918 11852
rect 25041 11849 25053 11852
rect 25087 11849 25099 11883
rect 25041 11843 25099 11849
rect 27893 11883 27951 11889
rect 27893 11849 27905 11883
rect 27939 11880 27951 11883
rect 28258 11880 28264 11892
rect 27939 11852 28264 11880
rect 27939 11849 27951 11852
rect 27893 11843 27951 11849
rect 28258 11840 28264 11852
rect 28316 11840 28322 11892
rect 17129 11815 17187 11821
rect 17129 11781 17141 11815
rect 17175 11781 17187 11815
rect 17129 11775 17187 11781
rect 17345 11815 17403 11821
rect 17345 11781 17357 11815
rect 17391 11812 17403 11815
rect 19242 11812 19248 11824
rect 17391 11784 19248 11812
rect 17391 11781 17403 11784
rect 17345 11775 17403 11781
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20714 11812 20720 11824
rect 20220 11784 20720 11812
rect 20220 11772 20226 11784
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 26234 11812 26240 11824
rect 21600 11784 26240 11812
rect 21600 11772 21606 11784
rect 26234 11772 26240 11784
rect 26292 11772 26298 11824
rect 27433 11815 27491 11821
rect 27433 11781 27445 11815
rect 27479 11812 27491 11815
rect 27522 11812 27528 11824
rect 27479 11784 27528 11812
rect 27479 11781 27491 11784
rect 27433 11775 27491 11781
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11744 14335 11747
rect 14826 11744 14832 11756
rect 14323 11716 14832 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 14918 11704 14924 11756
rect 14976 11744 14982 11756
rect 15562 11744 15568 11756
rect 14976 11716 15568 11744
rect 14976 11704 14982 11716
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15672 11716 15945 11744
rect 10284 11648 10548 11676
rect 11723 11648 11836 11676
rect 10284 11636 10290 11648
rect 8202 11608 8208 11620
rect 7944 11580 8208 11608
rect 8202 11568 8208 11580
rect 8260 11608 8266 11620
rect 11723 11608 11751 11648
rect 8260 11580 9812 11608
rect 8260 11568 8266 11580
rect 8294 11540 8300 11552
rect 7668 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11540 8358 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8352 11512 8769 11540
rect 8352 11500 8358 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8996 11512 9229 11540
rect 8996 11500 9002 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9784 11540 9812 11580
rect 9876 11580 11751 11608
rect 9876 11540 9904 11580
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 13688 11580 15240 11608
rect 13688 11568 13694 11580
rect 9784 11512 9904 11540
rect 9217 11503 9275 11509
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 13906 11540 13912 11552
rect 10284 11512 13912 11540
rect 10284 11500 10290 11512
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 15212 11540 15240 11580
rect 15378 11568 15384 11620
rect 15436 11608 15442 11620
rect 15672 11608 15700 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16758 11744 16764 11756
rect 16347 11716 16764 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16132 11676 16160 11707
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 17552 11716 18705 11744
rect 17552 11704 17558 11716
rect 18693 11713 18705 11716
rect 18739 11744 18751 11747
rect 19058 11744 19064 11756
rect 18739 11716 19064 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 19794 11744 19800 11756
rect 19659 11716 19800 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20329 11747 20387 11753
rect 20329 11744 20341 11747
rect 19904 11716 20341 11744
rect 18230 11676 18236 11688
rect 16132 11648 18236 11676
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18472 11648 18521 11676
rect 18472 11636 18478 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 19904 11676 19932 11716
rect 20329 11713 20341 11716
rect 20375 11713 20387 11747
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 20329 11707 20387 11713
rect 21928 11716 22109 11744
rect 18509 11639 18567 11645
rect 19352 11648 19932 11676
rect 15436 11580 15700 11608
rect 15841 11611 15899 11617
rect 15436 11568 15442 11580
rect 15841 11577 15853 11611
rect 15887 11608 15899 11611
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 15887 11580 17509 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 19352 11608 19380 11648
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 20036 11648 20085 11676
rect 20036 11636 20042 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 19886 11608 19892 11620
rect 18840 11580 19380 11608
rect 19444 11580 19892 11608
rect 18840 11568 18846 11580
rect 16025 11543 16083 11549
rect 16025 11540 16037 11543
rect 15212 11512 16037 11540
rect 16025 11509 16037 11512
rect 16071 11540 16083 11543
rect 16206 11540 16212 11552
rect 16071 11512 16212 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 19444 11540 19472 11580
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 21174 11568 21180 11620
rect 21232 11608 21238 11620
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 21232 11580 21465 11608
rect 21232 11568 21238 11580
rect 21453 11577 21465 11580
rect 21499 11577 21511 11611
rect 21453 11571 21511 11577
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 21928 11608 21956 11716
rect 22097 11713 22109 11716
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 23917 11747 23975 11753
rect 23917 11744 23929 11747
rect 23308 11716 23929 11744
rect 22002 11636 22008 11688
rect 22060 11676 22066 11688
rect 23308 11676 23336 11716
rect 23917 11713 23929 11716
rect 23963 11713 23975 11747
rect 23917 11707 23975 11713
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11744 26663 11747
rect 26694 11744 26700 11756
rect 26651 11716 26700 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 22060 11648 23336 11676
rect 22060 11636 22066 11648
rect 23658 11636 23664 11688
rect 23716 11636 23722 11688
rect 23106 11608 23112 11620
rect 21600 11580 23112 11608
rect 21600 11568 21606 11580
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 24670 11568 24676 11620
rect 24728 11608 24734 11620
rect 24728 11580 25268 11608
rect 24728 11568 24734 11580
rect 17359 11512 19472 11540
rect 22189 11543 22247 11549
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 22189 11509 22201 11543
rect 22235 11540 22247 11543
rect 22462 11540 22468 11552
rect 22235 11512 22468 11540
rect 22235 11509 22247 11512
rect 22189 11503 22247 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 23017 11543 23075 11549
rect 23017 11509 23029 11543
rect 23063 11540 23075 11543
rect 25130 11540 25136 11552
rect 23063 11512 25136 11540
rect 23063 11509 23075 11512
rect 23017 11503 23075 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 25240 11540 25268 11580
rect 27706 11568 27712 11620
rect 27764 11568 27770 11620
rect 26421 11543 26479 11549
rect 26421 11540 26433 11543
rect 25240 11512 26433 11540
rect 26421 11509 26433 11512
rect 26467 11509 26479 11543
rect 26421 11503 26479 11509
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 3970 11296 3976 11348
rect 4028 11296 4034 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 4948 11308 5549 11336
rect 4948 11296 4954 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 5718 11296 5724 11348
rect 5776 11296 5782 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 9950 11336 9956 11348
rect 7340 11308 9956 11336
rect 7340 11296 7346 11308
rect 3145 11271 3203 11277
rect 3145 11237 3157 11271
rect 3191 11268 3203 11271
rect 3234 11268 3240 11280
rect 3191 11240 3240 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 5169 11271 5227 11277
rect 3476 11240 4476 11268
rect 3476 11228 3482 11240
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 2225 11203 2283 11209
rect 1912 11172 1992 11200
rect 1912 11160 1918 11172
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 1964 11141 1992 11172
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 4246 11200 4252 11212
rect 2271 11172 4252 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 1995 11104 2639 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 1854 11024 1860 11076
rect 1912 11024 1918 11076
rect 2087 11067 2145 11073
rect 2087 11033 2099 11067
rect 2133 11064 2145 11067
rect 2314 11064 2320 11076
rect 2133 11036 2320 11064
rect 2133 11033 2145 11036
rect 2087 11027 2145 11033
rect 2314 11024 2320 11036
rect 2372 11024 2378 11076
rect 2611 11064 2639 11104
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 2866 11064 2872 11076
rect 2611 11036 2872 11064
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10996 1639 10999
rect 2958 10996 2964 11008
rect 1627 10968 2964 10996
rect 1627 10965 1639 10968
rect 1581 10959 1639 10965
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3252 10996 3280 11095
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4172 11064 4200 11095
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4448 11141 4476 11240
rect 5169 11237 5181 11271
rect 5215 11268 5227 11271
rect 5258 11268 5264 11280
rect 5215 11240 5264 11268
rect 5215 11237 5227 11240
rect 5169 11231 5227 11237
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 6181 11271 6239 11277
rect 6181 11237 6193 11271
rect 6227 11237 6239 11271
rect 6181 11231 6239 11237
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 6196 11200 6224 11231
rect 6454 11228 6460 11280
rect 6512 11268 6518 11280
rect 6917 11271 6975 11277
rect 6917 11268 6929 11271
rect 6512 11240 6929 11268
rect 6512 11228 6518 11240
rect 6917 11237 6929 11240
rect 6963 11237 6975 11271
rect 6917 11231 6975 11237
rect 7558 11228 7564 11280
rect 7616 11268 7622 11280
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 7616 11240 7849 11268
rect 7616 11228 7622 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 5868 11172 6224 11200
rect 5868 11160 5874 11172
rect 6270 11160 6276 11212
rect 6328 11160 6334 11212
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 6604 11172 7052 11200
rect 6604 11160 6610 11172
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 4890 11132 4896 11144
rect 4479 11104 4896 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 6288 11132 6316 11160
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 5316 11104 6469 11132
rect 5316 11092 5322 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6457 11095 6515 11101
rect 6564 11104 6929 11132
rect 6564 11076 6592 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 3528 11036 4200 11064
rect 3528 10996 3556 11036
rect 4172 11008 4200 11036
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 5500 11036 5549 11064
rect 5500 11024 5506 11036
rect 5537 11033 5549 11036
rect 5583 11033 5595 11067
rect 5537 11027 5595 11033
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 6086 11064 6092 11076
rect 5684 11036 6092 11064
rect 5684 11024 5690 11036
rect 6086 11024 6092 11036
rect 6144 11064 6150 11076
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 6144 11036 6193 11064
rect 6144 11024 6150 11036
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6181 11027 6239 11033
rect 6546 11024 6552 11076
rect 6604 11024 6610 11076
rect 3252 10968 3556 10996
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 5902 10996 5908 11008
rect 4488 10968 5908 10996
rect 4488 10956 4494 10968
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 6052 10968 6377 10996
rect 6052 10956 6058 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6932 10996 6960 11095
rect 7024 11064 7052 11172
rect 8294 11160 8300 11212
rect 8352 11160 8358 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 8588 11200 8616 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 10505 11339 10563 11345
rect 10505 11305 10517 11339
rect 10551 11336 10563 11339
rect 10870 11336 10876 11348
rect 10551 11308 10876 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11882 11296 11888 11348
rect 11940 11296 11946 11348
rect 12618 11336 12624 11348
rect 11992 11308 12624 11336
rect 9769 11271 9827 11277
rect 9769 11237 9781 11271
rect 9815 11268 9827 11271
rect 11992 11268 12020 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 13262 11296 13268 11348
rect 13320 11296 13326 11348
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13412 11308 13645 11336
rect 13412 11296 13418 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14918 11336 14924 11348
rect 13964 11308 14924 11336
rect 13964 11296 13970 11308
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15381 11339 15439 11345
rect 15381 11305 15393 11339
rect 15427 11336 15439 11339
rect 15470 11336 15476 11348
rect 15427 11308 15476 11336
rect 15427 11305 15439 11308
rect 15381 11299 15439 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 15930 11336 15936 11348
rect 15611 11308 15936 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16209 11339 16267 11345
rect 16209 11305 16221 11339
rect 16255 11336 16267 11339
rect 16666 11336 16672 11348
rect 16255 11308 16672 11336
rect 16255 11305 16267 11308
rect 16209 11299 16267 11305
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 16853 11339 16911 11345
rect 16853 11305 16865 11339
rect 16899 11305 16911 11339
rect 16853 11299 16911 11305
rect 9815 11240 12020 11268
rect 12253 11271 12311 11277
rect 9815 11237 9827 11240
rect 9769 11231 9827 11237
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12526 11268 12532 11280
rect 12299 11240 12532 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 12636 11240 14657 11268
rect 8527 11172 8616 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 10597 11203 10655 11209
rect 8720 11172 10364 11200
rect 8720 11160 8726 11172
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 10226 11132 10232 11144
rect 7147 11104 10232 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10336 11141 10364 11172
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 8205 11067 8263 11073
rect 8205 11064 8217 11067
rect 7024 11036 8217 11064
rect 8205 11033 8217 11036
rect 8251 11033 8263 11067
rect 8205 11027 8263 11033
rect 9398 11024 9404 11076
rect 9456 11024 9462 11076
rect 10612 11064 10640 11163
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 12032 11172 12173 11200
rect 12032 11160 12038 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12636 11200 12664 11240
rect 14645 11237 14657 11240
rect 14691 11268 14703 11271
rect 15654 11268 15660 11280
rect 14691 11240 15660 11268
rect 14691 11237 14703 11240
rect 14645 11231 14703 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 16393 11271 16451 11277
rect 16393 11268 16405 11271
rect 15896 11240 16405 11268
rect 15896 11228 15902 11240
rect 16393 11237 16405 11240
rect 16439 11237 16451 11271
rect 16393 11231 16451 11237
rect 12161 11163 12219 11169
rect 12452 11172 12664 11200
rect 13357 11203 13415 11209
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 11790 11132 11796 11144
rect 11471 11104 11796 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12452 11141 12480 11172
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13538 11200 13544 11212
rect 13403 11172 13544 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14734 11160 14740 11212
rect 14792 11160 14798 11212
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 16868 11200 16896 11299
rect 17310 11296 17316 11348
rect 17368 11296 17374 11348
rect 20162 11336 20168 11348
rect 18708 11308 20168 11336
rect 18230 11228 18236 11280
rect 18288 11268 18294 11280
rect 18708 11277 18736 11308
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20441 11339 20499 11345
rect 20441 11305 20453 11339
rect 20487 11336 20499 11339
rect 20487 11308 20760 11336
rect 20487 11305 20499 11308
rect 20441 11299 20499 11305
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 18288 11240 18705 11268
rect 18288 11228 18294 11240
rect 18693 11237 18705 11240
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 20625 11271 20683 11277
rect 20625 11268 20637 11271
rect 19392 11240 20637 11268
rect 19392 11228 19398 11240
rect 20625 11237 20637 11240
rect 20671 11237 20683 11271
rect 20732 11268 20760 11308
rect 24026 11296 24032 11348
rect 24084 11296 24090 11348
rect 26234 11296 26240 11348
rect 26292 11296 26298 11348
rect 21634 11268 21640 11280
rect 20732 11240 21640 11268
rect 20625 11231 20683 11237
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 22002 11228 22008 11280
rect 22060 11228 22066 11280
rect 22554 11228 22560 11280
rect 22612 11268 22618 11280
rect 22612 11240 22692 11268
rect 22612 11228 22618 11240
rect 14884 11172 16896 11200
rect 17037 11203 17095 11209
rect 14884 11160 14890 11172
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 17494 11200 17500 11212
rect 17083 11172 17500 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 22664 11209 22692 11240
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11169 22707 11203
rect 22649 11163 22707 11169
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11940 11104 12357 11132
rect 11940 11092 11946 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 12986 11132 12992 11144
rect 12667 11104 12992 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13096 11104 13461 11132
rect 9508 11036 10640 11064
rect 8570 10996 8576 11008
rect 6932 10968 8576 10996
rect 6365 10959 6423 10965
rect 8570 10956 8576 10968
rect 8628 10996 8634 11008
rect 9508 10996 9536 11036
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 13096 11064 13124 11104
rect 13449 11101 13461 11104
rect 13495 11132 13507 11135
rect 13630 11132 13636 11144
rect 13495 11104 13636 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 17129 11135 17187 11141
rect 14332 11104 16989 11132
rect 14332 11092 14338 11104
rect 11112 11036 13124 11064
rect 13173 11067 13231 11073
rect 11112 11024 11118 11036
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13722 11064 13728 11076
rect 13219 11036 13728 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 15194 11024 15200 11076
rect 15252 11073 15258 11076
rect 15252 11067 15281 11073
rect 15269 11033 15281 11067
rect 15252 11027 15281 11033
rect 15413 11067 15471 11073
rect 15413 11033 15425 11067
rect 15459 11064 15471 11067
rect 15930 11064 15936 11076
rect 15459 11036 15936 11064
rect 15459 11033 15471 11036
rect 15413 11027 15471 11033
rect 15252 11024 15258 11027
rect 15930 11024 15936 11036
rect 15988 11024 15994 11076
rect 16022 11024 16028 11076
rect 16080 11024 16086 11076
rect 16850 11024 16856 11076
rect 16908 11024 16914 11076
rect 16961 11064 16989 11104
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17770 11132 17776 11144
rect 17175 11104 17776 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18892 11132 18920 11163
rect 18003 11104 18920 11132
rect 19429 11135 19487 11141
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19794 11132 19800 11144
rect 19475 11104 19800 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20128 11107 20530 11132
rect 20128 11104 20545 11107
rect 20128 11092 20134 11104
rect 20487 11101 20545 11104
rect 18417 11067 18475 11073
rect 18417 11064 18429 11067
rect 16961 11036 18429 11064
rect 18417 11033 18429 11036
rect 18463 11033 18475 11067
rect 18417 11027 18475 11033
rect 19610 11024 19616 11076
rect 19668 11024 19674 11076
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 20346 11064 20352 11076
rect 20303 11036 20352 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 20487 11067 20499 11101
rect 20533 11067 20545 11101
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21174 11132 21180 11144
rect 20772 11104 21180 11132
rect 20772 11092 20778 11104
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 23198 11132 23204 11144
rect 22235 11104 23204 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 26694 11092 26700 11144
rect 26752 11132 26758 11144
rect 26881 11135 26939 11141
rect 26881 11132 26893 11135
rect 26752 11104 26893 11132
rect 26752 11092 26758 11104
rect 26881 11101 26893 11104
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 27137 11135 27195 11141
rect 27137 11132 27149 11135
rect 27028 11104 27149 11132
rect 27028 11092 27034 11104
rect 27137 11101 27149 11104
rect 27183 11101 27195 11135
rect 27137 11095 27195 11101
rect 20487 11061 20545 11067
rect 20898 11024 20904 11076
rect 20956 11064 20962 11076
rect 21082 11064 21088 11076
rect 20956 11036 21088 11064
rect 20956 11024 20962 11036
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 21266 11024 21272 11076
rect 21324 11024 21330 11076
rect 21450 11024 21456 11076
rect 21508 11024 21514 11076
rect 22916 11067 22974 11073
rect 22916 11033 22928 11067
rect 22962 11064 22974 11067
rect 24670 11064 24676 11076
rect 22962 11036 24676 11064
rect 22962 11033 22974 11036
rect 22916 11027 22974 11033
rect 24670 11024 24676 11036
rect 24728 11024 24734 11076
rect 25130 11073 25136 11076
rect 25124 11064 25136 11073
rect 25091 11036 25136 11064
rect 25124 11027 25136 11036
rect 25130 11024 25136 11027
rect 25188 11024 25194 11076
rect 8628 10968 9536 10996
rect 8628 10956 8634 10968
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 9861 10999 9919 11005
rect 9861 10996 9873 10999
rect 9732 10968 9873 10996
rect 9732 10956 9738 10968
rect 9861 10965 9873 10968
rect 9907 10965 9919 10999
rect 9861 10959 9919 10965
rect 11238 10956 11244 11008
rect 11296 10956 11302 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12986 10996 12992 11008
rect 12492 10968 12992 10996
rect 12492 10956 12498 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 16114 10996 16120 11008
rect 15896 10968 16120 10996
rect 15896 10956 15902 10968
rect 16114 10956 16120 10968
rect 16172 10996 16178 11008
rect 16235 10999 16293 11005
rect 16235 10996 16247 10999
rect 16172 10968 16247 10996
rect 16172 10956 16178 10968
rect 16235 10965 16247 10968
rect 16281 10996 16293 10999
rect 17034 10996 17040 11008
rect 16281 10968 17040 10996
rect 16281 10965 16293 10968
rect 16235 10959 16293 10965
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 17770 10956 17776 11008
rect 17828 10956 17834 11008
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 19242 10996 19248 11008
rect 18380 10968 19248 10996
rect 18380 10956 18386 10968
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 19797 10999 19855 11005
rect 19797 10965 19809 10999
rect 19843 10996 19855 10999
rect 19886 10996 19892 11008
rect 19843 10968 19892 10996
rect 19843 10965 19855 10968
rect 19797 10959 19855 10965
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 21284 10996 21312 11024
rect 28261 10999 28319 11005
rect 28261 10996 28273 10999
rect 21284 10968 28273 10996
rect 28261 10965 28273 10968
rect 28307 10965 28319 10999
rect 28261 10959 28319 10965
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1946 10752 1952 10804
rect 2004 10801 2010 10804
rect 2004 10795 2023 10801
rect 2011 10761 2023 10795
rect 2004 10755 2023 10761
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 3418 10792 3424 10804
rect 2179 10764 3424 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 2004 10752 2010 10755
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 5258 10752 5264 10804
rect 5316 10801 5322 10804
rect 5316 10795 5335 10801
rect 5323 10761 5335 10795
rect 5316 10755 5335 10761
rect 5316 10752 5322 10755
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 12802 10792 12808 10804
rect 5592 10764 7512 10792
rect 5592 10752 5598 10764
rect 7484 10736 7512 10764
rect 9876 10764 12808 10792
rect 1765 10727 1823 10733
rect 1765 10693 1777 10727
rect 1811 10724 1823 10727
rect 2222 10724 2228 10736
rect 1811 10696 2228 10724
rect 1811 10693 1823 10696
rect 1765 10687 1823 10693
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 2590 10684 2596 10736
rect 2648 10684 2654 10736
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 3292 10696 5089 10724
rect 3292 10684 3298 10696
rect 5077 10693 5089 10696
rect 5123 10724 5135 10727
rect 5994 10724 6000 10736
rect 5123 10696 6000 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 7466 10684 7472 10736
rect 7524 10724 7530 10736
rect 7561 10727 7619 10733
rect 7561 10724 7573 10727
rect 7524 10696 7573 10724
rect 7524 10684 7530 10696
rect 7561 10693 7573 10696
rect 7607 10693 7619 10727
rect 7561 10687 7619 10693
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 8754 10724 8760 10736
rect 8435 10696 8760 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 6730 10656 6736 10668
rect 5684 10628 6736 10656
rect 5684 10616 5690 10628
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6972 10628 7021 10656
rect 6972 10616 6978 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8662 10656 8668 10668
rect 8619 10628 8668 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9674 10656 9680 10668
rect 9447 10628 9680 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 9876 10665 9904 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 12952 10764 14289 10792
rect 12952 10752 12958 10764
rect 14277 10761 14289 10764
rect 14323 10792 14335 10795
rect 15194 10792 15200 10804
rect 14323 10764 15200 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15344 10764 16313 10792
rect 15344 10752 15350 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 17034 10752 17040 10804
rect 17092 10801 17098 10804
rect 17092 10795 17111 10801
rect 17099 10761 17111 10795
rect 17092 10755 17111 10761
rect 17092 10752 17098 10755
rect 17218 10752 17224 10804
rect 17276 10752 17282 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18341 10795 18399 10801
rect 18341 10792 18353 10795
rect 18288 10764 18353 10792
rect 18288 10752 18294 10764
rect 18341 10761 18353 10764
rect 18387 10761 18399 10795
rect 18341 10755 18399 10761
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 20165 10795 20223 10801
rect 18555 10764 20116 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 12406 10727 12464 10733
rect 12406 10724 12418 10727
rect 10928 10696 12418 10724
rect 10928 10684 10934 10696
rect 12406 10693 12418 10696
rect 12452 10693 12464 10727
rect 12406 10687 12464 10693
rect 13538 10684 13544 10736
rect 13596 10724 13602 10736
rect 15933 10727 15991 10733
rect 15933 10724 15945 10727
rect 13596 10696 15945 10724
rect 13596 10684 13602 10696
rect 15933 10693 15945 10696
rect 15979 10693 15991 10727
rect 15933 10687 15991 10693
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 10962 10616 10968 10668
rect 11020 10616 11026 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12250 10656 12256 10668
rect 12207 10628 12256 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 13630 10656 13636 10668
rect 12308 10628 13636 10656
rect 12308 10616 12314 10628
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13964 10628 14197 10656
rect 13964 10616 13970 10628
rect 14185 10625 14197 10628
rect 14231 10656 14243 10659
rect 14366 10656 14372 10668
rect 14231 10628 14372 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 3418 10588 3424 10600
rect 2464 10560 3424 10588
rect 2464 10548 2470 10560
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 5442 10588 5448 10600
rect 5276 10560 5448 10588
rect 1670 10480 1676 10532
rect 1728 10520 1734 10532
rect 3881 10523 3939 10529
rect 3881 10520 3893 10523
rect 1728 10492 3893 10520
rect 1728 10480 1734 10492
rect 3881 10489 3893 10492
rect 3927 10489 3939 10523
rect 3881 10483 3939 10489
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 2130 10452 2136 10464
rect 1995 10424 2136 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 5276 10461 5304 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 11146 10588 11152 10600
rect 8803 10560 11152 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 10781 10523 10839 10529
rect 9263 10492 10732 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 4396 10424 5273 10452
rect 4396 10412 4402 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 6086 10452 6092 10464
rect 5491 10424 6092 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 7834 10452 7840 10464
rect 7607 10424 7840 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 10704 10452 10732 10492
rect 10781 10489 10793 10523
rect 10827 10520 10839 10523
rect 10870 10520 10876 10532
rect 10827 10492 10876 10520
rect 10827 10489 10839 10492
rect 10781 10483 10839 10489
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 14844 10520 14872 10619
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15948 10656 15976 10687
rect 16114 10684 16120 10736
rect 16172 10733 16178 10736
rect 16172 10727 16191 10733
rect 16179 10693 16191 10727
rect 16853 10727 16911 10733
rect 16853 10724 16865 10727
rect 16172 10687 16191 10693
rect 16592 10696 16865 10724
rect 16172 10684 16178 10687
rect 16482 10656 16488 10668
rect 15436 10628 15884 10656
rect 15948 10628 16488 10656
rect 15436 10616 15442 10628
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15746 10588 15752 10600
rect 15059 10560 15752 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 15856 10588 15884 10628
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16592 10588 16620 10696
rect 16853 10693 16865 10696
rect 16899 10724 16911 10727
rect 16942 10724 16948 10736
rect 16899 10696 16948 10724
rect 16899 10693 16911 10696
rect 16853 10687 16911 10693
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 18138 10684 18144 10736
rect 18196 10684 18202 10736
rect 18356 10656 18384 10755
rect 18782 10684 18788 10736
rect 18840 10724 18846 10736
rect 18969 10727 19027 10733
rect 18969 10724 18981 10727
rect 18840 10696 18981 10724
rect 18840 10684 18846 10696
rect 18969 10693 18981 10696
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 19199 10693 19257 10699
rect 19199 10690 19211 10693
rect 19189 10659 19211 10690
rect 19245 10659 19257 10693
rect 19426 10684 19432 10736
rect 19484 10724 19490 10736
rect 19797 10727 19855 10733
rect 19797 10724 19809 10727
rect 19484 10696 19809 10724
rect 19484 10684 19490 10696
rect 19797 10693 19809 10696
rect 19843 10693 19855 10727
rect 19797 10687 19855 10693
rect 19978 10684 19984 10736
rect 20036 10733 20042 10736
rect 20036 10727 20055 10733
rect 20043 10693 20055 10727
rect 20088 10724 20116 10764
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20438 10792 20444 10804
rect 20211 10764 20444 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20438 10752 20444 10764
rect 20496 10752 20502 10804
rect 22465 10795 22523 10801
rect 22465 10761 22477 10795
rect 22511 10761 22523 10795
rect 22465 10755 22523 10761
rect 22480 10724 22508 10755
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 23658 10792 23664 10804
rect 22612 10764 23664 10792
rect 22612 10752 22618 10764
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 25038 10752 25044 10804
rect 25096 10752 25102 10804
rect 20088 10696 22094 10724
rect 22480 10696 25728 10724
rect 20036 10687 20055 10693
rect 20036 10684 20042 10687
rect 19189 10656 19257 10659
rect 18356 10653 19257 10656
rect 18356 10628 19217 10653
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 20530 10656 20536 10668
rect 19392 10628 20536 10656
rect 19392 10616 19398 10628
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 19518 10588 19524 10600
rect 15856 10560 16620 10588
rect 17696 10560 19524 10588
rect 17696 10520 17724 10560
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 19794 10548 19800 10600
rect 19852 10588 19858 10600
rect 20254 10588 20260 10600
rect 19852 10560 20260 10588
rect 19852 10548 19858 10560
rect 20254 10548 20260 10560
rect 20312 10588 20318 10600
rect 20640 10588 20668 10619
rect 20806 10616 20812 10668
rect 20864 10616 20870 10668
rect 22066 10656 22094 10696
rect 22646 10656 22652 10668
rect 22066 10628 22652 10656
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 22922 10616 22928 10668
rect 22980 10656 22986 10668
rect 25700 10665 25728 10696
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22980 10628 23029 10656
rect 22980 10616 22986 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23917 10659 23975 10665
rect 23917 10656 23929 10659
rect 23017 10619 23075 10625
rect 23124 10628 23929 10656
rect 21082 10588 21088 10600
rect 20312 10560 21088 10588
rect 20312 10548 20318 10560
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 22005 10591 22063 10597
rect 22005 10557 22017 10591
rect 22051 10588 22063 10591
rect 22094 10588 22100 10600
rect 22051 10560 22100 10588
rect 22051 10557 22063 10560
rect 22005 10551 22063 10557
rect 22094 10548 22100 10560
rect 22152 10548 22158 10600
rect 23124 10588 23152 10628
rect 23917 10625 23929 10628
rect 23963 10625 23975 10659
rect 23917 10619 23975 10625
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 22204 10560 23152 10588
rect 23201 10591 23259 10597
rect 14844 10492 17724 10520
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 22204 10520 22232 10560
rect 23201 10557 23213 10591
rect 23247 10588 23259 10591
rect 23658 10588 23664 10600
rect 23247 10560 23664 10588
rect 23247 10557 23259 10560
rect 23201 10551 23259 10557
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 17828 10492 22232 10520
rect 22373 10523 22431 10529
rect 17828 10480 17834 10492
rect 22373 10489 22385 10523
rect 22419 10520 22431 10523
rect 22554 10520 22560 10532
rect 22419 10492 22560 10520
rect 22419 10489 22431 10492
rect 22373 10483 22431 10489
rect 22554 10480 22560 10492
rect 22612 10480 22618 10532
rect 25501 10523 25559 10529
rect 22756 10492 23244 10520
rect 11790 10452 11796 10464
rect 10704 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 12400 10424 13553 10452
rect 12400 10412 12406 10424
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 13541 10415 13599 10421
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 15194 10452 15200 10464
rect 15151 10424 15200 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15286 10412 15292 10464
rect 15344 10412 15350 10464
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16942 10452 16948 10464
rect 16163 10424 16948 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 17310 10452 17316 10464
rect 17083 10424 17316 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18966 10452 18972 10464
rect 18371 10424 18972 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 19242 10452 19248 10464
rect 19199 10424 19248 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19334 10412 19340 10464
rect 19392 10412 19398 10464
rect 19978 10412 19984 10464
rect 20036 10412 20042 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 22756 10452 22784 10492
rect 21039 10424 22784 10452
rect 23216 10452 23244 10492
rect 25501 10489 25513 10523
rect 25547 10520 25559 10523
rect 26786 10520 26792 10532
rect 25547 10492 26792 10520
rect 25547 10489 25559 10492
rect 25501 10483 25559 10489
rect 26786 10480 26792 10492
rect 26844 10480 26850 10532
rect 23842 10452 23848 10464
rect 23216 10424 23848 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 26142 10412 26148 10464
rect 26200 10412 26206 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 4028 10220 5641 10248
rect 4028 10208 4034 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 7374 10248 7380 10260
rect 6135 10220 7380 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 8444 10220 9505 10248
rect 8444 10208 8450 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10502 10248 10508 10260
rect 10275 10220 10508 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10502 10208 10508 10220
rect 10560 10248 10566 10260
rect 11054 10248 11060 10260
rect 10560 10220 11060 10248
rect 10560 10208 10566 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11974 10248 11980 10260
rect 11655 10220 11980 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 13170 10208 13176 10260
rect 13228 10208 13234 10260
rect 15286 10248 15292 10260
rect 13372 10220 15292 10248
rect 2130 10140 2136 10192
rect 2188 10180 2194 10192
rect 2774 10180 2780 10192
rect 2188 10152 2780 10180
rect 2188 10140 2194 10152
rect 2774 10140 2780 10152
rect 2832 10180 2838 10192
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 2832 10152 6561 10180
rect 2832 10140 2838 10152
rect 6549 10149 6561 10152
rect 6595 10149 6607 10183
rect 6549 10143 6607 10149
rect 9214 10140 9220 10192
rect 9272 10180 9278 10192
rect 9858 10180 9864 10192
rect 9272 10152 9864 10180
rect 9272 10140 9278 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10321 10183 10379 10189
rect 10321 10149 10333 10183
rect 10367 10180 10379 10183
rect 13372 10180 13400 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15654 10208 15660 10260
rect 15712 10208 15718 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 16632 10220 17325 10248
rect 16632 10208 16638 10220
rect 17313 10217 17325 10220
rect 17359 10248 17371 10251
rect 17678 10248 17684 10260
rect 17359 10220 17684 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 20438 10248 20444 10260
rect 19300 10220 20444 10248
rect 19300 10208 19306 10220
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 28353 10251 28411 10257
rect 28353 10248 28365 10251
rect 20864 10220 28365 10248
rect 20864 10208 20870 10220
rect 28353 10217 28365 10220
rect 28399 10217 28411 10251
rect 28353 10211 28411 10217
rect 10367 10152 13400 10180
rect 10367 10149 10379 10152
rect 10321 10143 10379 10149
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 18782 10180 18788 10192
rect 17276 10152 18788 10180
rect 17276 10140 17282 10152
rect 18782 10140 18788 10152
rect 18840 10180 18846 10192
rect 19613 10183 19671 10189
rect 19613 10180 19625 10183
rect 18840 10152 19625 10180
rect 18840 10140 18846 10152
rect 19613 10149 19625 10152
rect 19659 10180 19671 10183
rect 20346 10180 20352 10192
rect 19659 10152 20352 10180
rect 19659 10149 19671 10152
rect 19613 10143 19671 10149
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 20990 10140 20996 10192
rect 21048 10140 21054 10192
rect 21082 10140 21088 10192
rect 21140 10180 21146 10192
rect 21542 10180 21548 10192
rect 21140 10152 21548 10180
rect 21140 10140 21146 10152
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 21726 10140 21732 10192
rect 21784 10180 21790 10192
rect 21913 10183 21971 10189
rect 21913 10180 21925 10183
rect 21784 10152 21925 10180
rect 21784 10140 21790 10152
rect 21913 10149 21925 10152
rect 21959 10149 21971 10183
rect 21913 10143 21971 10149
rect 22097 10183 22155 10189
rect 22097 10149 22109 10183
rect 22143 10149 22155 10183
rect 22097 10143 22155 10149
rect 22925 10183 22983 10189
rect 22925 10149 22937 10183
rect 22971 10149 22983 10183
rect 22925 10143 22983 10149
rect 23017 10183 23075 10189
rect 23017 10149 23029 10183
rect 23063 10180 23075 10183
rect 23198 10180 23204 10192
rect 23063 10152 23204 10180
rect 23063 10149 23075 10152
rect 23017 10143 23075 10149
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3053 10115 3111 10121
rect 3053 10112 3065 10115
rect 3016 10084 3065 10112
rect 3016 10072 3022 10084
rect 3053 10081 3065 10084
rect 3099 10081 3111 10115
rect 5626 10112 5632 10124
rect 3053 10075 3111 10081
rect 4632 10084 5632 10112
rect 474 10004 480 10056
rect 532 10044 538 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 532 10016 1593 10044
rect 532 10004 538 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3510 10044 3516 10056
rect 3283 10016 3516 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4338 10044 4344 10056
rect 3620 10016 4344 10044
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 3620 9976 3648 10016
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4632 10053 4660 10084
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10112 5871 10115
rect 5994 10112 6000 10124
rect 5859 10084 6000 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8202 10112 8208 10124
rect 7975 10084 8208 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 12434 10112 12440 10124
rect 8444 10084 9352 10112
rect 8444 10072 8450 10084
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5534 10044 5540 10056
rect 4939 10016 5540 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 2464 9948 3648 9976
rect 2464 9936 2470 9948
rect 3694 9936 3700 9988
rect 3752 9976 3758 9988
rect 4724 9976 4752 10007
rect 3752 9948 4752 9976
rect 4816 9976 4844 10007
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6730 10044 6736 10056
rect 6595 10016 6736 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 6914 10044 6920 10056
rect 6871 10016 6920 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 8478 10044 8484 10056
rect 8128 10016 8484 10044
rect 4816 9948 5396 9976
rect 3752 9936 3758 9948
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 2038 9908 2044 9920
rect 1636 9880 2044 9908
rect 1636 9868 1642 9880
rect 2038 9868 2044 9880
rect 2096 9908 2102 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 2096 9880 3433 9908
rect 2096 9868 2102 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 5258 9908 5264 9920
rect 4479 9880 5264 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5368 9908 5396 9948
rect 5626 9936 5632 9988
rect 5684 9936 5690 9988
rect 7190 9976 7196 9988
rect 5736 9948 7196 9976
rect 5736 9908 5764 9948
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 8128 9976 8156 10016
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 9324 10053 9352 10084
rect 10704 10084 12440 10112
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10704 10053 10732 10084
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12710 10072 12716 10124
rect 12768 10072 12774 10124
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 12943 10084 13400 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9916 10016 10425 10044
rect 9916 10004 9922 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11664 10016 11805 10044
rect 11664 10004 11670 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11974 10044 11980 10056
rect 11793 10007 11851 10013
rect 11972 10004 11980 10044
rect 12032 10004 12038 10056
rect 12250 10004 12256 10056
rect 12308 10004 12314 10056
rect 12728 10044 12756 10072
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12728 10016 13001 10044
rect 12989 10013 13001 10016
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 7392 9948 8156 9976
rect 5368 9880 5764 9908
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 6822 9908 6828 9920
rect 6779 9880 6828 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 6822 9868 6828 9880
rect 6880 9908 6886 9920
rect 7392 9908 7420 9948
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 8938 9976 8944 9988
rect 8352 9948 8944 9976
rect 8352 9936 8358 9948
rect 8938 9936 8944 9948
rect 8996 9976 9002 9988
rect 9125 9979 9183 9985
rect 9125 9976 9137 9979
rect 8996 9948 9137 9976
rect 8996 9936 9002 9948
rect 9125 9945 9137 9948
rect 9171 9945 9183 9979
rect 9125 9939 9183 9945
rect 10318 9936 10324 9988
rect 10376 9976 10382 9988
rect 10376 9948 11100 9976
rect 10376 9936 10382 9948
rect 6880 9880 7420 9908
rect 6880 9868 6886 9880
rect 7466 9868 7472 9920
rect 7524 9868 7530 9920
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 10042 9908 10048 9920
rect 8435 9880 10048 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10597 9911 10655 9917
rect 10597 9877 10609 9911
rect 10643 9908 10655 9911
rect 10870 9908 10876 9920
rect 10643 9880 10876 9908
rect 10643 9877 10655 9880
rect 10597 9871 10655 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11072 9908 11100 9948
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11204 9948 11897 9976
rect 11204 9936 11210 9948
rect 11885 9945 11897 9948
rect 11931 9945 11943 9979
rect 11885 9939 11943 9945
rect 11972 9908 12000 10004
rect 12158 9985 12164 9988
rect 12115 9979 12164 9985
rect 12115 9945 12127 9979
rect 12161 9945 12164 9979
rect 12115 9939 12164 9945
rect 12158 9936 12164 9939
rect 12216 9936 12222 9988
rect 12710 9936 12716 9988
rect 12768 9936 12774 9988
rect 13372 9976 13400 10084
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 14277 10115 14335 10121
rect 14277 10112 14289 10115
rect 13688 10084 14289 10112
rect 13688 10072 13694 10084
rect 14277 10081 14289 10084
rect 14323 10081 14335 10115
rect 14277 10075 14335 10081
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 19242 10112 19248 10124
rect 17000 10084 19248 10112
rect 17000 10072 17006 10084
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 21358 10072 21364 10124
rect 21416 10112 21422 10124
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21416 10084 21649 10112
rect 21416 10072 21422 10084
rect 21637 10081 21649 10084
rect 21683 10112 21695 10115
rect 21818 10112 21824 10124
rect 21683 10084 21824 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 22112 10112 22140 10143
rect 22830 10112 22836 10124
rect 22112 10084 22836 10112
rect 22830 10072 22836 10084
rect 22888 10072 22894 10124
rect 22931 10112 22959 10143
rect 23198 10140 23204 10152
rect 23256 10140 23262 10192
rect 23845 10183 23903 10189
rect 23845 10149 23857 10183
rect 23891 10180 23903 10183
rect 24026 10180 24032 10192
rect 23891 10152 24032 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 23290 10112 23296 10124
rect 22931 10084 23296 10112
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 14533 10047 14591 10053
rect 14533 10044 14545 10047
rect 13504 10016 14545 10044
rect 13504 10004 13510 10016
rect 14533 10013 14545 10016
rect 14579 10013 14591 10047
rect 14533 10007 14591 10013
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16298 10004 16304 10056
rect 16356 10004 16362 10056
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17092 10016 18153 10044
rect 17092 10004 17098 10016
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 19426 10044 19432 10056
rect 18141 10007 18199 10013
rect 19306 10016 19432 10044
rect 16942 9976 16948 9988
rect 13372 9948 16948 9976
rect 16942 9936 16948 9948
rect 17000 9936 17006 9988
rect 17218 9936 17224 9988
rect 17276 9936 17282 9988
rect 11072 9880 12000 9908
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13630 9908 13636 9920
rect 12492 9880 13636 9908
rect 12492 9868 12498 9880
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 15930 9868 15936 9920
rect 15988 9908 15994 9920
rect 16485 9911 16543 9917
rect 16485 9908 16497 9911
rect 15988 9880 16497 9908
rect 15988 9868 15994 9880
rect 16485 9877 16497 9880
rect 16531 9877 16543 9911
rect 16485 9871 16543 9877
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 16908 9880 18245 9908
rect 16908 9868 16914 9880
rect 18233 9877 18245 9880
rect 18279 9908 18291 9911
rect 19306 9908 19334 10016
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 19978 10004 19984 10056
rect 20036 10044 20042 10056
rect 22094 10044 22100 10056
rect 20036 10016 22100 10044
rect 20036 10004 20042 10016
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 22186 10004 22192 10056
rect 22244 10044 22250 10056
rect 22462 10044 22468 10056
rect 22244 10016 22468 10044
rect 22244 10004 22250 10016
rect 22462 10004 22468 10016
rect 22520 10044 22526 10056
rect 22520 10016 22692 10044
rect 22520 10004 22526 10016
rect 20622 9936 20628 9988
rect 20680 9936 20686 9988
rect 21008 9948 21680 9976
rect 18279 9880 19334 9908
rect 18279 9877 18291 9880
rect 18233 9871 18291 9877
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 21008 9908 21036 9948
rect 19760 9880 21036 9908
rect 21085 9911 21143 9917
rect 19760 9868 19766 9880
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 21542 9908 21548 9920
rect 21131 9880 21548 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 21652 9908 21680 9948
rect 21818 9936 21824 9988
rect 21876 9976 21882 9988
rect 22557 9979 22615 9985
rect 22557 9976 22569 9979
rect 21876 9948 22569 9976
rect 21876 9936 21882 9948
rect 22557 9945 22569 9948
rect 22603 9945 22615 9979
rect 22664 9976 22692 10016
rect 25130 10004 25136 10056
rect 25188 10004 25194 10056
rect 26694 10004 26700 10056
rect 26752 10044 26758 10056
rect 26973 10047 27031 10053
rect 26973 10044 26985 10047
rect 26752 10016 26985 10044
rect 26752 10004 26758 10016
rect 26973 10013 26985 10016
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 23477 9979 23535 9985
rect 23477 9976 23489 9979
rect 22664 9948 23489 9976
rect 22557 9939 22615 9945
rect 23477 9945 23489 9948
rect 23523 9945 23535 9979
rect 23477 9939 23535 9945
rect 23860 9948 24164 9976
rect 23860 9908 23888 9948
rect 21652 9880 23888 9908
rect 23934 9868 23940 9920
rect 23992 9868 23998 9920
rect 24136 9908 24164 9948
rect 24854 9936 24860 9988
rect 24912 9976 24918 9988
rect 25378 9979 25436 9985
rect 25378 9976 25390 9979
rect 24912 9948 25390 9976
rect 24912 9936 24918 9948
rect 25378 9945 25390 9948
rect 25424 9945 25436 9979
rect 25378 9939 25436 9945
rect 26234 9936 26240 9988
rect 26292 9976 26298 9988
rect 27218 9979 27276 9985
rect 27218 9976 27230 9979
rect 26292 9948 27230 9976
rect 26292 9936 26298 9948
rect 27218 9945 27230 9948
rect 27264 9945 27276 9979
rect 27218 9939 27276 9945
rect 26513 9911 26571 9917
rect 26513 9908 26525 9911
rect 24136 9880 26525 9908
rect 26513 9877 26525 9880
rect 26559 9877 26571 9911
rect 26513 9871 26571 9877
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3970 9704 3976 9716
rect 3016 9676 3976 9704
rect 3016 9664 3022 9676
rect 3970 9664 3976 9676
rect 4028 9704 4034 9716
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 4028 9676 4077 9704
rect 4028 9664 4034 9676
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 6914 9704 6920 9716
rect 4065 9667 4123 9673
rect 4172 9676 6920 9704
rect 1394 9596 1400 9648
rect 1452 9636 1458 9648
rect 1826 9639 1884 9645
rect 1826 9636 1838 9639
rect 1452 9608 1838 9636
rect 1452 9596 1458 9608
rect 1826 9605 1838 9608
rect 1872 9605 1884 9639
rect 1826 9599 1884 9605
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 3234 9636 3240 9648
rect 2832 9608 3240 9636
rect 2832 9596 2838 9608
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 3694 9596 3700 9648
rect 3752 9636 3758 9648
rect 4172 9636 4200 9676
rect 6914 9664 6920 9676
rect 6972 9664 6978 9716
rect 8297 9707 8355 9713
rect 8297 9673 8309 9707
rect 8343 9704 8355 9707
rect 8570 9704 8576 9716
rect 8343 9676 8576 9704
rect 8343 9673 8355 9676
rect 8297 9667 8355 9673
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 9217 9707 9275 9713
rect 9217 9673 9229 9707
rect 9263 9674 9275 9707
rect 9263 9673 9352 9674
rect 9217 9667 9352 9673
rect 3752 9608 4200 9636
rect 4709 9639 4767 9645
rect 3752 9596 3758 9608
rect 4709 9605 4721 9639
rect 4755 9636 4767 9639
rect 4982 9636 4988 9648
rect 4755 9608 4988 9636
rect 4755 9605 4767 9608
rect 4709 9599 4767 9605
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6604 9608 6653 9636
rect 6604 9596 6610 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7282 9636 7288 9648
rect 7055 9608 7288 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 9232 9646 9352 9667
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 9640 9676 12020 9704
rect 9640 9664 9646 9676
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 1670 9568 1676 9580
rect 1627 9540 1676 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 3881 9571 3939 9577
rect 2280 9540 2636 9568
rect 2280 9528 2286 9540
rect 2608 9432 2636 9540
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4062 9568 4068 9580
rect 3927 9540 4068 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 4172 9500 4200 9531
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4396 9540 4629 9568
rect 4396 9528 4402 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 3568 9472 4200 9500
rect 4816 9500 4844 9531
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5718 9568 5724 9580
rect 5491 9540 5724 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 7926 9528 7932 9580
rect 7984 9528 7990 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 9324 9568 9352 9646
rect 9398 9596 9404 9648
rect 9456 9636 9462 9648
rect 9950 9636 9956 9648
rect 9456 9608 9956 9636
rect 9456 9596 9462 9608
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 10192 9608 10333 9636
rect 10192 9596 10198 9608
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10321 9599 10379 9605
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 11606 9636 11612 9648
rect 10468 9608 11612 9636
rect 10468 9596 10474 9608
rect 11606 9596 11612 9608
rect 11664 9636 11670 9648
rect 11992 9636 12020 9676
rect 13096 9676 14044 9704
rect 12069 9639 12127 9645
rect 12069 9636 12081 9639
rect 11664 9608 11928 9636
rect 11992 9608 12081 9636
rect 11664 9596 11670 9608
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 8159 9540 9168 9568
rect 9324 9540 9873 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 4982 9500 4988 9512
rect 4816 9472 4988 9500
rect 3568 9460 3574 9472
rect 2608 9404 3556 9432
rect 3528 9376 3556 9404
rect 4080 9376 4108 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9140 9500 9168 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 10962 9568 10968 9580
rect 9861 9531 9919 9537
rect 10244 9540 10968 9568
rect 10244 9500 10272 9540
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11900 9577 11928 9608
rect 12069 9605 12081 9608
rect 12115 9605 12127 9639
rect 12069 9599 12127 9605
rect 12158 9596 12164 9648
rect 12216 9645 12222 9648
rect 12216 9639 12245 9645
rect 12233 9636 12245 9639
rect 12233 9608 12434 9636
rect 12233 9605 12245 9608
rect 12216 9599 12245 9605
rect 12216 9596 12222 9599
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12299 9571 12357 9577
rect 12299 9568 12311 9571
rect 12084 9540 12311 9568
rect 9140 9472 10272 9500
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 11716 9500 11744 9528
rect 12084 9500 12112 9540
rect 12299 9537 12311 9540
rect 12345 9537 12357 9571
rect 12299 9531 12357 9537
rect 11716 9472 12112 9500
rect 12406 9500 12434 9608
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 12860 9608 12909 9636
rect 12860 9596 12866 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 13096 9500 13124 9676
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 14016 9636 14044 9676
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 15470 9704 15476 9716
rect 14884 9676 15476 9704
rect 14884 9664 14890 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 20990 9664 20996 9716
rect 21048 9704 21054 9716
rect 24026 9704 24032 9716
rect 21048 9676 24032 9704
rect 21048 9664 21054 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 24486 9664 24492 9716
rect 24544 9704 24550 9716
rect 25130 9704 25136 9716
rect 24544 9676 25136 9704
rect 24544 9664 24550 9676
rect 25130 9664 25136 9676
rect 25188 9704 25194 9716
rect 26694 9704 26700 9716
rect 25188 9676 26700 9704
rect 25188 9664 25194 9676
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 14182 9636 14188 9648
rect 13228 9608 13952 9636
rect 14016 9608 14188 9636
rect 13228 9596 13234 9608
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13924 9577 13952 9608
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 14332 9608 14381 9636
rect 14332 9596 14338 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 14569 9639 14627 9645
rect 14569 9636 14581 9639
rect 14369 9599 14427 9605
rect 14476 9608 14581 9636
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13412 9540 13737 9568
rect 13412 9528 13418 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14476 9568 14504 9608
rect 14569 9605 14581 9608
rect 14615 9605 14627 9639
rect 14569 9599 14627 9605
rect 15102 9596 15108 9648
rect 15160 9596 15166 9648
rect 15321 9639 15379 9645
rect 15321 9605 15333 9639
rect 15367 9636 15379 9639
rect 15367 9608 17356 9636
rect 15367 9605 15379 9608
rect 15321 9599 15379 9605
rect 14056 9540 14504 9568
rect 14056 9528 14062 9540
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 15804 9540 16313 9568
rect 15804 9528 15810 9540
rect 16301 9537 16313 9540
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16540 9540 16957 9568
rect 16540 9528 16546 9540
rect 16945 9537 16957 9540
rect 16991 9568 17003 9571
rect 17218 9568 17224 9580
rect 16991 9540 17224 9568
rect 16991 9537 17003 9540
rect 16945 9531 17003 9537
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 17328 9568 17356 9608
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 17460 9608 17693 9636
rect 17460 9596 17466 9608
rect 17681 9605 17693 9608
rect 17727 9605 17739 9639
rect 17681 9599 17739 9605
rect 18248 9608 18828 9636
rect 17954 9568 17960 9580
rect 17328 9540 17960 9568
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18248 9577 18276 9608
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 14458 9500 14464 9512
rect 12406 9472 13124 9500
rect 13372 9472 14464 9500
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 10226 9432 10232 9444
rect 9171 9404 10232 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9401 10747 9435
rect 10689 9395 10747 9401
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 13372 9432 13400 9472
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14608 9472 14780 9500
rect 14608 9460 14614 9472
rect 11747 9404 13400 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 992 9336 2973 9364
rect 992 9324 998 9336
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 2961 9327 3019 9333
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3568 9336 3709 9364
rect 3568 9324 3574 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3697 9327 3755 9333
rect 4062 9324 4068 9376
rect 4120 9324 4126 9376
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4338 9364 4344 9376
rect 4212 9336 4344 9364
rect 4212 9324 4218 9336
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 5074 9364 5080 9376
rect 4948 9336 5080 9364
rect 4948 9324 4954 9336
rect 5074 9324 5080 9336
rect 5132 9364 5138 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5132 9336 5641 9364
rect 5132 9324 5138 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 5629 9327 5687 9333
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9582 9364 9588 9376
rect 8904 9336 9588 9364
rect 8904 9324 8910 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 10704 9364 10732 9395
rect 13446 9392 13452 9444
rect 13504 9432 13510 9444
rect 14752 9441 14780 9472
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15286 9500 15292 9512
rect 15160 9472 15292 9500
rect 15160 9460 15166 9472
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 18432 9500 18460 9531
rect 15988 9472 18460 9500
rect 18800 9500 18828 9608
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 18932 9608 19257 9636
rect 18932 9596 18938 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19245 9599 19303 9605
rect 19794 9596 19800 9648
rect 19852 9636 19858 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19852 9608 20269 9636
rect 19852 9596 19858 9608
rect 20257 9605 20269 9608
rect 20303 9636 20315 9639
rect 20622 9636 20628 9648
rect 20303 9608 20628 9636
rect 20303 9605 20315 9608
rect 20257 9599 20315 9605
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 21450 9596 21456 9648
rect 21508 9636 21514 9648
rect 22646 9636 22652 9648
rect 21508 9608 22652 9636
rect 21508 9596 21514 9608
rect 22646 9596 22652 9608
rect 22704 9596 22710 9648
rect 22738 9596 22744 9648
rect 22796 9636 22802 9648
rect 26234 9636 26240 9648
rect 22796 9608 26240 9636
rect 22796 9596 22802 9608
rect 26234 9596 26240 9608
rect 26292 9596 26298 9648
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9568 19119 9571
rect 19334 9568 19340 9580
rect 19107 9540 19340 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21269 9571 21327 9577
rect 21269 9568 21281 9571
rect 21140 9540 21281 9568
rect 21140 9528 21146 9540
rect 21269 9537 21281 9540
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9568 22247 9571
rect 22278 9568 22284 9580
rect 22235 9540 22284 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 22830 9528 22836 9580
rect 22888 9528 22894 9580
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 24486 9568 24492 9580
rect 23716 9540 24492 9568
rect 23716 9528 23722 9540
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 24756 9571 24814 9577
rect 24756 9537 24768 9571
rect 24802 9568 24814 9571
rect 24802 9540 26372 9568
rect 24802 9537 24814 9540
rect 24756 9531 24814 9537
rect 20070 9500 20076 9512
rect 18800 9472 20076 9500
rect 15988 9460 15994 9472
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 14737 9435 14795 9441
rect 13504 9404 14688 9432
rect 13504 9392 13510 9404
rect 12066 9364 12072 9376
rect 10704 9336 12072 9364
rect 12066 9324 12072 9336
rect 12124 9364 12130 9376
rect 12618 9364 12624 9376
rect 12124 9336 12624 9364
rect 12124 9324 12130 9336
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12952 9336 13001 9364
rect 12952 9324 12958 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13136 9336 13829 9364
rect 13136 9324 13142 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 13964 9336 14565 9364
rect 13964 9324 13970 9336
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 14660 9364 14688 9404
rect 14737 9401 14749 9435
rect 14783 9401 14795 9435
rect 15473 9435 15531 9441
rect 15473 9432 15485 9435
rect 14737 9395 14795 9401
rect 14844 9404 15485 9432
rect 14844 9364 14872 9404
rect 15473 9401 15485 9404
rect 15519 9401 15531 9435
rect 15473 9395 15531 9401
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 18141 9435 18199 9441
rect 18141 9432 18153 9435
rect 15896 9404 18153 9432
rect 15896 9392 15902 9404
rect 18141 9401 18153 9404
rect 18187 9401 18199 9435
rect 18141 9395 18199 9401
rect 19702 9392 19708 9444
rect 19760 9432 19766 9444
rect 20533 9435 20591 9441
rect 20533 9432 20545 9435
rect 19760 9404 20545 9432
rect 19760 9392 19766 9404
rect 20533 9401 20545 9404
rect 20579 9401 20591 9435
rect 20533 9395 20591 9401
rect 22002 9392 22008 9444
rect 22060 9392 22066 9444
rect 23385 9435 23443 9441
rect 23385 9401 23397 9435
rect 23431 9432 23443 9435
rect 24394 9432 24400 9444
rect 23431 9404 24400 9432
rect 23431 9401 23443 9404
rect 23385 9395 23443 9401
rect 24394 9392 24400 9404
rect 24452 9392 24458 9444
rect 26344 9441 26372 9540
rect 26510 9528 26516 9580
rect 26568 9528 26574 9580
rect 26329 9435 26387 9441
rect 26329 9401 26341 9435
rect 26375 9401 26387 9435
rect 26329 9395 26387 9401
rect 14660 9336 14872 9364
rect 14553 9327 14611 9333
rect 15286 9324 15292 9376
rect 15344 9324 15350 9376
rect 15746 9324 15752 9376
rect 15804 9324 15810 9376
rect 16114 9324 16120 9376
rect 16172 9324 16178 9376
rect 17034 9324 17040 9376
rect 17092 9324 17098 9376
rect 17954 9324 17960 9376
rect 18012 9324 18018 9376
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 20622 9364 20628 9376
rect 19475 9336 20628 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9364 20775 9367
rect 21266 9364 21272 9376
rect 20763 9336 21272 9364
rect 20763 9333 20775 9336
rect 20717 9327 20775 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21358 9324 21364 9376
rect 21416 9324 21422 9376
rect 22649 9367 22707 9373
rect 22649 9333 22661 9367
rect 22695 9364 22707 9367
rect 22738 9364 22744 9376
rect 22695 9336 22744 9364
rect 22695 9333 22707 9336
rect 22649 9327 22707 9333
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 25869 9367 25927 9373
rect 25869 9364 25881 9367
rect 23808 9336 25881 9364
rect 23808 9324 23814 9336
rect 25869 9333 25881 9336
rect 25915 9333 25927 9367
rect 25869 9327 25927 9333
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1762 9160 1768 9172
rect 1719 9132 1768 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2498 9120 2504 9172
rect 2556 9120 2562 9172
rect 3234 9120 3240 9172
rect 3292 9120 3298 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4706 9160 4712 9172
rect 3476 9132 4712 9160
rect 3476 9120 3482 9132
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 4856 9132 4905 9160
rect 4856 9120 4862 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 4893 9123 4951 9129
rect 6733 9163 6791 9169
rect 6733 9129 6745 9163
rect 6779 9160 6791 9163
rect 6822 9160 6828 9172
rect 6779 9132 6828 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7340 9132 7696 9160
rect 7340 9120 7346 9132
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 4341 9095 4399 9101
rect 4341 9092 4353 9095
rect 2740 9064 4353 9092
rect 2740 9052 2746 9064
rect 4341 9061 4353 9064
rect 4387 9092 4399 9095
rect 5074 9092 5080 9104
rect 4387 9064 5080 9092
rect 4387 9061 4399 9064
rect 4341 9055 4399 9061
rect 5074 9052 5080 9064
rect 5132 9052 5138 9104
rect 5718 9052 5724 9104
rect 5776 9092 5782 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 5776 9064 7481 9092
rect 5776 9052 5782 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 7469 9055 7527 9061
rect 2424 8996 2774 9024
rect 1026 8916 1032 8968
rect 1084 8956 1090 8968
rect 2424 8965 2452 8996
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1084 8928 1685 8956
rect 1084 8916 1090 8928
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 1872 8888 1900 8919
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 2746 8956 2774 8996
rect 3970 8984 3976 9036
rect 4028 8984 4034 9036
rect 4890 9024 4896 9036
rect 4080 8996 4896 9024
rect 4080 8956 4108 8996
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 7006 9024 7012 9036
rect 5460 8996 7012 9024
rect 2746 8928 4108 8956
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4522 8956 4528 8968
rect 4203 8928 4528 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 5460 8965 5488 8996
rect 7006 8984 7012 8996
rect 7064 9024 7070 9036
rect 7668 9024 7696 9132
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 7800 9132 8401 9160
rect 7800 9120 7806 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 9766 9120 9772 9172
rect 9824 9120 9830 9172
rect 10134 9160 10140 9172
rect 9876 9132 10140 9160
rect 8294 9052 8300 9104
rect 8352 9052 8358 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9876 9092 9904 9132
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11517 9163 11575 9169
rect 11517 9129 11529 9163
rect 11563 9160 11575 9163
rect 11606 9160 11612 9172
rect 11563 9132 11612 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 11882 9160 11888 9172
rect 11747 9132 11888 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 12526 9120 12532 9172
rect 12584 9120 12590 9172
rect 12986 9120 12992 9172
rect 13044 9120 13050 9172
rect 13446 9120 13452 9172
rect 13504 9120 13510 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 14458 9160 14464 9172
rect 13872 9132 14464 9160
rect 13872 9120 13878 9132
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 14642 9160 14648 9172
rect 14599 9132 14648 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 14918 9160 14924 9172
rect 14792 9132 14924 9160
rect 14792 9120 14798 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15580 9132 15669 9160
rect 8904 9064 9904 9092
rect 9953 9095 10011 9101
rect 8904 9052 8910 9064
rect 9953 9061 9965 9095
rect 9999 9061 10011 9095
rect 9953 9055 10011 9061
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 7064 8996 7420 9024
rect 7668 8996 8493 9024
rect 7064 8984 7070 8996
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 2682 8888 2688 8900
rect 1872 8860 2688 8888
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 3053 8891 3111 8897
rect 3053 8888 3065 8891
rect 2924 8860 3065 8888
rect 2924 8848 2930 8860
rect 3053 8857 3065 8860
rect 3099 8857 3111 8891
rect 3053 8851 3111 8857
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 4816 8888 4844 8919
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5592 8928 5641 8956
rect 5592 8916 5598 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7392 8965 7420 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 9968 9024 9996 9055
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 10686 9092 10692 9104
rect 10560 9064 10692 9092
rect 10560 9052 10566 9064
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 13265 9095 13323 9101
rect 11696 9064 12572 9092
rect 11696 9024 11724 9064
rect 9968 8996 11724 9024
rect 12544 9024 12572 9064
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 15580 9092 15608 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 17218 9120 17224 9172
rect 17276 9120 17282 9172
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9129 18199 9163
rect 18141 9123 18199 9129
rect 13311 9064 15608 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 12544 8996 13369 9024
rect 8481 8987 8539 8993
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 13872 8996 14381 9024
rect 13872 8984 13878 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15596 9024 15792 9032
rect 15068 9004 16252 9024
rect 15068 8996 15624 9004
rect 15764 8996 16252 9004
rect 15068 8984 15074 8996
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7708 8928 7757 8956
rect 7708 8916 7714 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 3660 8860 4844 8888
rect 3660 8848 3666 8860
rect 6454 8848 6460 8900
rect 6512 8848 6518 8900
rect 7668 8888 7696 8916
rect 6932 8860 7696 8888
rect 8220 8888 8248 8919
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 9088 8928 10425 8956
rect 9088 8916 9094 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10652 8928 12209 8956
rect 10652 8916 10658 8928
rect 11348 8900 11376 8928
rect 9398 8888 9404 8900
rect 8220 8860 9404 8888
rect 6932 8832 6960 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 9582 8848 9588 8900
rect 9640 8848 9646 8900
rect 10778 8888 10784 8900
rect 9692 8860 10784 8888
rect 3234 8780 3240 8832
rect 3292 8829 3298 8832
rect 3292 8823 3311 8829
rect 3299 8789 3311 8823
rect 3292 8783 3311 8789
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 4154 8820 4160 8832
rect 3467 8792 4160 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 3292 8780 3298 8783
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 4672 8792 5825 8820
rect 4672 8780 4678 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 6914 8780 6920 8832
rect 6972 8780 6978 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7064 8792 7481 8820
rect 7064 8780 7070 8792
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 7558 8780 7564 8832
rect 7616 8780 7622 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 9692 8820 9720 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 11330 8848 11336 8900
rect 11388 8848 11394 8900
rect 12181 8897 12209 8928
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 12676 8928 13553 8956
rect 12676 8916 12682 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13688 8928 13737 8956
rect 13688 8916 13694 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 14550 8916 14556 8968
rect 14608 8916 14614 8968
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15528 8928 16129 8956
rect 15528 8916 15534 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16224 8956 16252 8996
rect 16373 8959 16431 8965
rect 16373 8956 16385 8959
rect 16224 8928 16385 8956
rect 16117 8919 16175 8925
rect 16373 8925 16385 8928
rect 16419 8925 16431 8959
rect 17236 8956 17264 9120
rect 18156 9092 18184 9123
rect 19610 9120 19616 9172
rect 19668 9120 19674 9172
rect 20625 9163 20683 9169
rect 20625 9129 20637 9163
rect 20671 9160 20683 9163
rect 22830 9160 22836 9172
rect 20671 9132 22836 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 24026 9120 24032 9172
rect 24084 9120 24090 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 24820 9132 25973 9160
rect 24820 9120 24826 9132
rect 25961 9129 25973 9132
rect 26007 9129 26019 9163
rect 25961 9123 26019 9129
rect 27982 9120 27988 9172
rect 28040 9160 28046 9172
rect 28077 9163 28135 9169
rect 28077 9160 28089 9163
rect 28040 9132 28089 9160
rect 28040 9120 28046 9132
rect 28077 9129 28089 9132
rect 28123 9129 28135 9163
rect 28077 9123 28135 9129
rect 19797 9095 19855 9101
rect 18156 9064 19748 9092
rect 19426 8984 19432 9036
rect 19484 8984 19490 9036
rect 18874 8956 18880 8968
rect 17236 8928 18880 8956
rect 16373 8919 16431 8925
rect 11549 8891 11607 8897
rect 11549 8857 11561 8891
rect 11595 8888 11607 8891
rect 12161 8891 12219 8897
rect 11595 8860 11944 8888
rect 11595 8857 11607 8860
rect 11549 8851 11607 8857
rect 8352 8792 9720 8820
rect 9795 8823 9853 8829
rect 8352 8780 8358 8792
rect 9795 8789 9807 8823
rect 9841 8820 9853 8823
rect 10410 8820 10416 8832
rect 9841 8792 10416 8820
rect 9841 8789 9853 8792
rect 9795 8783 9853 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10652 8792 10885 8820
rect 10652 8780 10658 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 11916 8820 11944 8860
rect 12161 8857 12173 8891
rect 12207 8857 12219 8891
rect 12161 8851 12219 8857
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 12361 8891 12419 8897
rect 12361 8888 12373 8891
rect 12308 8860 12373 8888
rect 12308 8848 12314 8860
rect 12361 8857 12373 8860
rect 12407 8857 12419 8891
rect 12361 8851 12419 8857
rect 14274 8848 14280 8900
rect 14332 8848 14338 8900
rect 17972 8897 18000 8928
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8857 15347 8891
rect 15289 8851 15347 8857
rect 17957 8891 18015 8897
rect 17957 8857 17969 8891
rect 18003 8857 18015 8891
rect 17957 8851 18015 8857
rect 18173 8891 18231 8897
rect 18173 8857 18185 8891
rect 18219 8888 18231 8891
rect 19150 8888 19156 8900
rect 18219 8860 19156 8888
rect 18219 8857 18231 8860
rect 18173 8851 18231 8857
rect 13170 8820 13176 8832
rect 11916 8792 13176 8820
rect 10873 8783 10931 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 13780 8792 14749 8820
rect 13780 8780 13786 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 15304 8820 15332 8851
rect 19150 8848 19156 8860
rect 19208 8848 19214 8900
rect 19444 8897 19472 8984
rect 19720 8956 19748 9064
rect 19797 9061 19809 9095
rect 19843 9061 19855 9095
rect 19797 9055 19855 9061
rect 21085 9095 21143 9101
rect 21085 9061 21097 9095
rect 21131 9092 21143 9095
rect 21131 9064 22600 9092
rect 21131 9061 21143 9064
rect 21085 9055 21143 9061
rect 19812 9024 19840 9055
rect 22370 9024 22376 9036
rect 19812 8996 22376 9024
rect 22370 8984 22376 8996
rect 22428 8984 22434 9036
rect 19720 8928 20576 8956
rect 19429 8891 19487 8897
rect 19429 8857 19441 8891
rect 19475 8857 19487 8891
rect 19429 8851 19487 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 20254 8888 20260 8900
rect 19576 8860 20260 8888
rect 19576 8848 19582 8860
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 20438 8848 20444 8900
rect 20496 8848 20502 8900
rect 20548 8888 20576 8928
rect 21266 8916 21272 8968
rect 21324 8916 21330 8968
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21600 8928 21925 8956
rect 21600 8916 21606 8928
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 22370 8888 22376 8900
rect 20548 8860 22376 8888
rect 22370 8848 22376 8860
rect 22428 8848 22434 8900
rect 15160 8792 15332 8820
rect 15499 8823 15557 8829
rect 15160 8780 15166 8792
rect 15499 8789 15511 8823
rect 15545 8820 15557 8823
rect 16022 8820 16028 8832
rect 15545 8792 16028 8820
rect 15545 8789 15557 8792
rect 15499 8783 15557 8789
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 17497 8823 17555 8829
rect 17497 8820 17509 8823
rect 16356 8792 17509 8820
rect 16356 8780 16362 8792
rect 17497 8789 17509 8792
rect 17543 8789 17555 8823
rect 17497 8783 17555 8789
rect 18322 8780 18328 8832
rect 18380 8780 18386 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 19629 8823 19687 8829
rect 19629 8820 19641 8823
rect 19116 8792 19641 8820
rect 19116 8780 19122 8792
rect 19629 8789 19641 8792
rect 19675 8789 19687 8823
rect 20456 8820 20484 8848
rect 20898 8820 20904 8832
rect 20456 8792 20904 8820
rect 19629 8783 19687 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 21729 8823 21787 8829
rect 21729 8789 21741 8823
rect 21775 8820 21787 8823
rect 22462 8820 22468 8832
rect 21775 8792 22468 8820
rect 21775 8789 21787 8792
rect 21729 8783 21787 8789
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 22572 8820 22600 9064
rect 26694 8984 26700 9036
rect 26752 8984 26758 9036
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8956 22707 8959
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 22695 8928 24593 8956
rect 22695 8925 22707 8928
rect 22649 8919 22707 8925
rect 23124 8900 23152 8928
rect 24581 8925 24593 8928
rect 24627 8956 24639 8959
rect 24670 8956 24676 8968
rect 24627 8928 24676 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 26786 8916 26792 8968
rect 26844 8956 26850 8968
rect 26953 8959 27011 8965
rect 26953 8956 26965 8959
rect 26844 8928 26965 8956
rect 26844 8916 26850 8928
rect 26953 8925 26965 8928
rect 26999 8925 27011 8959
rect 26953 8919 27011 8925
rect 22738 8848 22744 8900
rect 22796 8888 22802 8900
rect 22894 8891 22952 8897
rect 22894 8888 22906 8891
rect 22796 8860 22906 8888
rect 22796 8848 22802 8860
rect 22894 8857 22906 8860
rect 22940 8857 22952 8891
rect 22894 8851 22952 8857
rect 23106 8848 23112 8900
rect 23164 8848 23170 8900
rect 23566 8848 23572 8900
rect 23624 8888 23630 8900
rect 24826 8891 24884 8897
rect 24826 8888 24838 8891
rect 23624 8860 24838 8888
rect 23624 8848 23630 8860
rect 24826 8857 24838 8860
rect 24872 8857 24884 8891
rect 24826 8851 24884 8857
rect 24946 8820 24952 8832
rect 22572 8792 24952 8820
rect 24946 8780 24952 8792
rect 25004 8780 25010 8832
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 658 8576 664 8628
rect 716 8616 722 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 716 8588 3617 8616
rect 716 8576 722 8588
rect 3605 8585 3617 8588
rect 3651 8585 3663 8619
rect 3605 8579 3663 8585
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 4522 8576 4528 8628
rect 4580 8576 4586 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 5960 8588 9137 8616
rect 5960 8576 5966 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 11054 8616 11060 8628
rect 9125 8579 9183 8585
rect 9324 8588 11060 8616
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 1826 8551 1884 8557
rect 1826 8548 1838 8551
rect 1360 8520 1838 8548
rect 1360 8508 1366 8520
rect 1826 8517 1838 8520
rect 1872 8517 1884 8551
rect 1826 8511 1884 8517
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 3786 8548 3792 8560
rect 2372 8520 2774 8548
rect 2372 8508 2378 8520
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1670 8480 1676 8492
rect 1627 8452 1676 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 2746 8412 2774 8520
rect 3528 8520 3792 8548
rect 3528 8489 3556 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 4356 8548 4384 8576
rect 5442 8548 5448 8560
rect 4356 8520 5448 8548
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5534 8508 5540 8560
rect 5592 8508 5598 8560
rect 5626 8508 5632 8560
rect 5684 8548 5690 8560
rect 5994 8548 6000 8560
rect 5684 8520 6000 8548
rect 5684 8508 5690 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6104 8520 7205 8548
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4264 8452 4537 8480
rect 4264 8412 4292 8452
rect 4525 8449 4537 8452
rect 4571 8480 4583 8483
rect 4614 8480 4620 8492
rect 4571 8452 4620 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4890 8480 4896 8492
rect 4764 8452 4896 8480
rect 4764 8440 4770 8452
rect 4890 8440 4896 8452
rect 4948 8480 4954 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 4948 8452 5365 8480
rect 4948 8440 4954 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 6104 8480 6132 8520
rect 7193 8517 7205 8520
rect 7239 8517 7251 8551
rect 7193 8511 7251 8517
rect 7653 8551 7711 8557
rect 7653 8517 7665 8551
rect 7699 8548 7711 8551
rect 8478 8548 8484 8560
rect 7699 8520 8484 8548
rect 7699 8517 7711 8520
rect 7653 8511 7711 8517
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 9030 8548 9036 8560
rect 8711 8520 9036 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 5353 8443 5411 8449
rect 5644 8452 6132 8480
rect 5644 8424 5672 8452
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 9324 8480 9352 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8585 11207 8619
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 11149 8579 11207 8585
rect 12406 8588 13093 8616
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 11164 8548 11192 8579
rect 9456 8520 11192 8548
rect 9456 8508 9462 8520
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11946 8551 12004 8557
rect 11946 8548 11958 8551
rect 11848 8520 11958 8548
rect 11848 8508 11854 8520
rect 11946 8517 11958 8520
rect 11992 8517 12004 8551
rect 11946 8511 12004 8517
rect 7668 8452 9352 8480
rect 2746 8384 4292 8412
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 4396 8384 4445 8412
rect 4396 8372 4402 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 7668 8412 7696 8452
rect 8113 8415 8171 8421
rect 8113 8412 8125 8415
rect 5767 8384 7696 8412
rect 7760 8384 8125 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 6178 8344 6184 8356
rect 3007 8316 6184 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7760 8344 7788 8384
rect 8113 8381 8125 8384
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 7616 8316 7788 8344
rect 8021 8347 8079 8353
rect 7616 8304 7622 8316
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8294 8344 8300 8356
rect 8067 8316 8300 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 8846 8344 8852 8356
rect 8536 8316 8852 8344
rect 8536 8304 8542 8316
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 9416 8344 9444 8508
rect 10036 8483 10094 8489
rect 10036 8449 10048 8483
rect 10082 8480 10094 8483
rect 10410 8480 10416 8492
rect 10082 8452 10416 8480
rect 10082 8449 10094 8452
rect 10036 8443 10094 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 12406 8480 12434 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14792 8588 14933 8616
rect 14792 8576 14798 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 15562 8576 15568 8628
rect 15620 8625 15626 8628
rect 15620 8619 15639 8625
rect 15627 8616 15639 8619
rect 15749 8619 15807 8625
rect 15627 8588 15700 8616
rect 15627 8585 15639 8588
rect 15620 8579 15639 8585
rect 15620 8576 15626 8579
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 14553 8551 14611 8557
rect 14553 8548 14565 8551
rect 14240 8520 14565 8548
rect 14240 8508 14246 8520
rect 14553 8517 14565 8520
rect 14599 8517 14611 8551
rect 14553 8511 14611 8517
rect 15378 8508 15384 8560
rect 15436 8508 15442 8560
rect 15672 8548 15700 8588
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 15838 8616 15844 8628
rect 15795 8588 15844 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16298 8616 16304 8628
rect 15948 8588 16304 8616
rect 15948 8548 15976 8588
rect 16298 8576 16304 8588
rect 16356 8616 16362 8628
rect 17053 8619 17111 8625
rect 17053 8616 17065 8619
rect 16356 8588 17065 8616
rect 16356 8576 16362 8588
rect 17053 8585 17065 8588
rect 17099 8585 17111 8619
rect 17053 8579 17111 8585
rect 17218 8576 17224 8628
rect 17276 8576 17282 8628
rect 17891 8619 17949 8625
rect 17891 8585 17903 8619
rect 17937 8616 17949 8619
rect 18138 8616 18144 8628
rect 17937 8588 18144 8616
rect 17937 8585 17949 8588
rect 17891 8579 17949 8585
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 21910 8616 21916 8628
rect 18708 8588 21916 8616
rect 15672 8520 15976 8548
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16850 8548 16856 8560
rect 16080 8520 16856 8548
rect 16080 8508 16086 8520
rect 16850 8508 16856 8520
rect 16908 8508 16914 8560
rect 17681 8551 17739 8557
rect 17681 8517 17693 8551
rect 17727 8548 17739 8551
rect 17770 8548 17776 8560
rect 17727 8520 17776 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 17770 8508 17776 8520
rect 17828 8508 17834 8560
rect 18708 8557 18736 8588
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 22005 8619 22063 8625
rect 22005 8585 22017 8619
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 17972 8520 18705 8548
rect 11020 8452 12434 8480
rect 11020 8440 11026 8452
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13504 8452 13553 8480
rect 13504 8440 13510 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9640 8384 9781 8412
rect 9640 8372 9646 8384
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 10836 8384 11713 8412
rect 10836 8372 10842 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 13556 8412 13584 8443
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14458 8489 14464 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 13688 8452 14289 8480
rect 13688 8440 13694 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14425 8483 14464 8489
rect 14425 8449 14437 8483
rect 14425 8443 14464 8449
rect 14458 8440 14464 8443
rect 14516 8440 14522 8492
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 14783 8483 14841 8489
rect 14783 8449 14795 8483
rect 14829 8449 14841 8483
rect 14783 8443 14841 8449
rect 14182 8412 14188 8424
rect 13556 8384 14188 8412
rect 11701 8375 11759 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14798 8412 14826 8443
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 17972 8480 18000 8520
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 18693 8511 18751 8517
rect 18877 8551 18935 8557
rect 18877 8517 18889 8551
rect 18923 8548 18935 8551
rect 22020 8548 22048 8579
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 24489 8619 24547 8625
rect 24489 8616 24501 8619
rect 22152 8588 24501 8616
rect 22152 8576 22158 8588
rect 24489 8585 24501 8588
rect 24535 8585 24547 8619
rect 24489 8579 24547 8585
rect 25222 8557 25228 8560
rect 23354 8551 23412 8557
rect 23354 8548 23366 8551
rect 18923 8520 20392 8548
rect 22020 8520 23366 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 15344 8452 18000 8480
rect 18509 8483 18567 8489
rect 15344 8440 15350 8452
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18782 8480 18788 8492
rect 18555 8452 18788 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18782 8440 18788 8452
rect 18840 8480 18846 8492
rect 19334 8480 19340 8492
rect 18840 8452 19340 8480
rect 18840 8440 18846 8452
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 20364 8489 20392 8520
rect 23354 8517 23366 8520
rect 23400 8517 23412 8551
rect 25216 8548 25228 8557
rect 25183 8520 25228 8548
rect 23354 8511 23412 8517
rect 25216 8511 25228 8520
rect 25222 8508 25228 8511
rect 25280 8508 25286 8560
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20680 8452 21005 8480
rect 20680 8440 20686 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 20993 8443 21051 8449
rect 22066 8452 22201 8480
rect 15930 8412 15936 8424
rect 14798 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17862 8412 17868 8424
rect 16724 8384 17868 8412
rect 16724 8372 16730 8384
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8412 19763 8415
rect 22066 8412 22094 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 19751 8384 22094 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 23106 8412 23112 8424
rect 22336 8384 23112 8412
rect 22336 8372 22342 8384
rect 23106 8372 23112 8384
rect 23164 8372 23170 8424
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 24949 8415 25007 8421
rect 24949 8412 24961 8415
rect 24728 8384 24961 8412
rect 24728 8372 24734 8384
rect 24949 8381 24961 8384
rect 24995 8381 25007 8415
rect 24949 8375 25007 8381
rect 9079 8316 9444 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 14458 8344 14464 8356
rect 13228 8316 14464 8344
rect 13228 8304 13234 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 14568 8316 18184 8344
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 4120 8248 4261 8276
rect 4120 8236 4126 8248
rect 4249 8245 4261 8248
rect 4295 8276 4307 8279
rect 6362 8276 6368 8288
rect 4295 8248 6368 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 11146 8276 11152 8288
rect 7892 8248 11152 8276
rect 7892 8236 7898 8248
rect 11146 8236 11152 8248
rect 11204 8276 11210 8288
rect 12618 8276 12624 8288
rect 11204 8248 12624 8276
rect 11204 8236 11210 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13538 8276 13544 8288
rect 12952 8248 13544 8276
rect 12952 8236 12958 8248
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 13725 8279 13783 8285
rect 13725 8276 13737 8279
rect 13596 8248 13737 8276
rect 13596 8236 13602 8248
rect 13725 8245 13737 8248
rect 13771 8276 13783 8279
rect 14568 8276 14596 8316
rect 13771 8248 14596 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 15562 8236 15568 8288
rect 15620 8236 15626 8288
rect 16758 8236 16764 8288
rect 16816 8276 16822 8288
rect 17037 8279 17095 8285
rect 17037 8276 17049 8279
rect 16816 8248 17049 8276
rect 16816 8236 16822 8248
rect 17037 8245 17049 8248
rect 17083 8245 17095 8279
rect 17037 8239 17095 8245
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17865 8279 17923 8285
rect 17865 8276 17877 8279
rect 17460 8248 17877 8276
rect 17460 8236 17466 8248
rect 17865 8245 17877 8248
rect 17911 8245 17923 8279
rect 17865 8239 17923 8245
rect 18046 8236 18052 8288
rect 18104 8236 18110 8288
rect 18156 8276 18184 8316
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 19794 8344 19800 8356
rect 19392 8316 19800 8344
rect 19392 8304 19398 8316
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 20162 8304 20168 8356
rect 20220 8304 20226 8356
rect 20809 8347 20867 8353
rect 20809 8313 20821 8347
rect 20855 8344 20867 8347
rect 20855 8316 23152 8344
rect 20855 8313 20867 8316
rect 20809 8307 20867 8313
rect 19426 8276 19432 8288
rect 18156 8248 19432 8276
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 21082 8276 21088 8288
rect 19576 8248 21088 8276
rect 19576 8236 19582 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 21542 8276 21548 8288
rect 21232 8248 21548 8276
rect 21232 8236 21238 8248
rect 21542 8236 21548 8248
rect 21600 8236 21606 8288
rect 23124 8276 23152 8316
rect 26326 8304 26332 8356
rect 26384 8304 26390 8356
rect 23474 8276 23480 8288
rect 23124 8248 23480 8276
rect 23474 8236 23480 8248
rect 23532 8236 23538 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4396 8044 4445 8072
rect 4396 8032 4402 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 6917 8075 6975 8081
rect 4948 8044 6868 8072
rect 4948 8032 4954 8044
rect 6178 8004 6184 8016
rect 5920 7976 6184 8004
rect 1670 7896 1676 7948
rect 1728 7896 1734 7948
rect 5626 7936 5632 7948
rect 4632 7908 5632 7936
rect 1940 7871 1998 7877
rect 1940 7837 1952 7871
rect 1986 7868 1998 7871
rect 2314 7868 2320 7880
rect 1986 7840 2320 7868
rect 1986 7837 1998 7840
rect 1940 7831 1998 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 4632 7877 4660 7908
rect 5626 7896 5632 7908
rect 5684 7936 5690 7948
rect 5684 7908 5856 7936
rect 5684 7896 5690 7908
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 4948 7840 5212 7868
rect 4948 7828 4954 7840
rect 5184 7800 5212 7840
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5316 7840 5549 7868
rect 5316 7828 5322 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 5828 7877 5856 7908
rect 5920 7877 5948 7976
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 6840 8004 6868 8044
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7098 8072 7104 8084
rect 6963 8044 7104 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 8754 8072 8760 8084
rect 7484 8044 8760 8072
rect 7484 8004 7512 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9582 8072 9588 8084
rect 9180 8044 9588 8072
rect 9180 8032 9186 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10410 8032 10416 8084
rect 10468 8032 10474 8084
rect 10686 8032 10692 8084
rect 10744 8072 10750 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 10744 8044 11897 8072
rect 10744 8032 10750 8044
rect 11885 8041 11897 8044
rect 11931 8041 11943 8075
rect 11885 8035 11943 8041
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 13630 8072 13636 8084
rect 12115 8044 13636 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 15102 8032 15108 8084
rect 15160 8072 15166 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15160 8044 15669 8072
rect 15160 8032 15166 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 18046 8072 18052 8084
rect 15979 8044 18052 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18782 8072 18788 8084
rect 18564 8044 18788 8072
rect 18564 8032 18570 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 19150 8032 19156 8084
rect 19208 8072 19214 8084
rect 19518 8072 19524 8084
rect 19208 8044 19524 8072
rect 19208 8032 19214 8044
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 20530 8072 20536 8084
rect 19659 8044 20536 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20772 8044 21496 8072
rect 20772 8032 20778 8044
rect 6840 7976 7512 8004
rect 7484 7945 7512 7976
rect 7834 7964 7840 8016
rect 7892 7964 7898 8016
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 11974 8004 11980 8016
rect 9907 7976 11980 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 16022 8004 16028 8016
rect 12406 7976 16028 8004
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 9953 7939 10011 7945
rect 9953 7936 9965 7939
rect 7469 7899 7527 7905
rect 8588 7908 9965 7936
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 5920 7800 5948 7831
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 8588 7877 8616 7908
rect 9953 7905 9965 7908
rect 9999 7905 10011 7939
rect 12406 7936 12434 7976
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 16117 8007 16175 8013
rect 16117 7973 16129 8007
rect 16163 8004 16175 8007
rect 16206 8004 16212 8016
rect 16163 7976 16212 8004
rect 16163 7973 16175 7976
rect 16117 7967 16175 7973
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 19797 8007 19855 8013
rect 19797 8004 19809 8007
rect 18012 7976 19809 8004
rect 18012 7964 18018 7976
rect 19797 7973 19809 7976
rect 19843 7973 19855 8007
rect 21468 8004 21496 8044
rect 21542 8032 21548 8084
rect 21600 8072 21606 8084
rect 23106 8072 23112 8084
rect 21600 8044 23112 8072
rect 21600 8032 21606 8044
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 23293 8075 23351 8081
rect 23293 8041 23305 8075
rect 23339 8072 23351 8075
rect 24854 8072 24860 8084
rect 23339 8044 24860 8072
rect 23339 8041 23351 8044
rect 23293 8035 23351 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 24964 8044 26740 8072
rect 22741 8007 22799 8013
rect 22741 8004 22753 8007
rect 21468 7976 22753 8004
rect 19797 7967 19855 7973
rect 22741 7973 22753 7976
rect 22787 8004 22799 8007
rect 24964 8004 24992 8044
rect 22787 7976 24992 8004
rect 26712 8004 26740 8044
rect 27154 8032 27160 8084
rect 27212 8032 27218 8084
rect 28350 8004 28356 8016
rect 26712 7976 28356 8004
rect 22787 7973 22799 7976
rect 22741 7967 22799 7973
rect 28350 7964 28356 7976
rect 28408 7964 28414 8016
rect 9953 7899 10011 7905
rect 11716 7908 12434 7936
rect 12805 7939 12863 7945
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6052 7840 6745 7868
rect 6052 7828 6058 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9456 7840 9674 7868
rect 9456 7828 9462 7840
rect 5184 7772 5948 7800
rect 6546 7760 6552 7812
rect 6604 7760 6610 7812
rect 8754 7760 8760 7812
rect 8812 7800 8818 7812
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 8812 7772 9505 7800
rect 8812 7760 8818 7772
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 9646 7800 9674 7840
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11204 7840 11253 7868
rect 11204 7828 11210 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11716 7809 11744 7908
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 15838 7936 15844 7948
rect 12851 7908 15844 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16666 7936 16672 7948
rect 15988 7908 16672 7936
rect 15988 7896 15994 7908
rect 13078 7868 13084 7880
rect 11808 7840 13084 7868
rect 11701 7803 11759 7809
rect 9646 7772 11376 7800
rect 9493 7763 9551 7769
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 5258 7732 5264 7744
rect 4847 7704 5264 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 6089 7735 6147 7741
rect 6089 7701 6101 7735
rect 6135 7732 6147 7735
rect 7374 7732 7380 7744
rect 6135 7704 7380 7732
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 7742 7692 7748 7744
rect 7800 7732 7806 7744
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7800 7704 7941 7732
rect 7800 7692 7806 7704
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 7929 7695 7987 7701
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7732 8447 7735
rect 9582 7732 9588 7744
rect 8435 7704 9588 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11238 7732 11244 7744
rect 11103 7704 11244 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11348 7732 11376 7772
rect 11701 7769 11713 7803
rect 11747 7769 11759 7803
rect 11701 7763 11759 7769
rect 11808 7732 11836 7840
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 11917 7803 11975 7809
rect 11917 7769 11929 7803
rect 11963 7800 11975 7803
rect 12158 7800 12164 7812
rect 11963 7772 12164 7800
rect 11963 7769 11975 7772
rect 11917 7763 11975 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 12621 7803 12679 7809
rect 12621 7769 12633 7803
rect 12667 7800 12679 7803
rect 12802 7800 12808 7812
rect 12667 7772 12808 7800
rect 12667 7769 12679 7772
rect 12621 7763 12679 7769
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 13740 7800 13768 7831
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 14240 7840 14289 7868
rect 14240 7828 14246 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 15514 7840 15976 7868
rect 15514 7800 15542 7840
rect 13740 7772 15542 7800
rect 15948 7800 15976 7840
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16408 7877 16436 7908
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 18923 7908 20668 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 16172 7840 16221 7868
rect 16172 7828 16178 7840
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16482 7828 16488 7880
rect 16540 7868 16546 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 16540 7840 17601 7868
rect 16540 7828 16546 7840
rect 17589 7837 17601 7840
rect 17635 7868 17647 7871
rect 18693 7871 18751 7877
rect 17635 7840 18644 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17126 7800 17132 7812
rect 15948 7772 17132 7800
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 17405 7803 17463 7809
rect 17405 7769 17417 7803
rect 17451 7800 17463 7803
rect 18506 7800 18512 7812
rect 17451 7772 18512 7800
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 11348 7704 11836 7732
rect 13538 7692 13544 7744
rect 13596 7692 13602 7744
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 13688 7704 14657 7732
rect 13688 7692 13694 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 17420 7732 17448 7763
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 18616 7800 18644 7840
rect 18693 7837 18705 7871
rect 18739 7868 18751 7871
rect 19610 7868 19616 7880
rect 18739 7840 19616 7868
rect 18739 7837 18751 7840
rect 18693 7831 18751 7837
rect 19610 7828 19616 7840
rect 19668 7868 19674 7880
rect 19886 7868 19892 7880
rect 19668 7840 19892 7868
rect 19668 7828 19674 7840
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20036 7840 20545 7868
rect 20036 7828 20042 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20640 7868 20668 7908
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 22373 7939 22431 7945
rect 22373 7936 22385 7939
rect 21600 7908 22385 7936
rect 21600 7896 21606 7908
rect 22373 7905 22385 7908
rect 22419 7905 22431 7939
rect 22373 7899 22431 7905
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 25130 7936 25136 7948
rect 22520 7908 25136 7936
rect 22520 7896 22526 7908
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 22554 7868 22560 7880
rect 20640 7840 22560 7868
rect 20533 7831 20591 7837
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 23477 7871 23535 7877
rect 23477 7837 23489 7871
rect 23523 7868 23535 7871
rect 23842 7868 23848 7880
rect 23523 7840 23848 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 23992 7840 24777 7868
rect 23992 7828 23998 7840
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7868 25835 7871
rect 26418 7868 26424 7880
rect 25823 7840 26424 7868
rect 25823 7837 25835 7840
rect 25777 7831 25835 7837
rect 26418 7828 26424 7840
rect 26476 7828 26482 7880
rect 18616 7772 19012 7800
rect 15896 7704 17448 7732
rect 17773 7735 17831 7741
rect 15896 7692 15902 7704
rect 17773 7701 17785 7735
rect 17819 7732 17831 7735
rect 18874 7732 18880 7744
rect 17819 7704 18880 7732
rect 17819 7701 17831 7704
rect 17773 7695 17831 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 18984 7732 19012 7772
rect 19426 7760 19432 7812
rect 19484 7760 19490 7812
rect 19536 7772 19748 7800
rect 19536 7732 19564 7772
rect 18984 7704 19564 7732
rect 19610 7692 19616 7744
rect 19668 7741 19674 7744
rect 19668 7735 19687 7741
rect 19675 7701 19687 7735
rect 19720 7732 19748 7772
rect 20622 7760 20628 7812
rect 20680 7800 20686 7812
rect 20778 7803 20836 7809
rect 20778 7800 20790 7803
rect 20680 7772 20790 7800
rect 20680 7760 20686 7772
rect 20778 7769 20790 7772
rect 20824 7769 20836 7803
rect 24486 7800 24492 7812
rect 20778 7763 20836 7769
rect 20916 7772 24492 7800
rect 20916 7732 20944 7772
rect 24486 7760 24492 7772
rect 24544 7760 24550 7812
rect 26022 7803 26080 7809
rect 26022 7800 26034 7803
rect 24596 7772 26034 7800
rect 19720 7704 20944 7732
rect 19668 7695 19687 7701
rect 19668 7692 19674 7695
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 21600 7704 21925 7732
rect 21600 7692 21606 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 21913 7695 21971 7701
rect 22833 7735 22891 7741
rect 22833 7701 22845 7735
rect 22879 7732 22891 7735
rect 23198 7732 23204 7744
rect 22879 7704 23204 7732
rect 22879 7701 22891 7704
rect 22833 7695 22891 7701
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 24596 7741 24624 7772
rect 26022 7769 26034 7772
rect 26068 7769 26080 7803
rect 26022 7763 26080 7769
rect 24581 7735 24639 7741
rect 24581 7701 24593 7735
rect 24627 7701 24639 7735
rect 24581 7695 24639 7701
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 5534 7528 5540 7540
rect 3191 7500 5540 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6270 7528 6276 7540
rect 5951 7500 6276 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 7064 7500 7113 7528
rect 7064 7488 7070 7500
rect 7101 7497 7113 7500
rect 7147 7497 7159 7531
rect 9030 7528 9036 7540
rect 7101 7491 7159 7497
rect 7208 7500 9036 7528
rect 1670 7420 1676 7472
rect 1728 7460 1734 7472
rect 1728 7432 2774 7460
rect 1728 7420 1734 7432
rect 1780 7401 1808 7432
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 2021 7395 2079 7401
rect 2021 7392 2033 7395
rect 1765 7355 1823 7361
rect 1872 7364 2033 7392
rect 750 7284 756 7336
rect 808 7324 814 7336
rect 1872 7324 1900 7364
rect 2021 7361 2033 7364
rect 2067 7361 2079 7395
rect 2746 7392 2774 7432
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 6914 7460 6920 7472
rect 5316 7432 6920 7460
rect 5316 7420 5322 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 3970 7401 3976 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 2746 7364 3709 7392
rect 2021 7355 2079 7361
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3964 7355 3976 7401
rect 3970 7352 3976 7355
rect 4028 7352 4034 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5684 7364 5733 7392
rect 5684 7352 5690 7364
rect 5721 7361 5733 7364
rect 5767 7392 5779 7395
rect 5767 7364 6408 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 808 7296 1900 7324
rect 808 7284 814 7296
rect 4706 7216 4712 7268
rect 4764 7256 4770 7268
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 4764 7228 5089 7256
rect 4764 7216 4770 7228
rect 5077 7225 5089 7228
rect 5123 7225 5135 7259
rect 5077 7219 5135 7225
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 4724 7188 4752 7216
rect 3752 7160 4752 7188
rect 6380 7188 6408 7364
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6696 7364 6837 7392
rect 6696 7352 6702 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6512 7296 6929 7324
rect 6512 7284 6518 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 7116 7256 7144 7287
rect 6788 7228 7144 7256
rect 6788 7216 6794 7228
rect 7208 7188 7236 7500
rect 9030 7488 9036 7500
rect 9088 7528 9094 7540
rect 12802 7528 12808 7540
rect 9088 7500 12808 7528
rect 9088 7488 9094 7500
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 16022 7528 16028 7540
rect 13311 7500 16028 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 17000 7500 17325 7528
rect 17000 7488 17006 7500
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 17313 7491 17371 7497
rect 18138 7488 18144 7540
rect 18196 7528 18202 7540
rect 18995 7531 19053 7537
rect 18995 7528 19007 7531
rect 18196 7500 19007 7528
rect 18196 7488 18202 7500
rect 18995 7497 19007 7500
rect 19041 7528 19053 7531
rect 19610 7528 19616 7540
rect 19041 7500 19616 7528
rect 19041 7497 19053 7500
rect 18995 7491 19053 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20533 7531 20591 7537
rect 20533 7497 20545 7531
rect 20579 7528 20591 7531
rect 20622 7528 20628 7540
rect 20579 7500 20628 7528
rect 20579 7497 20591 7500
rect 20533 7491 20591 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 20956 7500 21496 7528
rect 20956 7488 20962 7500
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 7340 7432 9536 7460
rect 7340 7420 7346 7432
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 7524 7364 7573 7392
rect 7524 7352 7530 7364
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7708 7364 7757 7392
rect 7708 7352 7714 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9381 7395 9439 7401
rect 9381 7392 9393 7395
rect 8444 7364 9393 7392
rect 8444 7352 8450 7364
rect 9381 7361 9393 7364
rect 9427 7361 9439 7395
rect 9508 7392 9536 7432
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 9732 7432 12434 7460
rect 9732 7420 9738 7432
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 9508 7364 11161 7392
rect 9381 7355 9439 7361
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12250 7392 12256 7404
rect 11931 7364 12256 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12406 7392 12434 7432
rect 12894 7420 12900 7472
rect 12952 7420 12958 7472
rect 13113 7463 13171 7469
rect 13113 7429 13125 7463
rect 13159 7460 13171 7463
rect 14642 7460 14648 7472
rect 13159 7432 14648 7460
rect 13159 7429 13171 7432
rect 13113 7423 13171 7429
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 14826 7420 14832 7472
rect 14884 7460 14890 7472
rect 14884 7432 16252 7460
rect 14884 7420 14890 7432
rect 14441 7395 14499 7401
rect 14441 7392 14453 7395
rect 12406 7364 14453 7392
rect 14441 7361 14453 7364
rect 14487 7361 14499 7395
rect 14441 7355 14499 7361
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 15068 7364 16129 7392
rect 15068 7352 15074 7364
rect 16117 7361 16129 7364
rect 16163 7361 16175 7395
rect 16224 7392 16252 7432
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 17954 7460 17960 7472
rect 16448 7432 17960 7460
rect 16448 7420 16454 7432
rect 17954 7420 17960 7432
rect 18012 7460 18018 7472
rect 18012 7432 18092 7460
rect 18012 7420 18018 7432
rect 17589 7395 17647 7401
rect 17589 7392 17601 7395
rect 16224 7364 17601 7392
rect 16117 7355 16175 7361
rect 17589 7361 17601 7364
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 8168 7296 8217 7324
rect 8168 7284 8174 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 9122 7284 9128 7336
rect 9180 7284 9186 7336
rect 14182 7284 14188 7336
rect 14240 7284 14246 7336
rect 16132 7324 16160 7355
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18064 7401 18092 7432
rect 18782 7420 18788 7472
rect 18840 7420 18846 7472
rect 19886 7420 19892 7472
rect 19944 7460 19950 7472
rect 21468 7460 21496 7500
rect 21726 7488 21732 7540
rect 21784 7528 21790 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 21784 7500 22201 7528
rect 21784 7488 21790 7500
rect 22189 7497 22201 7500
rect 22235 7528 22247 7531
rect 22278 7528 22284 7540
rect 22235 7500 22284 7528
rect 22235 7497 22247 7500
rect 22189 7491 22247 7497
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 22738 7488 22744 7540
rect 22796 7488 22802 7540
rect 25961 7531 26019 7537
rect 25961 7528 25973 7531
rect 22848 7500 25973 7528
rect 22848 7460 22876 7500
rect 25961 7497 25973 7500
rect 26007 7497 26019 7531
rect 25961 7491 26019 7497
rect 19944 7432 21404 7460
rect 21468 7432 22876 7460
rect 19944 7420 19950 7432
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 19150 7392 19156 7404
rect 18656 7364 19156 7392
rect 18656 7352 18662 7364
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19978 7392 19984 7404
rect 19484 7364 19984 7392
rect 19484 7352 19490 7364
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20714 7352 20720 7404
rect 20772 7352 20778 7404
rect 21376 7401 21404 7432
rect 23474 7420 23480 7472
rect 23532 7460 23538 7472
rect 24826 7463 24884 7469
rect 24826 7460 24838 7463
rect 23532 7432 24838 7460
rect 23532 7420 23538 7432
rect 24826 7429 24838 7432
rect 24872 7429 24884 7463
rect 24826 7423 24884 7429
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7392 22155 7395
rect 22186 7392 22192 7404
rect 22143 7364 22192 7392
rect 22143 7361 22155 7364
rect 22097 7355 22155 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 22925 7395 22983 7401
rect 22925 7392 22937 7395
rect 22704 7364 22937 7392
rect 22704 7352 22710 7364
rect 22925 7361 22937 7364
rect 22971 7361 22983 7395
rect 22925 7355 22983 7361
rect 23198 7352 23204 7404
rect 23256 7392 23262 7404
rect 23569 7395 23627 7401
rect 23569 7392 23581 7395
rect 23256 7364 23581 7392
rect 23256 7352 23262 7364
rect 23569 7361 23581 7364
rect 23615 7361 23627 7395
rect 23569 7355 23627 7361
rect 24670 7352 24676 7404
rect 24728 7352 24734 7404
rect 17681 7327 17739 7333
rect 16132 7296 17632 7324
rect 8478 7216 8484 7268
rect 8536 7256 8542 7268
rect 8536 7228 8892 7256
rect 8536 7216 8542 7228
rect 6380 7160 7236 7188
rect 3752 7148 3758 7160
rect 7650 7148 7656 7200
rect 7708 7148 7714 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8628 7160 8677 7188
rect 8628 7148 8634 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8864 7188 8892 7228
rect 10502 7216 10508 7268
rect 10560 7216 10566 7268
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 17604 7256 17632 7296
rect 17681 7293 17693 7327
rect 17727 7324 17739 7327
rect 18230 7324 18236 7336
rect 17727 7296 18236 7324
rect 17727 7293 17739 7296
rect 17681 7287 17739 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 19610 7284 19616 7336
rect 19668 7284 19674 7336
rect 22278 7324 22284 7336
rect 19904 7296 22284 7324
rect 17773 7259 17831 7265
rect 15344 7228 16160 7256
rect 17604 7228 17724 7256
rect 15344 7216 15350 7228
rect 16132 7200 16160 7228
rect 9490 7188 9496 7200
rect 8864 7160 9496 7188
rect 8665 7151 8723 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10468 7160 10977 7188
rect 10468 7148 10474 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 11698 7148 11704 7200
rect 11756 7148 11762 7200
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 15565 7191 15623 7197
rect 15565 7188 15577 7191
rect 14424 7160 15577 7188
rect 14424 7148 14430 7160
rect 15565 7157 15577 7160
rect 15611 7157 15623 7191
rect 15565 7151 15623 7157
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16172 7160 16221 7188
rect 16172 7148 16178 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 17696 7188 17724 7228
rect 17773 7225 17785 7259
rect 17819 7256 17831 7259
rect 19153 7259 19211 7265
rect 19153 7256 19165 7259
rect 17819 7228 19165 7256
rect 17819 7225 17831 7228
rect 17773 7219 17831 7225
rect 19153 7225 19165 7228
rect 19199 7225 19211 7259
rect 19153 7219 19211 7225
rect 18230 7188 18236 7200
rect 17696 7160 18236 7188
rect 16209 7151 16267 7157
rect 18230 7148 18236 7160
rect 18288 7188 18294 7200
rect 18598 7188 18604 7200
rect 18288 7160 18604 7188
rect 18288 7148 18294 7160
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18969 7191 19027 7197
rect 18969 7157 18981 7191
rect 19015 7188 19027 7191
rect 19904 7188 19932 7296
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22554 7284 22560 7336
rect 22612 7324 22618 7336
rect 23750 7324 23756 7336
rect 22612 7296 23756 7324
rect 22612 7284 22618 7296
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 24581 7327 24639 7333
rect 24581 7293 24593 7327
rect 24627 7324 24639 7327
rect 24688 7324 24716 7352
rect 24627 7296 24716 7324
rect 24627 7293 24639 7296
rect 24581 7287 24639 7293
rect 19978 7216 19984 7268
rect 20036 7216 20042 7268
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 21542 7256 21548 7268
rect 20588 7228 21548 7256
rect 20588 7216 20594 7228
rect 21542 7216 21548 7228
rect 21600 7216 21606 7268
rect 23566 7256 23572 7268
rect 22066 7228 23572 7256
rect 19015 7160 19932 7188
rect 20073 7191 20131 7197
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 20073 7157 20085 7191
rect 20119 7188 20131 7191
rect 20254 7188 20260 7200
rect 20119 7160 20260 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 21177 7191 21235 7197
rect 21177 7157 21189 7191
rect 21223 7188 21235 7191
rect 22066 7188 22094 7228
rect 23566 7216 23572 7228
rect 23624 7216 23630 7268
rect 26510 7256 26516 7268
rect 25884 7228 26516 7256
rect 21223 7160 22094 7188
rect 23385 7191 23443 7197
rect 21223 7157 21235 7160
rect 21177 7151 21235 7157
rect 23385 7157 23397 7191
rect 23431 7188 23443 7191
rect 25884 7188 25912 7228
rect 26510 7216 26516 7228
rect 26568 7216 26574 7268
rect 23431 7160 25912 7188
rect 23431 7157 23443 7160
rect 23385 7151 23443 7157
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 4617 6987 4675 6993
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 4890 6984 4896 6996
rect 4663 6956 4896 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 8386 6944 8392 6996
rect 8444 6944 8450 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9214 6984 9220 6996
rect 8812 6956 9220 6984
rect 8812 6944 8818 6956
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 9950 6984 9956 6996
rect 9907 6956 9956 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 11977 6987 12035 6993
rect 11977 6984 11989 6987
rect 10560 6956 11989 6984
rect 10560 6944 10566 6956
rect 11977 6953 11989 6956
rect 12023 6953 12035 6987
rect 11977 6947 12035 6953
rect 12158 6944 12164 6996
rect 12216 6944 12222 6996
rect 12621 6987 12679 6993
rect 12621 6953 12633 6987
rect 12667 6984 12679 6987
rect 12710 6984 12716 6996
rect 12667 6956 12716 6984
rect 12667 6953 12679 6956
rect 12621 6947 12679 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13504 6956 14412 6984
rect 13504 6944 13510 6956
rect 4801 6919 4859 6925
rect 4801 6916 4813 6919
rect 4172 6888 4813 6916
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 4172 6848 4200 6888
rect 4801 6885 4813 6888
rect 4847 6916 4859 6919
rect 6733 6919 6791 6925
rect 4847 6888 5856 6916
rect 4847 6885 4859 6888
rect 4801 6879 4859 6885
rect 5718 6848 5724 6860
rect 3292 6820 4200 6848
rect 4264 6820 5724 6848
rect 3292 6808 3298 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 1670 6780 1676 6792
rect 1627 6752 1676 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 4264 6789 4292 6820
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5828 6848 5856 6888
rect 6733 6885 6745 6919
rect 6779 6885 6791 6919
rect 6733 6879 6791 6885
rect 6748 6848 6776 6879
rect 10962 6876 10968 6928
rect 11020 6876 11026 6928
rect 12894 6916 12900 6928
rect 11809 6888 12900 6916
rect 7466 6848 7472 6860
rect 5828 6820 6500 6848
rect 6748 6820 7472 6848
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5258 6780 5264 6792
rect 4663 6752 5264 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5552 6752 6377 6780
rect 842 6672 848 6724
rect 900 6712 906 6724
rect 1826 6715 1884 6721
rect 1826 6712 1838 6715
rect 900 6684 1838 6712
rect 900 6672 906 6684
rect 1826 6681 1838 6684
rect 1872 6681 1884 6715
rect 1826 6675 1884 6681
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5552 6721 5580 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6472 6780 6500 6820
rect 7466 6808 7472 6820
rect 7524 6848 7530 6860
rect 9766 6848 9772 6860
rect 7524 6820 9772 6848
rect 7524 6808 7530 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 10980 6848 11008 6876
rect 10888 6820 11008 6848
rect 7190 6780 7196 6792
rect 6472 6752 7196 6780
rect 6365 6743 6423 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7800 6752 7941 6780
rect 7800 6740 7806 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 10686 6789 10692 6792
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 9272 6752 10517 6780
rect 9272 6740 9278 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10653 6783 10692 6789
rect 10653 6749 10665 6783
rect 10653 6743 10692 6749
rect 10686 6740 10692 6743
rect 10744 6740 10750 6792
rect 10888 6789 10916 6820
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11011 6783 11069 6789
rect 11011 6749 11023 6783
rect 11057 6780 11069 6783
rect 11238 6780 11244 6792
rect 11057 6752 11244 6780
rect 11057 6749 11069 6752
rect 11011 6743 11069 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 4856 6684 5549 6712
rect 4856 6672 4862 6684
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 5537 6675 5595 6681
rect 5721 6715 5779 6721
rect 5721 6681 5733 6715
rect 5767 6712 5779 6715
rect 5767 6684 6408 6712
rect 5767 6681 5779 6684
rect 5721 6675 5779 6681
rect 6380 6656 6408 6684
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 9306 6712 9312 6724
rect 8444 6684 9312 6712
rect 8444 6672 8450 6684
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 10318 6712 10324 6724
rect 9723 6684 10324 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 11809 6721 11837 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 13998 6916 14004 6928
rect 13004 6888 14004 6916
rect 13004 6848 13032 6888
rect 13998 6876 14004 6888
rect 14056 6876 14062 6928
rect 14384 6916 14412 6956
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 14516 6956 14657 6984
rect 14516 6944 14522 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 14826 6944 14832 6996
rect 14884 6944 14890 6996
rect 15470 6944 15476 6996
rect 15528 6944 15534 6996
rect 17034 6984 17040 6996
rect 15596 6956 17040 6984
rect 15010 6916 15016 6928
rect 14384 6888 15016 6916
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15102 6876 15108 6928
rect 15160 6916 15166 6928
rect 15596 6916 15624 6956
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17184 6956 17601 6984
rect 17184 6944 17190 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 20530 6984 20536 6996
rect 17589 6947 17647 6953
rect 18340 6956 20536 6984
rect 15160 6888 15624 6916
rect 15657 6919 15715 6925
rect 15160 6876 15166 6888
rect 15657 6885 15669 6919
rect 15703 6885 15715 6919
rect 15657 6879 15715 6885
rect 12176 6820 13032 6848
rect 13081 6851 13139 6857
rect 11793 6715 11851 6721
rect 11793 6681 11805 6715
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 12009 6715 12067 6721
rect 12009 6681 12021 6715
rect 12055 6712 12067 6715
rect 12176 6712 12204 6820
rect 13081 6817 13093 6851
rect 13127 6848 13139 6851
rect 15672 6848 15700 6879
rect 16482 6876 16488 6928
rect 16540 6876 16546 6928
rect 17218 6876 17224 6928
rect 17276 6916 17282 6928
rect 17405 6919 17463 6925
rect 17405 6916 17417 6919
rect 17276 6888 17417 6916
rect 17276 6876 17282 6888
rect 17405 6885 17417 6888
rect 17451 6916 17463 6919
rect 18340 6916 18368 6956
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 20714 6944 20720 6996
rect 20772 6984 20778 6996
rect 20809 6987 20867 6993
rect 20809 6984 20821 6987
rect 20772 6956 20821 6984
rect 20772 6944 20778 6956
rect 20809 6953 20821 6956
rect 20855 6953 20867 6987
rect 20809 6947 20867 6953
rect 23106 6944 23112 6996
rect 23164 6944 23170 6996
rect 17451 6888 18368 6916
rect 18417 6919 18475 6925
rect 17451 6885 17463 6888
rect 17405 6879 17463 6885
rect 18417 6885 18429 6919
rect 18463 6885 18475 6919
rect 18417 6879 18475 6885
rect 19705 6919 19763 6925
rect 19705 6885 19717 6919
rect 19751 6885 19763 6919
rect 19705 6879 19763 6885
rect 13127 6820 15700 6848
rect 18432 6848 18460 6879
rect 18690 6848 18696 6860
rect 18432 6820 18696 6848
rect 13127 6817 13139 6820
rect 13081 6811 13139 6817
rect 18690 6808 18696 6820
rect 18748 6848 18754 6860
rect 19150 6848 19156 6860
rect 18748 6820 19156 6848
rect 18748 6808 18754 6820
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19720 6848 19748 6879
rect 20622 6876 20628 6928
rect 20680 6876 20686 6928
rect 19300 6820 19748 6848
rect 19300 6808 19306 6820
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 20036 6820 20361 6848
rect 20036 6808 20042 6820
rect 20349 6817 20361 6820
rect 20395 6817 20407 6851
rect 20349 6811 20407 6817
rect 21726 6808 21732 6860
rect 21784 6808 21790 6860
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13630 6780 13636 6792
rect 13403 6752 13636 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 15102 6780 15108 6792
rect 14476 6752 15108 6780
rect 13280 6712 13308 6740
rect 12055 6684 12204 6712
rect 12406 6684 13308 6712
rect 12055 6681 12067 6684
rect 12009 6675 12067 6681
rect 2958 6604 2964 6656
rect 3016 6604 3022 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5626 6644 5632 6656
rect 4764 6616 5632 6644
rect 4764 6604 4770 6616
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5905 6647 5963 6653
rect 5905 6613 5917 6647
rect 5951 6644 5963 6647
rect 5994 6644 6000 6656
rect 5951 6616 6000 6644
rect 5951 6613 5963 6616
rect 5905 6607 5963 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6362 6604 6368 6656
rect 6420 6604 6426 6656
rect 6822 6604 6828 6656
rect 6880 6604 6886 6656
rect 7742 6604 7748 6656
rect 7800 6604 7806 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 9877 6647 9935 6653
rect 9877 6644 9889 6647
rect 9824 6616 9889 6644
rect 9824 6604 9830 6616
rect 9877 6613 9889 6616
rect 9923 6613 9935 6647
rect 9877 6607 9935 6613
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 11054 6644 11060 6656
rect 10091 6616 11060 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 12406 6644 12434 6684
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 14476 6721 14504 6752
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 15160 6752 15332 6780
rect 15160 6740 15166 6752
rect 15304 6721 15332 6752
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16850 6780 16856 6792
rect 15896 6752 16856 6780
rect 15896 6740 15902 6752
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18095 6752 20116 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 14461 6715 14519 6721
rect 14461 6712 14473 6715
rect 13780 6684 14473 6712
rect 13780 6672 13786 6684
rect 14461 6681 14473 6684
rect 14507 6681 14519 6715
rect 14461 6675 14519 6681
rect 15289 6715 15347 6721
rect 15289 6681 15301 6715
rect 15335 6681 15347 6715
rect 15289 6675 15347 6681
rect 15470 6672 15476 6724
rect 15528 6721 15534 6724
rect 15528 6715 15547 6721
rect 15535 6681 15547 6715
rect 15528 6675 15547 6681
rect 15528 6672 15534 6675
rect 16114 6672 16120 6724
rect 16172 6712 16178 6724
rect 17129 6715 17187 6721
rect 16172 6684 16712 6712
rect 16172 6672 16178 6684
rect 11195 6616 12434 6644
rect 13265 6647 13323 6653
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 14366 6644 14372 6656
rect 13311 6616 14372 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14642 6604 14648 6656
rect 14700 6653 14706 6656
rect 14700 6647 14719 6653
rect 14707 6613 14719 6647
rect 14700 6607 14719 6613
rect 14700 6604 14706 6607
rect 15654 6604 15660 6656
rect 15712 6644 15718 6656
rect 16577 6647 16635 6653
rect 16577 6644 16589 6647
rect 15712 6616 16589 6644
rect 15712 6604 15718 6616
rect 16577 6613 16589 6616
rect 16623 6613 16635 6647
rect 16684 6644 16712 6684
rect 17129 6681 17141 6715
rect 17175 6712 17187 6715
rect 17862 6712 17868 6724
rect 17175 6684 17868 6712
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 19334 6712 19340 6724
rect 17972 6684 19340 6712
rect 16942 6644 16948 6656
rect 16684 6616 16948 6644
rect 16577 6607 16635 6613
rect 16942 6604 16948 6616
rect 17000 6644 17006 6656
rect 17972 6644 18000 6684
rect 19334 6672 19340 6684
rect 19392 6712 19398 6724
rect 19429 6715 19487 6721
rect 19429 6712 19441 6715
rect 19392 6684 19441 6712
rect 19392 6672 19398 6684
rect 19429 6681 19441 6684
rect 19475 6681 19487 6715
rect 19429 6675 19487 6681
rect 17000 6616 18000 6644
rect 18509 6647 18567 6653
rect 17000 6604 17006 6616
rect 18509 6613 18521 6647
rect 18555 6644 18567 6647
rect 19518 6644 19524 6656
rect 18555 6616 19524 6644
rect 18555 6613 18567 6616
rect 18509 6607 18567 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 20088 6644 20116 6752
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 21985 6783 22043 6789
rect 21985 6780 21997 6783
rect 20220 6752 21997 6780
rect 20220 6740 20226 6752
rect 21985 6749 21997 6752
rect 22031 6749 22043 6783
rect 21985 6743 22043 6749
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24670 6780 24676 6792
rect 24627 6752 24676 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 24780 6752 26096 6780
rect 21634 6672 21640 6724
rect 21692 6712 21698 6724
rect 24780 6712 24808 6752
rect 21692 6684 24808 6712
rect 24848 6715 24906 6721
rect 21692 6672 21698 6684
rect 24848 6681 24860 6715
rect 24894 6712 24906 6715
rect 24946 6712 24952 6724
rect 24894 6684 24952 6712
rect 24894 6681 24906 6684
rect 24848 6675 24906 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 25130 6672 25136 6724
rect 25188 6712 25194 6724
rect 25188 6684 26004 6712
rect 25188 6672 25194 6684
rect 20714 6644 20720 6656
rect 20088 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 23569 6647 23627 6653
rect 23569 6613 23581 6647
rect 23615 6644 23627 6647
rect 24762 6644 24768 6656
rect 23615 6616 24768 6644
rect 23615 6613 23627 6616
rect 23569 6607 23627 6613
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 25976 6653 26004 6684
rect 25961 6647 26019 6653
rect 25961 6613 25973 6647
rect 26007 6613 26019 6647
rect 26068 6644 26096 6752
rect 26418 6740 26424 6792
rect 26476 6740 26482 6792
rect 26510 6740 26516 6792
rect 26568 6780 26574 6792
rect 26677 6783 26735 6789
rect 26677 6780 26689 6783
rect 26568 6752 26689 6780
rect 26568 6740 26574 6752
rect 26677 6749 26689 6752
rect 26723 6749 26735 6783
rect 26677 6743 26735 6749
rect 27801 6647 27859 6653
rect 27801 6644 27813 6647
rect 26068 6616 27813 6644
rect 25961 6607 26019 6613
rect 27801 6613 27813 6616
rect 27847 6613 27859 6647
rect 27801 6607 27859 6613
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 4614 6440 4620 6452
rect 4111 6412 4620 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 5258 6440 5264 6452
rect 4856 6412 5264 6440
rect 4856 6400 4862 6412
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5408 6412 5457 6440
rect 5408 6400 5414 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 8386 6440 8392 6452
rect 6420 6412 8392 6440
rect 6420 6400 6426 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9364 6412 12112 6440
rect 9364 6400 9370 6412
rect 3694 6332 3700 6384
rect 3752 6332 3758 6384
rect 3913 6375 3971 6381
rect 3913 6341 3925 6375
rect 3959 6372 3971 6375
rect 4338 6372 4344 6384
rect 3959 6344 4344 6372
rect 3959 6341 3971 6344
rect 3913 6335 3971 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 4706 6332 4712 6384
rect 4764 6332 4770 6384
rect 4982 6332 4988 6384
rect 5040 6372 5046 6384
rect 8849 6375 8907 6381
rect 5040 6344 5580 6372
rect 5040 6332 5046 6344
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1728 6276 1777 6304
rect 1728 6264 1734 6276
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2032 6307 2090 6313
rect 2032 6273 2044 6307
rect 2078 6304 2090 6307
rect 4246 6304 4252 6316
rect 2078 6276 4252 6304
rect 2078 6273 2090 6276
rect 2032 6267 2090 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4724 6304 4752 6332
rect 4356 6276 4752 6304
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 4356 6236 4384 6276
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5074 6304 5080 6316
rect 4948 6276 5080 6304
rect 4948 6264 4954 6276
rect 5074 6264 5080 6276
rect 5132 6304 5138 6316
rect 5552 6313 5580 6344
rect 8849 6341 8861 6375
rect 8895 6372 8907 6375
rect 8938 6372 8944 6384
rect 8895 6344 8944 6372
rect 8895 6341 8907 6344
rect 8849 6335 8907 6341
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 9065 6375 9123 6381
rect 9065 6341 9077 6375
rect 9111 6372 9123 6375
rect 9766 6372 9772 6384
rect 9111 6344 9772 6372
rect 9111 6341 9123 6344
rect 9065 6335 9123 6341
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 10042 6381 10048 6384
rect 10036 6372 10048 6381
rect 10003 6344 10048 6372
rect 10036 6335 10048 6344
rect 10042 6332 10048 6335
rect 10100 6332 10106 6384
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5132 6276 5365 6304
rect 5132 6264 5138 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 6730 6264 6736 6316
rect 6788 6264 6794 6316
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 8956 6304 8984 6332
rect 10318 6304 10324 6316
rect 8956 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11112 6276 11713 6304
rect 11112 6264 11118 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 12084 6313 12112 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 13354 6440 13360 6452
rect 12216 6412 13360 6440
rect 12216 6400 12222 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 15381 6443 15439 6449
rect 15381 6440 15393 6443
rect 15252 6412 15393 6440
rect 15252 6400 15258 6412
rect 15381 6409 15393 6412
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17586 6440 17592 6452
rect 17083 6412 17592 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 17920 6412 18337 6440
rect 17920 6400 17926 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 12434 6332 12440 6384
rect 12492 6372 12498 6384
rect 14093 6375 14151 6381
rect 14093 6372 14105 6375
rect 12492 6344 14105 6372
rect 12492 6332 12498 6344
rect 14093 6341 14105 6344
rect 14139 6372 14151 6375
rect 15286 6372 15292 6384
rect 14139 6344 15292 6372
rect 14139 6341 14151 6344
rect 14093 6335 14151 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 15657 6375 15715 6381
rect 15657 6372 15669 6375
rect 15396 6344 15669 6372
rect 11977 6307 12035 6313
rect 11848 6276 11893 6304
rect 11848 6264 11854 6276
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12207 6307 12265 6313
rect 12207 6273 12219 6307
rect 12253 6304 12265 6307
rect 12342 6304 12348 6316
rect 12253 6276 12348 6304
rect 12253 6273 12265 6276
rect 12207 6267 12265 6273
rect 3016 6208 4384 6236
rect 3016 6196 3022 6208
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 6512 6208 8309 6236
rect 6512 6196 6518 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9180 6208 9781 6236
rect 9180 6196 9186 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 11992 6236 12020 6267
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6304 12955 6307
rect 13446 6304 13452 6316
rect 12943 6276 13452 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 15396 6304 15424 6344
rect 15657 6341 15669 6344
rect 15703 6341 15715 6375
rect 15657 6335 15715 6341
rect 15887 6375 15945 6381
rect 15887 6341 15899 6375
rect 15933 6372 15945 6375
rect 16666 6372 16672 6384
rect 15933 6344 16672 6372
rect 15933 6341 15945 6344
rect 15887 6335 15945 6341
rect 16666 6332 16672 6344
rect 16724 6332 16730 6384
rect 17313 6375 17371 6381
rect 17313 6341 17325 6375
rect 17359 6372 17371 6375
rect 17678 6372 17684 6384
rect 17359 6344 17684 6372
rect 17359 6341 17371 6344
rect 17313 6335 17371 6341
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 18230 6332 18236 6384
rect 18288 6332 18294 6384
rect 18340 6372 18368 6403
rect 18966 6400 18972 6452
rect 19024 6440 19030 6452
rect 25130 6440 25136 6452
rect 19024 6412 25136 6440
rect 19024 6400 19030 6412
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 25280 6412 25452 6440
rect 25280 6400 25286 6412
rect 19610 6372 19616 6384
rect 18340 6344 19616 6372
rect 19610 6332 19616 6344
rect 19668 6372 19674 6384
rect 19978 6372 19984 6384
rect 19668 6344 19984 6372
rect 19668 6332 19674 6344
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 21358 6372 21364 6384
rect 20732 6344 21364 6372
rect 20732 6316 20760 6344
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 22094 6332 22100 6384
rect 22152 6372 22158 6384
rect 22830 6372 22836 6384
rect 22152 6344 22836 6372
rect 22152 6332 22158 6344
rect 22830 6332 22836 6344
rect 22888 6332 22894 6384
rect 23382 6332 23388 6384
rect 23440 6332 23446 6384
rect 15252 6276 15424 6304
rect 15252 6264 15258 6276
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15528 6276 15577 6304
rect 15528 6264 15534 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16264 6276 17233 6304
rect 16264 6264 16270 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17543 6307 17601 6313
rect 17543 6273 17555 6307
rect 17589 6304 17601 6307
rect 17954 6304 17960 6316
rect 17589 6276 17960 6304
rect 17589 6273 17601 6276
rect 17543 6267 17601 6273
rect 13630 6236 13636 6248
rect 10836 6208 12020 6236
rect 10836 6196 10842 6208
rect 3145 6171 3203 6177
rect 3145 6137 3157 6171
rect 3191 6168 3203 6171
rect 3191 6140 4292 6168
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 4264 6100 4292 6140
rect 4338 6128 4344 6180
rect 4396 6168 4402 6180
rect 4396 6140 9168 6168
rect 4396 6128 4402 6140
rect 4982 6100 4988 6112
rect 4264 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 5592 6072 6561 6100
rect 5592 6060 5598 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7374 6100 7380 6112
rect 7248 6072 7380 6100
rect 7248 6060 7254 6072
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8996 6072 9045 6100
rect 8996 6060 9002 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9140 6100 9168 6140
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 11149 6171 11207 6177
rect 11149 6168 11161 6171
rect 10928 6140 11161 6168
rect 10928 6128 10934 6140
rect 11149 6137 11161 6140
rect 11195 6137 11207 6171
rect 11992 6168 12020 6208
rect 12268 6208 13636 6236
rect 12268 6168 12296 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6236 14611 6239
rect 14826 6236 14832 6248
rect 14599 6208 14832 6236
rect 14599 6205 14611 6208
rect 14553 6199 14611 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15344 6208 16037 6236
rect 15344 6196 15350 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17126 6236 17132 6248
rect 16908 6208 17132 6236
rect 16908 6196 16914 6208
rect 17126 6196 17132 6208
rect 17184 6236 17190 6248
rect 17420 6236 17448 6267
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18748 6276 18889 6304
rect 18748 6264 18754 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 19058 6264 19064 6316
rect 19116 6264 19122 6316
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19300 6276 20208 6304
rect 19300 6264 19306 6276
rect 17184 6208 17448 6236
rect 17681 6239 17739 6245
rect 17184 6196 17190 6208
rect 17681 6205 17693 6239
rect 17727 6236 17739 6239
rect 19702 6236 19708 6248
rect 17727 6208 19708 6236
rect 17727 6205 17739 6208
rect 17681 6199 17739 6205
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 20180 6236 20208 6276
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 20714 6264 20720 6316
rect 20772 6264 20778 6316
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22244 6276 22293 6304
rect 22244 6264 22250 6276
rect 22281 6273 22293 6276
rect 22327 6304 22339 6307
rect 23198 6304 23204 6316
rect 22327 6276 23204 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 23198 6264 23204 6276
rect 23256 6304 23262 6316
rect 23400 6304 23428 6332
rect 23256 6276 23428 6304
rect 23256 6264 23262 6276
rect 24210 6264 24216 6316
rect 24268 6264 24274 6316
rect 25424 6304 25452 6412
rect 26602 6400 26608 6452
rect 26660 6400 26666 6452
rect 25481 6307 25539 6313
rect 25481 6304 25493 6307
rect 25424 6276 25493 6304
rect 25481 6273 25493 6276
rect 25527 6273 25539 6307
rect 25481 6267 25539 6273
rect 21082 6236 21088 6248
rect 20180 6208 21088 6236
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 22002 6236 22008 6248
rect 21324 6208 22008 6236
rect 21324 6196 21330 6208
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 25038 6236 25044 6248
rect 24728 6208 25044 6236
rect 24728 6196 24734 6208
rect 25038 6196 25044 6208
rect 25096 6236 25102 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25096 6208 25237 6236
rect 25096 6196 25102 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 11992 6140 12296 6168
rect 11149 6131 11207 6137
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13081 6171 13139 6177
rect 13081 6168 13093 6171
rect 12768 6140 13093 6168
rect 12768 6128 12774 6140
rect 13081 6137 13093 6140
rect 13127 6137 13139 6171
rect 13081 6131 13139 6137
rect 14461 6171 14519 6177
rect 14461 6137 14473 6171
rect 14507 6137 14519 6171
rect 14461 6131 14519 6137
rect 12158 6100 12164 6112
rect 9140 6072 12164 6100
rect 9033 6063 9091 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12345 6103 12403 6109
rect 12345 6069 12357 6103
rect 12391 6100 12403 6103
rect 14090 6100 14096 6112
rect 12391 6072 14096 6100
rect 12391 6069 12403 6072
rect 12345 6063 12403 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14476 6100 14504 6131
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 16206 6168 16212 6180
rect 14700 6140 16212 6168
rect 14700 6128 14706 6140
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 17586 6168 17592 6180
rect 17368 6140 17592 6168
rect 17368 6128 17374 6140
rect 17586 6128 17592 6140
rect 17644 6128 17650 6180
rect 18046 6128 18052 6180
rect 18104 6168 18110 6180
rect 20622 6168 20628 6180
rect 18104 6140 20628 6168
rect 18104 6128 18110 6140
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 20990 6128 20996 6180
rect 21048 6128 21054 6180
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 24210 6168 24216 6180
rect 21223 6140 24216 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 14550 6100 14556 6112
rect 14476 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6100 14614 6112
rect 17862 6100 17868 6112
rect 14608 6072 17868 6100
rect 14608 6060 14614 6072
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 18877 6103 18935 6109
rect 18877 6100 18889 6103
rect 18840 6072 18889 6100
rect 18840 6060 18846 6072
rect 18877 6069 18889 6072
rect 18923 6069 18935 6103
rect 18877 6063 18935 6069
rect 20073 6103 20131 6109
rect 20073 6069 20085 6103
rect 20119 6100 20131 6103
rect 23382 6100 23388 6112
rect 20119 6072 23388 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 23566 6100 23572 6112
rect 23523 6072 23572 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 24029 6103 24087 6109
rect 24029 6069 24041 6103
rect 24075 6100 24087 6103
rect 27062 6100 27068 6112
rect 24075 6072 27068 6100
rect 24075 6069 24087 6072
rect 24029 6063 24087 6069
rect 27062 6060 27068 6072
rect 27120 6060 27126 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 2958 5896 2964 5908
rect 2547 5868 2964 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3326 5896 3332 5908
rect 3099 5868 3332 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 6730 5896 6736 5908
rect 3896 5868 6736 5896
rect 1210 5788 1216 5840
rect 1268 5828 1274 5840
rect 3896 5828 3924 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 9766 5896 9772 5908
rect 7024 5868 9772 5896
rect 1268 5800 3924 5828
rect 3973 5831 4031 5837
rect 1268 5788 1274 5800
rect 3973 5797 3985 5831
rect 4019 5828 4031 5831
rect 4062 5828 4068 5840
rect 4019 5800 4068 5828
rect 4019 5797 4031 5800
rect 3973 5791 4031 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 7024 5837 7052 5868
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 10100 5868 11897 5896
rect 10100 5856 10106 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 12894 5896 12900 5908
rect 12115 5868 12900 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 14461 5899 14519 5905
rect 13044 5868 13492 5896
rect 13044 5856 13050 5868
rect 5537 5831 5595 5837
rect 5537 5828 5549 5831
rect 5500 5800 5549 5828
rect 5500 5788 5506 5800
rect 5537 5797 5549 5800
rect 5583 5797 5595 5831
rect 5537 5791 5595 5797
rect 7009 5831 7067 5837
rect 7009 5797 7021 5831
rect 7055 5797 7067 5831
rect 8202 5828 8208 5840
rect 7009 5791 7067 5797
rect 7116 5800 8208 5828
rect 566 5720 572 5772
rect 624 5760 630 5772
rect 624 5732 1808 5760
rect 624 5720 630 5732
rect 474 5652 480 5704
rect 532 5692 538 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 532 5664 1685 5692
rect 532 5652 538 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1780 5692 1808 5732
rect 1854 5720 1860 5772
rect 1912 5720 1918 5772
rect 7116 5760 7144 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8573 5831 8631 5837
rect 8573 5828 8585 5831
rect 8444 5800 8585 5828
rect 8444 5788 8450 5800
rect 8573 5797 8585 5800
rect 8619 5828 8631 5831
rect 9122 5828 9128 5840
rect 8619 5800 9128 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 9122 5788 9128 5800
rect 9180 5788 9186 5840
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10505 5831 10563 5837
rect 10505 5828 10517 5831
rect 10284 5800 10517 5828
rect 10284 5788 10290 5800
rect 10505 5797 10517 5800
rect 10551 5797 10563 5831
rect 10505 5791 10563 5797
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10928 5800 10977 5828
rect 10928 5788 10934 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 13464 5828 13492 5868
rect 14461 5865 14473 5899
rect 14507 5896 14519 5899
rect 17218 5896 17224 5908
rect 14507 5868 17224 5896
rect 14507 5865 14519 5868
rect 14461 5859 14519 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 21266 5896 21272 5908
rect 17420 5868 21272 5896
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 13464 5800 14657 5828
rect 10965 5791 11023 5797
rect 14645 5797 14657 5800
rect 14691 5797 14703 5831
rect 14645 5791 14703 5797
rect 15381 5831 15439 5837
rect 15381 5797 15393 5831
rect 15427 5828 15439 5831
rect 15746 5828 15752 5840
rect 15427 5800 15752 5828
rect 15427 5797 15439 5800
rect 15381 5791 15439 5797
rect 15746 5788 15752 5800
rect 15804 5828 15810 5840
rect 17420 5828 17448 5868
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 23109 5899 23167 5905
rect 23109 5896 23121 5899
rect 21744 5868 23121 5896
rect 15804 5800 17448 5828
rect 17497 5831 17555 5837
rect 15804 5788 15810 5800
rect 17497 5797 17509 5831
rect 17543 5828 17555 5831
rect 17586 5828 17592 5840
rect 17543 5800 17592 5828
rect 17543 5797 17555 5800
rect 17497 5791 17555 5797
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 20809 5831 20867 5837
rect 20809 5828 20821 5831
rect 20680 5800 20821 5828
rect 20680 5788 20686 5800
rect 20809 5797 20821 5800
rect 20855 5797 20867 5831
rect 20809 5791 20867 5797
rect 21082 5788 21088 5840
rect 21140 5828 21146 5840
rect 21744 5828 21772 5868
rect 23109 5865 23121 5868
rect 23155 5865 23167 5899
rect 23109 5859 23167 5865
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23934 5896 23940 5908
rect 23532 5868 23940 5896
rect 23532 5856 23538 5868
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 24486 5856 24492 5908
rect 24544 5896 24550 5908
rect 25961 5899 26019 5905
rect 25961 5896 25973 5899
rect 24544 5868 25973 5896
rect 24544 5856 24550 5868
rect 25961 5865 25973 5868
rect 26007 5865 26019 5899
rect 25961 5859 26019 5865
rect 21140 5800 21772 5828
rect 21140 5788 21146 5800
rect 22738 5788 22744 5840
rect 22796 5828 22802 5840
rect 23845 5831 23903 5837
rect 23845 5828 23857 5831
rect 22796 5800 23857 5828
rect 22796 5788 22802 5800
rect 23845 5797 23857 5800
rect 23891 5828 23903 5831
rect 28353 5831 28411 5837
rect 28353 5828 28365 5831
rect 23891 5800 24624 5828
rect 23891 5797 23903 5800
rect 23845 5791 23903 5797
rect 4908 5732 7144 5760
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 1780 5664 3249 5692
rect 1673 5655 1731 5661
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 3936 5664 4261 5692
rect 3936 5652 3942 5664
rect 4249 5661 4261 5664
rect 4295 5692 4307 5695
rect 4338 5692 4344 5704
rect 4295 5664 4344 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4908 5701 4936 5732
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 12897 5763 12955 5769
rect 7248 5732 9260 5760
rect 7248 5720 7254 5732
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6086 5692 6092 5704
rect 6043 5664 6092 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7616 5664 7849 5692
rect 7616 5652 7622 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8754 5692 8760 5704
rect 8435 5664 8760 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 9232 5692 9260 5732
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13170 5760 13176 5772
rect 12943 5732 13176 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 13538 5720 13544 5772
rect 13596 5720 13602 5772
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 14826 5760 14832 5772
rect 14608 5732 14832 5760
rect 14608 5720 14614 5732
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 16206 5760 16212 5772
rect 16040 5732 16212 5760
rect 10870 5692 10876 5704
rect 9232 5664 10876 5692
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 11112 5664 11161 5692
rect 11112 5652 11118 5664
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13280 5692 13492 5702
rect 13127 5674 14228 5692
rect 13127 5664 13308 5674
rect 13464 5664 14228 5674
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 2406 5584 2412 5636
rect 2464 5584 2470 5636
rect 3786 5584 3792 5636
rect 3844 5624 3850 5636
rect 3973 5627 4031 5633
rect 3973 5624 3985 5627
rect 3844 5596 3985 5624
rect 3844 5584 3850 5596
rect 3973 5593 3985 5596
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5624 4767 5627
rect 5258 5624 5264 5636
rect 4755 5596 5264 5624
rect 4755 5593 4767 5596
rect 4709 5587 4767 5593
rect 5258 5584 5264 5596
rect 5316 5624 5322 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 5316 5596 6653 5624
rect 5316 5584 5322 5596
rect 6641 5593 6653 5596
rect 6687 5593 6699 5627
rect 6641 5587 6699 5593
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9370 5627 9428 5633
rect 9370 5624 9382 5627
rect 8628 5596 9382 5624
rect 8628 5584 8634 5596
rect 9370 5593 9382 5596
rect 9416 5593 9428 5627
rect 9370 5587 9428 5593
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 10594 5624 10600 5636
rect 9824 5596 10600 5624
rect 9824 5584 9830 5596
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 12986 5624 12992 5636
rect 11747 5596 12992 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13170 5584 13176 5636
rect 13228 5584 13234 5636
rect 13262 5584 13268 5636
rect 13320 5584 13326 5636
rect 13403 5627 13461 5633
rect 13403 5593 13415 5627
rect 13449 5624 13461 5627
rect 14090 5624 14096 5636
rect 13449 5596 14096 5624
rect 13449 5593 13461 5596
rect 13403 5587 13461 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 3752 5528 4169 5556
rect 3752 5516 3758 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 5074 5516 5080 5568
rect 5132 5516 5138 5568
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7101 5559 7159 5565
rect 7101 5556 7113 5559
rect 7064 5528 7113 5556
rect 7064 5516 7070 5528
rect 7101 5525 7113 5528
rect 7147 5525 7159 5559
rect 7101 5519 7159 5525
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 11901 5559 11959 5565
rect 11901 5556 11913 5559
rect 9732 5528 11913 5556
rect 9732 5516 9738 5528
rect 11901 5525 11913 5528
rect 11947 5556 11959 5559
rect 13998 5556 14004 5568
rect 11947 5528 14004 5556
rect 11947 5525 11959 5528
rect 11901 5519 11959 5525
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 14200 5556 14228 5664
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 16040 5701 16068 5732
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 16531 5732 19564 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16347 5695 16405 5701
rect 16347 5661 16359 5695
rect 16393 5692 16405 5695
rect 17954 5692 17960 5704
rect 16393 5664 17960 5692
rect 16393 5661 16405 5664
rect 16347 5655 16405 5661
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5692 18659 5695
rect 18966 5692 18972 5704
rect 18647 5664 18972 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 18966 5652 18972 5664
rect 19024 5652 19030 5704
rect 19426 5652 19432 5704
rect 19484 5652 19490 5704
rect 19536 5692 19564 5732
rect 22922 5720 22928 5772
rect 22980 5760 22986 5772
rect 24596 5760 24624 5800
rect 28000 5800 28365 5828
rect 22980 5732 24348 5760
rect 24596 5732 24716 5760
rect 22980 5720 22986 5732
rect 20622 5692 20628 5704
rect 19536 5664 20628 5692
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 21729 5695 21787 5701
rect 21729 5661 21741 5695
rect 21775 5692 21787 5695
rect 22738 5692 22744 5704
rect 21775 5664 22744 5692
rect 21775 5661 21787 5664
rect 21729 5655 21787 5661
rect 22738 5652 22744 5664
rect 22796 5692 22802 5704
rect 23382 5692 23388 5704
rect 22796 5664 23388 5692
rect 22796 5652 22802 5664
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 14274 5584 14280 5636
rect 14332 5584 14338 5636
rect 16114 5584 16120 5636
rect 16172 5584 16178 5636
rect 16209 5627 16267 5633
rect 16209 5593 16221 5627
rect 16255 5624 16267 5627
rect 16574 5624 16580 5636
rect 16255 5596 16580 5624
rect 16255 5593 16267 5596
rect 16209 5587 16267 5593
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 16942 5584 16948 5636
rect 17000 5624 17006 5636
rect 17129 5627 17187 5633
rect 17129 5624 17141 5627
rect 17000 5596 17141 5624
rect 17000 5584 17006 5596
rect 17129 5593 17141 5596
rect 17175 5593 17187 5627
rect 17129 5587 17187 5593
rect 18414 5584 18420 5636
rect 18472 5584 18478 5636
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19674 5627 19732 5633
rect 19674 5624 19686 5627
rect 19392 5596 19686 5624
rect 19392 5584 19398 5596
rect 19674 5593 19686 5596
rect 19720 5593 19732 5627
rect 19674 5587 19732 5593
rect 19794 5584 19800 5636
rect 19852 5624 19858 5636
rect 21974 5627 22032 5633
rect 21974 5624 21986 5627
rect 19852 5596 21986 5624
rect 19852 5584 19858 5596
rect 21974 5593 21986 5596
rect 22020 5593 22032 5627
rect 21974 5587 22032 5593
rect 22186 5584 22192 5636
rect 22244 5624 22250 5636
rect 23569 5627 23627 5633
rect 23569 5624 23581 5627
rect 22244 5596 23581 5624
rect 22244 5584 22250 5596
rect 23569 5593 23581 5596
rect 23615 5593 23627 5627
rect 24210 5624 24216 5636
rect 23569 5587 23627 5593
rect 23952 5596 24216 5624
rect 14487 5559 14545 5565
rect 14487 5556 14499 5559
rect 14200 5528 14499 5556
rect 14487 5525 14499 5528
rect 14533 5556 14545 5559
rect 15470 5556 15476 5568
rect 14533 5528 15476 5556
rect 14533 5525 14545 5528
rect 14487 5519 14545 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16022 5556 16028 5568
rect 15887 5528 16028 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 17034 5516 17040 5568
rect 17092 5556 17098 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 17092 5528 17601 5556
rect 17092 5516 17098 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 17589 5519 17647 5525
rect 18785 5559 18843 5565
rect 18785 5525 18797 5559
rect 18831 5556 18843 5559
rect 20162 5556 20168 5568
rect 18831 5528 20168 5556
rect 18831 5525 18843 5528
rect 18785 5519 18843 5525
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 23952 5556 23980 5596
rect 24210 5584 24216 5596
rect 24268 5584 24274 5636
rect 24320 5624 24348 5732
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24688 5692 24716 5732
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 26973 5763 27031 5769
rect 26973 5760 26985 5763
rect 26476 5732 26985 5760
rect 26476 5720 26482 5732
rect 26973 5729 26985 5732
rect 27019 5729 27031 5763
rect 26973 5723 27031 5729
rect 28000 5692 28028 5800
rect 28353 5797 28365 5800
rect 28399 5797 28411 5831
rect 28353 5791 28411 5797
rect 24688 5664 28028 5692
rect 24854 5633 24860 5636
rect 24320 5596 24808 5624
rect 20588 5528 23980 5556
rect 24029 5559 24087 5565
rect 20588 5516 20594 5528
rect 24029 5525 24041 5559
rect 24075 5556 24087 5559
rect 24670 5556 24676 5568
rect 24075 5528 24676 5556
rect 24075 5525 24087 5528
rect 24029 5519 24087 5525
rect 24670 5516 24676 5528
rect 24728 5516 24734 5568
rect 24780 5556 24808 5596
rect 24848 5587 24860 5633
rect 24912 5624 24918 5636
rect 24912 5596 24948 5624
rect 24854 5584 24860 5587
rect 24912 5584 24918 5596
rect 26142 5584 26148 5636
rect 26200 5624 26206 5636
rect 27218 5627 27276 5633
rect 27218 5624 27230 5627
rect 26200 5596 27230 5624
rect 26200 5584 26206 5596
rect 27218 5593 27230 5596
rect 27264 5593 27276 5627
rect 27218 5587 27276 5593
rect 26234 5556 26240 5568
rect 24780 5528 26240 5556
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3786 5352 3792 5364
rect 3191 5324 3792 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 3881 5355 3939 5361
rect 3881 5321 3893 5355
rect 3927 5352 3939 5355
rect 3970 5352 3976 5364
rect 3927 5324 3976 5352
rect 3927 5321 3939 5324
rect 3881 5315 3939 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4798 5352 4804 5364
rect 4295 5324 4804 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5408 5324 7420 5352
rect 5408 5312 5414 5324
rect 2032 5287 2090 5293
rect 2032 5253 2044 5287
rect 2078 5284 2090 5287
rect 5442 5284 5448 5296
rect 2078 5256 5448 5284
rect 2078 5253 2090 5256
rect 2032 5247 2090 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 5902 5284 5908 5296
rect 5552 5256 5908 5284
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1728 5188 1777 5216
rect 1728 5176 1734 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4154 5216 4160 5228
rect 4111 5188 4160 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5552 5216 5580 5256
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 7392 5293 7420 5324
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 10244 5324 10916 5352
rect 7377 5287 7435 5293
rect 7377 5253 7389 5287
rect 7423 5253 7435 5287
rect 7377 5247 7435 5253
rect 8389 5287 8447 5293
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 8846 5284 8852 5296
rect 8435 5256 8852 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 9582 5244 9588 5296
rect 9640 5284 9646 5296
rect 10244 5284 10272 5324
rect 9640 5256 10272 5284
rect 10367 5287 10425 5293
rect 9640 5244 9646 5256
rect 10367 5253 10379 5287
rect 10413 5284 10425 5287
rect 10778 5284 10784 5296
rect 10413 5256 10784 5284
rect 10413 5253 10425 5256
rect 10367 5247 10425 5253
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 10888 5284 10916 5324
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 12676 5324 13277 5352
rect 12676 5312 12682 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14148 5324 14749 5352
rect 14148 5312 14154 5324
rect 12130 5287 12188 5293
rect 12130 5284 12142 5287
rect 10888 5256 12142 5284
rect 12130 5253 12142 5256
rect 12176 5253 12188 5287
rect 12130 5247 12188 5253
rect 13630 5244 13636 5296
rect 13688 5284 13694 5296
rect 14614 5287 14672 5293
rect 14614 5284 14626 5287
rect 13688 5256 14626 5284
rect 13688 5244 13694 5256
rect 14614 5253 14626 5256
rect 14660 5253 14672 5287
rect 14721 5284 14749 5324
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 14884 5324 15761 5352
rect 14884 5312 14890 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 15749 5315 15807 5321
rect 16853 5355 16911 5361
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 18693 5355 18751 5361
rect 16899 5324 18276 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 16666 5284 16672 5296
rect 14721 5256 16672 5284
rect 14614 5247 14672 5253
rect 16666 5244 16672 5256
rect 16724 5244 16730 5296
rect 17310 5244 17316 5296
rect 17368 5284 17374 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 17368 5256 17785 5284
rect 17368 5244 17374 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 17954 5244 17960 5296
rect 18012 5293 18018 5296
rect 18012 5287 18041 5293
rect 18029 5253 18041 5287
rect 18248 5284 18276 5324
rect 18693 5321 18705 5355
rect 18739 5352 18751 5355
rect 19794 5352 19800 5364
rect 18739 5324 19800 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 19981 5355 20039 5361
rect 19981 5321 19993 5355
rect 20027 5321 20039 5355
rect 19981 5315 20039 5321
rect 22005 5355 22063 5361
rect 22005 5321 22017 5355
rect 22051 5352 22063 5355
rect 22051 5324 23796 5352
rect 22051 5321 22063 5324
rect 22005 5315 22063 5321
rect 19334 5284 19340 5296
rect 18248 5256 19340 5284
rect 18012 5247 18041 5253
rect 18012 5244 18018 5247
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19996 5284 20024 5315
rect 22894 5287 22952 5293
rect 22894 5284 22906 5287
rect 19996 5256 22906 5284
rect 22894 5253 22906 5256
rect 22940 5253 22952 5287
rect 23768 5284 23796 5324
rect 24026 5312 24032 5364
rect 24084 5312 24090 5364
rect 24489 5355 24547 5361
rect 24489 5321 24501 5355
rect 24535 5352 24547 5355
rect 26786 5352 26792 5364
rect 24535 5324 26792 5352
rect 24535 5321 24547 5324
rect 24489 5315 24547 5321
rect 26786 5312 26792 5324
rect 26844 5312 26850 5364
rect 27246 5312 27252 5364
rect 27304 5312 27310 5364
rect 25470 5287 25528 5293
rect 25470 5284 25482 5287
rect 23768 5256 25482 5284
rect 22894 5247 22952 5253
rect 25470 5253 25482 5256
rect 25516 5253 25528 5287
rect 25470 5247 25528 5253
rect 6736 5228 6788 5234
rect 5031 5188 5580 5216
rect 5629 5219 5687 5225
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 6086 5216 6092 5228
rect 5675 5188 6092 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9180 5188 9720 5216
rect 9180 5176 9186 5188
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 4982 5040 4988 5092
rect 5040 5080 5046 5092
rect 5350 5080 5356 5092
rect 5040 5052 5356 5080
rect 5040 5040 5046 5052
rect 5350 5040 5356 5052
rect 5408 5080 5414 5092
rect 5460 5080 5488 5111
rect 5408 5052 5488 5080
rect 5408 5040 5414 5052
rect 5810 5040 5816 5092
rect 5868 5040 5874 5092
rect 6104 5080 6132 5176
rect 6736 5170 6788 5176
rect 6638 5080 6644 5092
rect 6104 5052 6644 5080
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 8757 5083 8815 5089
rect 8757 5049 8769 5083
rect 8803 5080 8815 5083
rect 9122 5080 9128 5092
rect 8803 5052 9128 5080
rect 8803 5049 8815 5052
rect 8757 5043 8815 5049
rect 9122 5040 9128 5052
rect 9180 5080 9186 5092
rect 9306 5080 9312 5092
rect 9180 5052 9312 5080
rect 9180 5040 9186 5052
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9692 5080 9720 5188
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 9916 5188 10057 5216
rect 9916 5176 9922 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 10134 5176 10140 5228
rect 10192 5176 10198 5228
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10284 5188 11100 5216
rect 10284 5176 10290 5188
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 9824 5120 10517 5148
rect 9824 5108 9830 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 11072 5148 11100 5188
rect 11146 5176 11152 5228
rect 11204 5176 11210 5228
rect 13354 5216 13360 5228
rect 11256 5188 13360 5216
rect 11256 5148 11284 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 15654 5216 15660 5228
rect 13955 5188 15660 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17681 5219 17739 5225
rect 17681 5185 17693 5219
rect 17727 5185 17739 5219
rect 17681 5179 17739 5185
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 11072 5120 11284 5148
rect 11885 5151 11943 5157
rect 10505 5111 10563 5117
rect 11885 5117 11897 5151
rect 11931 5117 11943 5151
rect 14182 5148 14188 5160
rect 11885 5111 11943 5117
rect 13188 5120 14188 5148
rect 11900 5080 11928 5111
rect 9692 5052 11928 5080
rect 4801 5015 4859 5021
rect 4801 4981 4813 5015
rect 4847 5012 4859 5015
rect 6454 5012 6460 5024
rect 4847 4984 6460 5012
rect 4847 4981 4859 4984
rect 4801 4975 4859 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 8846 4972 8852 5024
rect 8904 4972 8910 5024
rect 10962 4972 10968 5024
rect 11020 4972 11026 5024
rect 11900 5012 11928 5052
rect 13188 5012 13216 5120
rect 14182 5108 14188 5120
rect 14240 5148 14246 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14240 5120 14381 5148
rect 14240 5108 14246 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 17696 5148 17724 5179
rect 15528 5120 17724 5148
rect 15528 5108 15534 5120
rect 17126 5040 17132 5092
rect 17184 5080 17190 5092
rect 17880 5080 17908 5179
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 20162 5176 20168 5228
rect 20220 5176 20226 5228
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 20809 5219 20867 5225
rect 20809 5216 20821 5219
rect 20772 5188 20821 5216
rect 20772 5176 20778 5188
rect 20809 5185 20821 5188
rect 20855 5216 20867 5219
rect 21634 5216 21640 5228
rect 20855 5188 21640 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 22066 5188 22201 5216
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5148 18199 5151
rect 20438 5148 20444 5160
rect 18187 5120 20444 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 22066 5148 22094 5188
rect 22189 5185 22201 5188
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 22738 5216 22744 5228
rect 22695 5188 22744 5216
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 22738 5176 22744 5188
rect 22796 5216 22802 5228
rect 22796 5188 24348 5216
rect 22796 5176 22802 5188
rect 21315 5120 22094 5148
rect 24320 5148 24348 5188
rect 24670 5176 24676 5228
rect 24728 5176 24734 5228
rect 26234 5176 26240 5228
rect 26292 5216 26298 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26292 5188 27169 5216
rect 26292 5176 26298 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27338 5176 27344 5228
rect 27396 5176 27402 5228
rect 25130 5148 25136 5160
rect 24320 5120 25136 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 25130 5108 25136 5120
rect 25188 5148 25194 5160
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 25188 5120 25237 5148
rect 25188 5108 25194 5120
rect 25225 5117 25237 5120
rect 25271 5117 25283 5151
rect 25225 5111 25283 5117
rect 17184 5052 17908 5080
rect 17184 5040 17190 5052
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 20530 5080 20536 5092
rect 20128 5052 20536 5080
rect 20128 5040 20134 5052
rect 20530 5040 20536 5052
rect 20588 5080 20594 5092
rect 21085 5083 21143 5089
rect 21085 5080 21097 5083
rect 20588 5052 21097 5080
rect 20588 5040 20594 5052
rect 21085 5049 21097 5052
rect 21131 5049 21143 5083
rect 21085 5043 21143 5049
rect 23952 5052 24624 5080
rect 11900 4984 13216 5012
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 15654 5012 15660 5024
rect 13771 4984 15660 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 18414 5012 18420 5024
rect 16908 4984 18420 5012
rect 16908 4972 16914 4984
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19337 5015 19395 5021
rect 19337 4981 19349 5015
rect 19383 5012 19395 5015
rect 20714 5012 20720 5024
rect 19383 4984 20720 5012
rect 19383 4981 19395 4984
rect 19337 4975 19395 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 20990 4972 20996 5024
rect 21048 5012 21054 5024
rect 23952 5012 23980 5052
rect 21048 4984 23980 5012
rect 24596 5012 24624 5052
rect 26605 5015 26663 5021
rect 26605 5012 26617 5015
rect 24596 4984 26617 5012
rect 21048 4972 21054 4984
rect 26605 4981 26617 4984
rect 26651 4981 26663 5015
rect 26605 4975 26663 4981
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 382 4768 388 4820
rect 440 4808 446 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 440 4780 3157 4808
rect 440 4768 446 4780
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 3145 4771 3203 4777
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 4396 4780 4445 4808
rect 4396 4768 4402 4780
rect 4433 4777 4445 4780
rect 4479 4777 4491 4811
rect 4433 4771 4491 4777
rect 4982 4768 4988 4820
rect 5040 4768 5046 4820
rect 5629 4811 5687 4817
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 8570 4808 8576 4820
rect 5675 4780 8576 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10594 4808 10600 4820
rect 10551 4780 10600 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 11204 4780 13737 4808
rect 11204 4768 11210 4780
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 13725 4771 13783 4777
rect 17586 4768 17592 4820
rect 17644 4808 17650 4820
rect 17644 4780 19748 4808
rect 17644 4768 17650 4780
rect 5534 4740 5540 4752
rect 3620 4712 5540 4740
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1728 4644 1777 4672
rect 1728 4632 1734 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 1765 4635 1823 4641
rect 2032 4607 2090 4613
rect 2032 4573 2044 4607
rect 2078 4604 2090 4607
rect 3620 4604 3648 4712
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 8662 4740 8668 4752
rect 8435 4712 8668 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 11790 4700 11796 4752
rect 11848 4700 11854 4752
rect 13633 4743 13691 4749
rect 13633 4709 13645 4743
rect 13679 4740 13691 4743
rect 15562 4740 15568 4752
rect 13679 4712 15568 4740
rect 13679 4709 13691 4712
rect 13633 4703 13691 4709
rect 15562 4700 15568 4712
rect 15620 4740 15626 4752
rect 16390 4740 16396 4752
rect 15620 4712 16396 4740
rect 15620 4700 15626 4712
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 17218 4700 17224 4752
rect 17276 4740 17282 4752
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 17276 4712 17325 4740
rect 17276 4700 17282 4712
rect 17313 4709 17325 4712
rect 17359 4709 17371 4743
rect 17313 4703 17371 4709
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18233 4743 18291 4749
rect 18233 4740 18245 4743
rect 18104 4712 18245 4740
rect 18104 4700 18110 4712
rect 18233 4709 18245 4712
rect 18279 4709 18291 4743
rect 18233 4703 18291 4709
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 6549 4675 6607 4681
rect 3752 4644 4292 4672
rect 3752 4632 3758 4644
rect 2078 4576 3648 4604
rect 2078 4573 2090 4576
rect 2032 4567 2090 4573
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 4264 4545 4292 4644
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6595 4644 7144 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4604 5871 4607
rect 6822 4604 6828 4616
rect 5859 4576 6828 4604
rect 5859 4573 5871 4576
rect 5813 4567 5871 4573
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7116 4604 7144 4644
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11808 4672 11836 4700
rect 15378 4672 15384 4684
rect 11204 4644 11836 4672
rect 12636 4644 15384 4672
rect 11204 4632 11210 4644
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 7116 4576 9137 4604
rect 9125 4573 9137 4576
rect 9171 4604 9183 4607
rect 9171 4576 9536 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9508 4548 9536 4576
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12636 4613 12664 4644
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 17000 4644 17049 4672
rect 17000 4632 17006 4644
rect 17037 4641 17049 4644
rect 17083 4672 17095 4675
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17083 4644 17969 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 19720 4672 19748 4780
rect 20530 4768 20536 4820
rect 20588 4808 20594 4820
rect 27157 4811 27215 4817
rect 27157 4808 27169 4811
rect 20588 4780 27169 4808
rect 20588 4768 20594 4780
rect 27157 4777 27169 4780
rect 27203 4777 27215 4811
rect 27157 4771 27215 4777
rect 27706 4768 27712 4820
rect 27764 4768 27770 4820
rect 21545 4743 21603 4749
rect 21545 4709 21557 4743
rect 21591 4709 21603 4743
rect 21545 4703 21603 4709
rect 18463 4644 19656 4672
rect 19720 4644 20300 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11940 4576 12633 4604
rect 11940 4564 11946 4576
rect 12621 4573 12633 4576
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12768 4576 13277 4604
rect 12768 4564 12774 4576
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 14424 4576 14473 4604
rect 14424 4564 14430 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15289 4607 15347 4613
rect 15289 4604 15301 4607
rect 14608 4576 15301 4604
rect 14608 4564 14614 4576
rect 15289 4573 15301 4576
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4604 16083 4607
rect 18874 4604 18880 4616
rect 16071 4576 18880 4604
rect 16071 4573 16083 4576
rect 16025 4567 16083 4573
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 3936 4508 4077 4536
rect 3936 4496 3942 4508
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 4065 4499 4123 4505
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4505 4307 4539
rect 4249 4499 4307 4505
rect 6365 4539 6423 4545
rect 6365 4505 6377 4539
rect 6411 4505 6423 4539
rect 6365 4499 6423 4505
rect 4080 4468 4108 4499
rect 4338 4468 4344 4480
rect 4080 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 6380 4468 6408 4499
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7254 4539 7312 4545
rect 7254 4536 7266 4539
rect 7156 4508 7266 4536
rect 7156 4496 7162 4508
rect 7254 4505 7266 4508
rect 7300 4505 7312 4539
rect 7254 4499 7312 4505
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 9370 4539 9428 4545
rect 9370 4536 9382 4539
rect 7800 4508 9382 4536
rect 7800 4496 7806 4508
rect 9370 4505 9382 4508
rect 9416 4505 9428 4539
rect 9370 4499 9428 4505
rect 9490 4496 9496 4548
rect 9548 4496 9554 4548
rect 11517 4539 11575 4545
rect 11517 4505 11529 4539
rect 11563 4536 11575 4539
rect 11790 4536 11796 4548
rect 11563 4508 11796 4536
rect 11563 4505 11575 4508
rect 11517 4499 11575 4505
rect 11790 4496 11796 4508
rect 11848 4536 11854 4548
rect 12342 4536 12348 4548
rect 11848 4508 12348 4536
rect 11848 4496 11854 4508
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 12437 4539 12495 4545
rect 12437 4505 12449 4539
rect 12483 4536 12495 4539
rect 13722 4536 13728 4548
rect 12483 4508 13728 4536
rect 12483 4505 12495 4508
rect 12437 4499 12495 4505
rect 13722 4496 13728 4508
rect 13780 4536 13786 4548
rect 14277 4539 14335 4545
rect 14277 4536 14289 4539
rect 13780 4508 14289 4536
rect 13780 4496 13786 4508
rect 14277 4505 14289 4508
rect 14323 4505 14335 4539
rect 15470 4536 15476 4548
rect 14277 4499 14335 4505
rect 14384 4508 15476 4536
rect 8386 4468 8392 4480
rect 6380 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12158 4468 12164 4480
rect 12023 4440 12164 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12805 4471 12863 4477
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 12894 4468 12900 4480
rect 12851 4440 12900 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14384 4468 14412 4508
rect 15470 4496 15476 4508
rect 15528 4536 15534 4548
rect 16040 4536 16068 4567
rect 18874 4564 18880 4576
rect 18932 4604 18938 4616
rect 19426 4604 19432 4616
rect 18932 4576 19432 4604
rect 18932 4564 18938 4576
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19628 4613 19656 4644
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 20162 4564 20168 4616
rect 20220 4564 20226 4616
rect 20272 4604 20300 4644
rect 21560 4604 21588 4703
rect 22370 4700 22376 4752
rect 22428 4700 22434 4752
rect 21634 4632 21640 4684
rect 21692 4672 21698 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21692 4644 22017 4672
rect 21692 4632 21698 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4672 22523 4675
rect 22511 4644 24808 4672
rect 22511 4641 22523 4644
rect 22465 4635 22523 4641
rect 20272 4576 21588 4604
rect 23198 4564 23204 4616
rect 23256 4564 23262 4616
rect 23474 4564 23480 4616
rect 23532 4564 23538 4616
rect 24780 4613 24808 4644
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 25188 4644 25789 4672
rect 25188 4632 25194 4644
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 25777 4635 25835 4641
rect 27246 4632 27252 4684
rect 27304 4672 27310 4684
rect 27304 4644 27844 4672
rect 27304 4632 27310 4644
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 27614 4564 27620 4616
rect 27672 4564 27678 4616
rect 27816 4613 27844 4644
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 15528 4508 16068 4536
rect 15528 4496 15534 4508
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 20410 4539 20468 4545
rect 20410 4536 20422 4539
rect 19392 4508 20422 4536
rect 19392 4496 19398 4508
rect 20410 4505 20422 4508
rect 20456 4505 20468 4539
rect 26022 4539 26080 4545
rect 26022 4536 26034 4539
rect 20410 4499 20468 4505
rect 24596 4508 26034 4536
rect 13872 4440 14412 4468
rect 13872 4428 13878 4440
rect 14642 4428 14648 4480
rect 14700 4428 14706 4480
rect 14734 4428 14740 4480
rect 14792 4468 14798 4480
rect 15105 4471 15163 4477
rect 15105 4468 15117 4471
rect 14792 4440 15117 4468
rect 14792 4428 14798 4440
rect 15105 4437 15117 4440
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 17497 4471 17555 4477
rect 17497 4437 17509 4471
rect 17543 4468 17555 4471
rect 18230 4468 18236 4480
rect 17543 4440 18236 4468
rect 17543 4437 17555 4440
rect 17497 4431 17555 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 21266 4468 21272 4480
rect 19475 4440 21272 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 24596 4477 24624 4508
rect 26022 4505 26034 4508
rect 26068 4505 26080 4539
rect 26022 4499 26080 4505
rect 24581 4471 24639 4477
rect 24581 4437 24593 4471
rect 24627 4437 24639 4471
rect 24581 4431 24639 4437
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 10134 4264 10140 4276
rect 3896 4236 10140 4264
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 3896 4205 3924 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 15749 4267 15807 4273
rect 15749 4264 15761 4267
rect 15436 4236 15761 4264
rect 15436 4224 15442 4236
rect 15749 4233 15761 4236
rect 15795 4233 15807 4267
rect 15749 4227 15807 4233
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 21634 4264 21640 4276
rect 16172 4236 21640 4264
rect 16172 4224 16178 4236
rect 3881 4199 3939 4205
rect 3881 4196 3893 4199
rect 3568 4168 3893 4196
rect 3568 4156 3574 4168
rect 3881 4165 3893 4168
rect 3927 4165 3939 4199
rect 6270 4196 6276 4208
rect 3881 4159 3939 4165
rect 3988 4168 6276 4196
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1728 4100 1777 4128
rect 1728 4088 1734 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 2021 4131 2079 4137
rect 2021 4128 2033 4131
rect 1765 4091 1823 4097
rect 1872 4100 2033 4128
rect 1118 4020 1124 4072
rect 1176 4060 1182 4072
rect 1872 4060 1900 4100
rect 2021 4097 2033 4100
rect 2067 4097 2079 4131
rect 2021 4091 2079 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 3988 4128 4016 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 6880 4168 7236 4196
rect 6880 4156 6886 4168
rect 3743 4100 4016 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4212 4100 4537 4128
rect 4212 4088 4218 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 1176 4032 1900 4060
rect 1176 4020 1182 4032
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 5000 4060 5028 4091
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7081 4131 7139 4137
rect 7081 4128 7093 4131
rect 6512 4100 7093 4128
rect 6512 4088 6518 4100
rect 7081 4097 7093 4100
rect 7127 4097 7139 4131
rect 7208 4128 7236 4168
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 7742 4196 7748 4208
rect 7524 4168 7748 4196
rect 7524 4156 7530 4168
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 9493 4199 9551 4205
rect 9493 4165 9505 4199
rect 9539 4196 9551 4199
rect 12526 4196 12532 4208
rect 9539 4168 12532 4196
rect 9539 4165 9551 4168
rect 9493 4159 9551 4165
rect 12526 4156 12532 4168
rect 12584 4196 12590 4208
rect 13725 4199 13783 4205
rect 12584 4168 13676 4196
rect 12584 4156 12590 4168
rect 8754 4128 8760 4140
rect 7208 4100 8760 4128
rect 7081 4091 7139 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 13648 4128 13676 4168
rect 13725 4165 13737 4199
rect 13771 4196 13783 4199
rect 13814 4196 13820 4208
rect 13771 4168 13820 4196
rect 13771 4165 13783 4168
rect 13725 4159 13783 4165
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 14636 4199 14694 4205
rect 14636 4165 14648 4199
rect 14682 4196 14694 4199
rect 14734 4196 14740 4208
rect 14682 4168 14740 4196
rect 14682 4165 14694 4168
rect 14636 4159 14694 4165
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 16850 4156 16856 4208
rect 16908 4156 16914 4208
rect 17052 4205 17080 4236
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 24670 4264 24676 4276
rect 22066 4236 24676 4264
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4165 17095 4199
rect 17037 4159 17095 4165
rect 17862 4156 17868 4208
rect 17920 4196 17926 4208
rect 17920 4168 18644 4196
rect 17920 4156 17926 4168
rect 16942 4128 16948 4140
rect 9640 4100 12664 4128
rect 13648 4100 16948 4128
rect 9640 4088 9646 4100
rect 4396 4032 5028 4060
rect 6825 4063 6883 4069
rect 4396 4020 4402 4032
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 2774 3952 2780 4004
rect 2832 3992 2838 4004
rect 3145 3995 3203 4001
rect 3145 3992 3157 3995
rect 2832 3964 3157 3992
rect 2832 3952 2838 3964
rect 3145 3961 3157 3964
rect 3191 3961 3203 3995
rect 3145 3955 3203 3961
rect 4246 3952 4252 4004
rect 4304 3992 4310 4004
rect 4801 3995 4859 4001
rect 4801 3992 4813 3995
rect 4304 3964 4813 3992
rect 4304 3952 4310 3964
rect 4801 3961 4813 3964
rect 4847 3961 4859 3995
rect 4801 3955 4859 3961
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5445 3995 5503 4001
rect 5445 3992 5457 3995
rect 5224 3964 5457 3992
rect 5224 3952 5230 3964
rect 5445 3961 5457 3964
rect 5491 3961 5503 3995
rect 5445 3955 5503 3961
rect 474 3884 480 3936
rect 532 3924 538 3936
rect 2406 3924 2412 3936
rect 532 3896 2412 3924
rect 532 3884 538 3896
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 4028 3896 4077 3924
rect 4028 3884 4034 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 6730 3924 6736 3936
rect 5408 3896 6736 3924
rect 5408 3884 5414 3896
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6840 3924 6868 4023
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9272 4032 10149 4060
rect 9272 4020 9278 4032
rect 10137 4029 10149 4032
rect 10183 4060 10195 4063
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 10183 4032 12173 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 12161 4029 12173 4032
rect 12207 4060 12219 4063
rect 12342 4060 12348 4072
rect 12207 4032 12348 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 12636 4069 12664 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 18489 4131 18547 4137
rect 18489 4128 18501 4131
rect 17144 4100 18501 4128
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 13320 4032 14381 4060
rect 13320 4020 13326 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 17144 4060 17172 4100
rect 18489 4097 18501 4100
rect 18535 4097 18547 4131
rect 18616 4128 18644 4168
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 22066 4196 22094 4236
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 20772 4168 22094 4196
rect 23124 4168 23336 4196
rect 20772 4156 20778 4168
rect 21177 4132 21235 4137
rect 21100 4131 21235 4132
rect 18616 4100 19288 4128
rect 18489 4091 18547 4097
rect 15436 4032 17172 4060
rect 18233 4063 18291 4069
rect 15436 4020 15442 4032
rect 18233 4029 18245 4063
rect 18279 4029 18291 4063
rect 19260 4060 19288 4100
rect 21100 4104 21189 4131
rect 19260 4032 19656 4060
rect 18233 4023 18291 4029
rect 9950 3992 9956 4004
rect 7760 3964 9956 3992
rect 7006 3924 7012 3936
rect 6840 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7760 3924 7788 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10502 3952 10508 4004
rect 10560 3952 10566 4004
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3992 12587 3995
rect 13906 3992 13912 4004
rect 12575 3964 13912 3992
rect 12575 3961 12587 3964
rect 12529 3955 12587 3961
rect 13906 3952 13912 3964
rect 13964 3992 13970 4004
rect 14274 3992 14280 4004
rect 13964 3964 14280 3992
rect 13964 3952 13970 3964
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 18248 3992 18276 4023
rect 15580 3964 18276 3992
rect 15580 3936 15608 3964
rect 7524 3896 7788 3924
rect 7524 3884 7530 3896
rect 8202 3884 8208 3936
rect 8260 3884 8266 3936
rect 8662 3884 8668 3936
rect 8720 3884 8726 3936
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 15562 3924 15568 3936
rect 13863 3896 15568 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 17221 3927 17279 3933
rect 17221 3893 17233 3927
rect 17267 3924 17279 3927
rect 17770 3924 17776 3936
rect 17267 3896 17776 3924
rect 17267 3893 17279 3896
rect 17221 3887 17279 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18248 3924 18276 3964
rect 19518 3924 19524 3936
rect 18248 3896 19524 3924
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19628 3933 19656 4032
rect 20070 4020 20076 4072
rect 20128 4020 20134 4072
rect 20533 4063 20591 4069
rect 20533 4029 20545 4063
rect 20579 4060 20591 4063
rect 21100 4060 21128 4104
rect 21177 4097 21189 4104
rect 21223 4097 21235 4131
rect 21177 4091 21235 4097
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21600 4100 22017 4128
rect 21600 4088 21606 4100
rect 22005 4097 22017 4100
rect 22051 4128 22063 4131
rect 22186 4128 22192 4140
rect 22051 4100 22192 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22186 4088 22192 4100
rect 22244 4088 22250 4140
rect 22646 4088 22652 4140
rect 22704 4128 22710 4140
rect 23124 4128 23152 4168
rect 23198 4137 23204 4140
rect 22704 4100 23152 4128
rect 22704 4088 22710 4100
rect 23192 4091 23204 4137
rect 23198 4088 23204 4091
rect 23256 4088 23262 4140
rect 23308 4128 23336 4168
rect 23382 4156 23388 4208
rect 23440 4196 23446 4208
rect 25590 4196 25596 4208
rect 23440 4168 25596 4196
rect 23440 4156 23446 4168
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 23474 4128 23480 4140
rect 23308 4100 23480 4128
rect 23474 4088 23480 4100
rect 23532 4128 23538 4140
rect 24762 4128 24768 4140
rect 23532 4100 24768 4128
rect 23532 4088 23538 4100
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 25021 4131 25079 4137
rect 25021 4128 25033 4131
rect 24863 4100 25033 4128
rect 22830 4060 22836 4072
rect 20579 4032 21128 4060
rect 22066 4032 22836 4060
rect 20579 4029 20591 4032
rect 20533 4023 20591 4029
rect 20438 3952 20444 4004
rect 20496 3952 20502 4004
rect 20993 3995 21051 4001
rect 20993 3961 21005 3995
rect 21039 3992 21051 3995
rect 22066 3992 22094 4032
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 22925 4063 22983 4069
rect 22925 4029 22937 4063
rect 22971 4029 22983 4063
rect 22925 4023 22983 4029
rect 21039 3964 22094 3992
rect 21039 3961 21051 3964
rect 20993 3955 21051 3961
rect 22278 3952 22284 4004
rect 22336 3952 22342 4004
rect 22738 3952 22744 4004
rect 22796 3992 22802 4004
rect 22940 3992 22968 4023
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24863 4060 24891 4100
rect 25021 4097 25033 4100
rect 25067 4097 25079 4131
rect 25021 4091 25079 4097
rect 27338 4088 27344 4140
rect 27396 4088 27402 4140
rect 23992 4032 24891 4060
rect 23992 4020 23998 4032
rect 22796 3964 22968 3992
rect 22796 3952 22802 3964
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 24268 3964 24440 3992
rect 24268 3952 24274 3964
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 20588 3896 22477 3924
rect 20588 3884 20594 3896
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 22465 3887 22523 3893
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 24305 3927 24363 3933
rect 24305 3924 24317 3927
rect 22612 3896 24317 3924
rect 22612 3884 22618 3896
rect 24305 3893 24317 3896
rect 24351 3893 24363 3927
rect 24412 3924 24440 3964
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 24412 3896 26157 3924
rect 24305 3887 24363 3893
rect 26145 3893 26157 3896
rect 26191 3893 26203 3927
rect 26145 3887 26203 3893
rect 26694 3884 26700 3936
rect 26752 3924 26758 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 26752 3896 27169 3924
rect 26752 3884 26758 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27157 3887 27215 3893
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 2556 3692 3157 3720
rect 2556 3680 2562 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 4856 3692 7021 3720
rect 4856 3680 4862 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 12713 3723 12771 3729
rect 7009 3683 7067 3689
rect 8588 3692 12434 3720
rect 5718 3652 5724 3664
rect 3988 3624 5724 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1728 3556 1777 3584
rect 1728 3544 1734 3556
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2032 3519 2090 3525
rect 2032 3485 2044 3519
rect 2078 3516 2090 3519
rect 3988 3516 4016 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 6546 3612 6552 3664
rect 6604 3612 6610 3664
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 6788 3624 7236 3652
rect 6788 3612 6794 3624
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4120 3556 5580 3584
rect 4120 3544 4126 3556
rect 5552 3525 5580 3556
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 6178 3584 6184 3596
rect 5868 3556 6184 3584
rect 5868 3544 5874 3556
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 6696 3556 7052 3584
rect 6696 3544 6702 3556
rect 2078 3488 4016 3516
rect 5261 3519 5319 3525
rect 2078 3485 2090 3488
rect 2032 3479 2090 3485
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 4065 3451 4123 3457
rect 4065 3448 4077 3451
rect 3016 3420 4077 3448
rect 3016 3408 3022 3420
rect 4065 3417 4077 3420
rect 4111 3448 4123 3451
rect 4982 3448 4988 3460
rect 4111 3420 4988 3448
rect 4111 3417 4123 3420
rect 4065 3411 4123 3417
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 5074 3408 5080 3460
rect 5132 3448 5138 3460
rect 5276 3448 5304 3479
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5776 3488 6377 3516
rect 5776 3476 5782 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6914 3516 6920 3528
rect 6365 3479 6423 3485
rect 6472 3488 6920 3516
rect 6472 3448 6500 3488
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7024 3525 7052 3556
rect 7208 3525 7236 3624
rect 7282 3612 7288 3664
rect 7340 3652 7346 3664
rect 8021 3655 8079 3661
rect 8021 3652 8033 3655
rect 7340 3624 8033 3652
rect 7340 3612 7346 3624
rect 8021 3621 8033 3624
rect 8067 3621 8079 3655
rect 8021 3615 8079 3621
rect 8588 3584 8616 3692
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 12066 3652 12072 3664
rect 11839 3624 12072 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 12406 3652 12434 3692
rect 12713 3689 12725 3723
rect 12759 3720 12771 3723
rect 16482 3720 16488 3732
rect 12759 3692 16488 3720
rect 12759 3689 12771 3692
rect 12713 3683 12771 3689
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 16942 3680 16948 3732
rect 17000 3680 17006 3732
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 19334 3720 19340 3732
rect 18371 3692 19340 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 20162 3720 20168 3732
rect 19576 3692 20168 3720
rect 19576 3680 19582 3692
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 24029 3723 24087 3729
rect 24029 3720 24041 3723
rect 22066 3692 24041 3720
rect 12802 3652 12808 3664
rect 12406 3624 12808 3652
rect 12802 3612 12808 3624
rect 12860 3652 12866 3664
rect 13078 3652 13084 3664
rect 12860 3624 13084 3652
rect 12860 3612 12866 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 17678 3612 17684 3664
rect 17736 3652 17742 3664
rect 17862 3652 17868 3664
rect 17736 3624 17868 3652
rect 17736 3612 17742 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 19794 3612 19800 3664
rect 19852 3612 19858 3664
rect 20622 3612 20628 3664
rect 20680 3612 20686 3664
rect 20806 3612 20812 3664
rect 20864 3652 20870 3664
rect 21545 3655 21603 3661
rect 21545 3652 21557 3655
rect 20864 3624 21557 3652
rect 20864 3612 20870 3624
rect 21545 3621 21557 3624
rect 21591 3652 21603 3655
rect 22066 3652 22094 3692
rect 24029 3689 24041 3692
rect 24075 3689 24087 3723
rect 24029 3683 24087 3689
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 25096 3692 27016 3720
rect 25096 3680 25102 3692
rect 21591 3624 22094 3652
rect 21591 3621 21603 3624
rect 21545 3615 21603 3621
rect 7852 3556 8616 3584
rect 7852 3525 7880 3556
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8720 3556 10548 3584
rect 8720 3544 8726 3556
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7837 3519 7895 3525
rect 7193 3479 7251 3485
rect 7300 3488 7788 3516
rect 5132 3420 6500 3448
rect 5132 3408 5138 3420
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 7300 3448 7328 3488
rect 7653 3451 7711 3457
rect 7653 3448 7665 3451
rect 6696 3420 7328 3448
rect 7392 3420 7665 3448
rect 6696 3408 6702 3420
rect 4154 3340 4160 3392
rect 4212 3340 4218 3392
rect 5442 3340 5448 3392
rect 5500 3340 5506 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 7392 3380 7420 3420
rect 7653 3417 7665 3420
rect 7699 3417 7711 3451
rect 7760 3448 7788 3488
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 9088 3488 9229 3516
rect 9088 3476 9094 3488
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 10134 3516 10140 3528
rect 9548 3488 10140 3516
rect 9548 3476 9554 3488
rect 10134 3476 10140 3488
rect 10192 3516 10198 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10192 3488 10425 3516
rect 10192 3476 10198 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10520 3516 10548 3556
rect 15562 3544 15568 3596
rect 15620 3544 15626 3596
rect 20640 3584 20668 3612
rect 22554 3584 22560 3596
rect 20640 3556 22560 3584
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 24394 3544 24400 3596
rect 24452 3584 24458 3596
rect 24762 3584 24768 3596
rect 24452 3556 24768 3584
rect 24452 3544 24458 3556
rect 24762 3544 24768 3556
rect 24820 3584 24826 3596
rect 26988 3593 27016 3692
rect 28350 3680 28356 3732
rect 28408 3680 28414 3732
rect 25133 3587 25191 3593
rect 25133 3584 25145 3587
rect 24820 3556 25145 3584
rect 24820 3544 24826 3556
rect 25133 3553 25145 3556
rect 25179 3553 25191 3587
rect 25133 3547 25191 3553
rect 26973 3587 27031 3593
rect 26973 3553 26985 3587
rect 27019 3553 27031 3587
rect 26973 3547 27031 3553
rect 10669 3519 10727 3525
rect 10669 3516 10681 3519
rect 10520 3488 10681 3516
rect 10413 3479 10471 3485
rect 10669 3485 10681 3488
rect 10715 3485 10727 3519
rect 10669 3479 10727 3485
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13538 3516 13544 3528
rect 13228 3488 13544 3516
rect 13228 3476 13234 3488
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13780 3488 14289 3516
rect 13780 3476 13786 3488
rect 14277 3485 14289 3488
rect 14323 3516 14335 3519
rect 15470 3516 15476 3528
rect 14323 3488 15476 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15821 3519 15879 3525
rect 15821 3516 15833 3519
rect 15712 3488 15833 3516
rect 15712 3476 15718 3488
rect 15821 3485 15833 3488
rect 15867 3485 15879 3519
rect 15821 3479 15879 3485
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18288 3488 18521 3516
rect 18288 3476 18294 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 22646 3476 22652 3528
rect 22704 3476 22710 3528
rect 27062 3476 27068 3528
rect 27120 3516 27126 3528
rect 27229 3519 27287 3525
rect 27229 3516 27241 3519
rect 27120 3488 27241 3516
rect 27120 3476 27126 3488
rect 27229 3485 27241 3488
rect 27275 3485 27287 3519
rect 27229 3479 27287 3485
rect 7760 3420 8156 3448
rect 7653 3411 7711 3417
rect 6328 3352 7420 3380
rect 8128 3380 8156 3420
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 9401 3451 9459 3457
rect 9401 3448 9413 3451
rect 9364 3420 9413 3448
rect 9364 3408 9370 3420
rect 9401 3417 9413 3420
rect 9447 3448 9459 3451
rect 10318 3448 10324 3460
rect 9447 3420 10324 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10318 3408 10324 3420
rect 10376 3448 10382 3460
rect 13357 3451 13415 3457
rect 13357 3448 13369 3451
rect 10376 3420 13369 3448
rect 10376 3408 10382 3420
rect 13357 3417 13369 3420
rect 13403 3448 13415 3451
rect 13740 3448 13768 3476
rect 13403 3420 13768 3448
rect 14461 3451 14519 3457
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 14461 3417 14473 3451
rect 14507 3448 14519 3451
rect 14507 3420 15884 3448
rect 14507 3417 14519 3420
rect 14461 3411 14519 3417
rect 10410 3380 10416 3392
rect 8128 3352 10416 3380
rect 6328 3340 6334 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 13722 3340 13728 3392
rect 13780 3340 13786 3392
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15286 3380 15292 3392
rect 14691 3352 15292 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15856 3380 15884 3420
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 17405 3451 17463 3457
rect 17405 3448 17417 3451
rect 15988 3420 17417 3448
rect 15988 3408 15994 3420
rect 17405 3417 17417 3420
rect 17451 3417 17463 3451
rect 17405 3411 17463 3417
rect 19429 3451 19487 3457
rect 19429 3417 19441 3451
rect 19475 3448 19487 3451
rect 20070 3448 20076 3460
rect 19475 3420 20076 3448
rect 19475 3417 19487 3420
rect 19429 3411 19487 3417
rect 20070 3408 20076 3420
rect 20128 3448 20134 3460
rect 20349 3451 20407 3457
rect 20349 3448 20361 3451
rect 20128 3420 20361 3448
rect 20128 3408 20134 3420
rect 20349 3417 20361 3420
rect 20395 3448 20407 3451
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 20395 3420 21281 3448
rect 20395 3417 20407 3420
rect 20349 3411 20407 3417
rect 21269 3417 21281 3420
rect 21315 3448 21327 3451
rect 21542 3448 21548 3460
rect 21315 3420 21548 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 21542 3408 21548 3420
rect 21600 3408 21606 3460
rect 21910 3408 21916 3460
rect 21968 3448 21974 3460
rect 22894 3451 22952 3457
rect 22894 3448 22906 3451
rect 21968 3420 22906 3448
rect 21968 3408 21974 3420
rect 22894 3417 22906 3420
rect 22940 3417 22952 3451
rect 22894 3411 22952 3417
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 24854 3448 24860 3460
rect 23072 3420 24860 3448
rect 23072 3408 23078 3420
rect 24854 3408 24860 3420
rect 24912 3408 24918 3460
rect 25038 3408 25044 3460
rect 25096 3448 25102 3460
rect 25378 3451 25436 3457
rect 25378 3448 25390 3451
rect 25096 3420 25390 3448
rect 25096 3408 25102 3420
rect 25378 3417 25390 3420
rect 25424 3417 25436 3451
rect 25378 3411 25436 3417
rect 16758 3380 16764 3392
rect 15856 3352 16764 3380
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17092 3352 17877 3380
rect 17092 3340 17098 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19668 3352 19901 3380
rect 19668 3340 19674 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 19889 3343 19947 3349
rect 20809 3383 20867 3389
rect 20809 3349 20821 3383
rect 20855 3380 20867 3383
rect 21358 3380 21364 3392
rect 20855 3352 21364 3380
rect 20855 3349 20867 3352
rect 20809 3343 20867 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 21729 3383 21787 3389
rect 21729 3380 21741 3383
rect 21508 3352 21741 3380
rect 21508 3340 21514 3352
rect 21729 3349 21741 3352
rect 21775 3349 21787 3383
rect 21729 3343 21787 3349
rect 22278 3340 22284 3392
rect 22336 3380 22342 3392
rect 24026 3380 24032 3392
rect 22336 3352 24032 3380
rect 22336 3340 22342 3352
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 26510 3340 26516 3392
rect 26568 3340 26574 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 3602 3176 3608 3188
rect 1811 3148 3608 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 7561 3179 7619 3185
rect 4387 3148 6960 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 2130 3108 2136 3120
rect 1780 3080 2136 3108
rect 1578 3000 1584 3052
rect 1636 3000 1642 3052
rect 1780 3049 1808 3080
rect 2130 3068 2136 3080
rect 2188 3068 2194 3120
rect 4154 3108 4160 3120
rect 2976 3080 4160 3108
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2976 3049 3004 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 6546 3108 6552 3120
rect 5552 3080 6552 3108
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1912 3012 2237 3040
rect 1912 3000 1918 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 3228 3043 3286 3049
rect 3228 3009 3240 3043
rect 3274 3040 3286 3043
rect 4062 3040 4068 3052
rect 3274 3012 4068 3040
rect 3274 3009 3286 3012
rect 3228 3003 3286 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 5350 3040 5356 3052
rect 4847 3012 5356 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5552 3049 5580 3080
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 6932 3108 6960 3148
rect 7561 3145 7573 3179
rect 7607 3176 7619 3179
rect 11977 3179 12035 3185
rect 7607 3148 11928 3176
rect 7607 3145 7619 3148
rect 7561 3139 7619 3145
rect 7466 3108 7472 3120
rect 6932 3080 7472 3108
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5074 2932 5080 2984
rect 5132 2932 5138 2984
rect 6546 2932 6552 2984
rect 6604 2932 6610 2984
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 2958 2904 2964 2916
rect 2455 2876 2964 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 3896 2876 5365 2904
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3896 2836 3924 2876
rect 5353 2873 5365 2876
rect 5399 2873 5411 2907
rect 5353 2867 5411 2873
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 6932 2904 6960 3080
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 9582 3108 9588 3120
rect 7760 3080 9588 3108
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 7760 3049 7788 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 11900 3108 11928 3148
rect 11977 3145 11989 3179
rect 12023 3176 12035 3179
rect 12023 3148 12434 3176
rect 12023 3145 12035 3148
rect 11977 3139 12035 3145
rect 12406 3108 12434 3148
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 13630 3176 13636 3188
rect 12768 3148 13636 3176
rect 12768 3136 12774 3148
rect 13630 3136 13636 3148
rect 13688 3176 13694 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13688 3148 14013 3176
rect 13688 3136 13694 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 14001 3139 14059 3145
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 14424 3148 15853 3176
rect 14424 3136 14430 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 20254 3176 20260 3188
rect 17460 3148 20260 3176
rect 17460 3136 17466 3148
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 20349 3179 20407 3185
rect 20349 3145 20361 3179
rect 20395 3176 20407 3179
rect 20438 3176 20444 3188
rect 20395 3148 20444 3176
rect 20395 3145 20407 3148
rect 20349 3139 20407 3145
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 26510 3176 26516 3188
rect 21784 3148 26516 3176
rect 21784 3136 21790 3148
rect 26510 3136 26516 3148
rect 26568 3136 26574 3188
rect 14706 3111 14764 3117
rect 14706 3108 14718 3111
rect 9732 3080 11100 3108
rect 11900 3080 12296 3108
rect 12406 3080 14718 3108
rect 9732 3068 9738 3080
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8472 3043 8530 3049
rect 8472 3009 8484 3043
rect 8518 3040 8530 3043
rect 10413 3043 10471 3049
rect 8518 3012 9812 3040
rect 8518 3009 8530 3012
rect 8472 3003 8530 3009
rect 7024 2972 7052 3000
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7024 2944 8217 2972
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 9784 2972 9812 3012
rect 10413 3009 10425 3043
rect 10459 3040 10471 3043
rect 10594 3040 10600 3052
rect 10459 3012 10600 3040
rect 10459 3009 10471 3012
rect 10413 3003 10471 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11072 3049 11100 3080
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 12158 3000 12164 3052
rect 12216 3000 12222 3052
rect 12268 3040 12296 3080
rect 14706 3077 14718 3080
rect 14752 3077 14764 3111
rect 14706 3071 14764 3077
rect 15470 3068 15476 3120
rect 15528 3108 15534 3120
rect 15654 3108 15660 3120
rect 15528 3080 15660 3108
rect 15528 3068 15534 3080
rect 15654 3068 15660 3080
rect 15712 3108 15718 3120
rect 16850 3108 16856 3120
rect 15712 3080 16856 3108
rect 15712 3068 15718 3080
rect 16850 3068 16856 3080
rect 16908 3108 16914 3120
rect 17129 3111 17187 3117
rect 17129 3108 17141 3111
rect 16908 3080 17141 3108
rect 16908 3068 16914 3080
rect 17129 3077 17141 3080
rect 17175 3077 17187 3111
rect 17129 3071 17187 3077
rect 17310 3068 17316 3120
rect 17368 3068 17374 3120
rect 17497 3111 17555 3117
rect 17497 3077 17509 3111
rect 17543 3108 17555 3111
rect 20898 3108 20904 3120
rect 17543 3080 20904 3108
rect 17543 3077 17555 3080
rect 17497 3071 17555 3077
rect 20898 3068 20904 3080
rect 20956 3068 20962 3120
rect 20993 3111 21051 3117
rect 20993 3077 21005 3111
rect 21039 3108 21051 3111
rect 21542 3108 21548 3120
rect 21039 3080 21548 3108
rect 21039 3077 21051 3080
rect 20993 3071 21051 3077
rect 21542 3068 21548 3080
rect 21600 3068 21606 3120
rect 24118 3068 24124 3120
rect 24176 3108 24182 3120
rect 24176 3080 26464 3108
rect 24176 3068 24182 3080
rect 12877 3043 12935 3049
rect 12877 3040 12889 3043
rect 12268 3012 12889 3040
rect 12877 3009 12889 3012
rect 12923 3009 12935 3043
rect 12877 3003 12935 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 13320 3012 14473 3040
rect 13320 3000 13326 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 18489 3043 18547 3049
rect 18489 3040 18501 3043
rect 14461 3003 14519 3009
rect 17236 3012 18501 3040
rect 11238 2972 11244 2984
rect 9784 2944 11244 2972
rect 8205 2935 8263 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 12618 2932 12624 2984
rect 12676 2932 12682 2984
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 17236 2972 17264 3012
rect 18489 3009 18501 3012
rect 18535 3009 18547 3043
rect 18489 3003 18547 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 26436 3049 26464 3080
rect 22261 3043 22319 3049
rect 22261 3040 22273 3043
rect 21968 3012 22273 3040
rect 21968 3000 21974 3012
rect 22261 3009 22273 3012
rect 22307 3009 22319 3043
rect 24653 3043 24711 3049
rect 24653 3040 24665 3043
rect 22261 3003 22319 3009
rect 23492 3012 24665 3040
rect 15528 2944 17264 2972
rect 15528 2932 15534 2944
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 17644 2944 18245 2972
rect 17644 2932 17650 2944
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 22002 2932 22008 2984
rect 22060 2932 22066 2984
rect 6871 2876 6960 2904
rect 7009 2907 7067 2913
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7009 2873 7021 2907
rect 7055 2904 7067 2907
rect 9585 2907 9643 2913
rect 7055 2876 8248 2904
rect 7055 2873 7067 2876
rect 7009 2867 7067 2873
rect 2832 2808 3924 2836
rect 2832 2796 2838 2808
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 6730 2836 6736 2848
rect 5040 2808 6736 2836
rect 5040 2796 5046 2808
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 8220 2836 8248 2876
rect 9585 2873 9597 2907
rect 9631 2904 9643 2907
rect 9766 2904 9772 2916
rect 9631 2876 9772 2904
rect 9631 2873 9643 2876
rect 9585 2867 9643 2873
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 10229 2907 10287 2913
rect 10229 2873 10241 2907
rect 10275 2904 10287 2907
rect 12526 2904 12532 2916
rect 10275 2876 12532 2904
rect 10275 2873 10287 2876
rect 10229 2867 10287 2873
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 17954 2904 17960 2916
rect 15396 2876 17960 2904
rect 9490 2836 9496 2848
rect 8220 2808 9496 2836
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10870 2796 10876 2848
rect 10928 2796 10934 2848
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 15396 2836 15424 2876
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 21361 2907 21419 2913
rect 21361 2904 21373 2907
rect 20312 2876 21373 2904
rect 20312 2864 20318 2876
rect 21361 2873 21373 2876
rect 21407 2904 21419 2907
rect 21726 2904 21732 2916
rect 21407 2876 21732 2904
rect 21407 2873 21419 2876
rect 21361 2867 21419 2873
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 23382 2864 23388 2916
rect 23440 2864 23446 2916
rect 13596 2808 15424 2836
rect 13596 2796 13602 2808
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 19613 2839 19671 2845
rect 19613 2836 19625 2839
rect 15896 2808 19625 2836
rect 15896 2796 15902 2808
rect 19613 2805 19625 2808
rect 19659 2805 19671 2839
rect 19613 2799 19671 2805
rect 21453 2839 21511 2845
rect 21453 2805 21465 2839
rect 21499 2836 21511 2839
rect 22278 2836 22284 2848
rect 21499 2808 22284 2836
rect 21499 2805 21511 2808
rect 21453 2799 21511 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 23492 2836 23520 3012
rect 24653 3009 24665 3012
rect 24699 3009 24711 3043
rect 24653 3003 24711 3009
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 24394 2932 24400 2984
rect 24452 2932 24458 2984
rect 25774 2864 25780 2916
rect 25832 2864 25838 2916
rect 26234 2864 26240 2916
rect 26292 2864 26298 2916
rect 22704 2808 23520 2836
rect 22704 2796 22710 2808
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 2958 2592 2964 2644
rect 3016 2592 3022 2644
rect 6546 2632 6552 2644
rect 4356 2604 6552 2632
rect 4356 2505 4384 2604
rect 6546 2592 6552 2604
rect 6604 2632 6610 2644
rect 6604 2604 6914 2632
rect 6604 2592 6610 2604
rect 4706 2524 4712 2576
rect 4764 2524 4770 2576
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 6886 2496 6914 2604
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 7432 2604 8493 2632
rect 7432 2592 7438 2604
rect 8481 2601 8493 2604
rect 8527 2632 8539 2635
rect 9950 2632 9956 2644
rect 8527 2604 9956 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10560 2604 10977 2632
rect 10560 2592 10566 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11296 2604 12664 2632
rect 11296 2592 11302 2604
rect 12636 2576 12664 2604
rect 12802 2592 12808 2644
rect 12860 2592 12866 2644
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 15378 2632 15384 2644
rect 14323 2604 15384 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16448 2604 17141 2632
rect 16448 2592 16454 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17678 2632 17684 2644
rect 17460 2604 17684 2632
rect 17460 2592 17466 2604
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18233 2635 18291 2641
rect 18233 2601 18245 2635
rect 18279 2632 18291 2635
rect 21174 2632 21180 2644
rect 18279 2604 21180 2632
rect 18279 2601 18291 2604
rect 18233 2595 18291 2601
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 22204 2604 24041 2632
rect 12618 2524 12624 2576
rect 12676 2564 12682 2576
rect 13262 2564 13268 2576
rect 12676 2536 13268 2564
rect 12676 2524 12682 2536
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 13541 2567 13599 2573
rect 13541 2533 13553 2567
rect 13587 2564 13599 2567
rect 15470 2564 15476 2576
rect 13587 2536 15476 2564
rect 13587 2533 13599 2536
rect 13541 2527 13599 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 17494 2524 17500 2576
rect 17552 2564 17558 2576
rect 18690 2564 18696 2576
rect 17552 2536 18696 2564
rect 17552 2524 17558 2536
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 19426 2524 19432 2576
rect 19484 2524 19490 2576
rect 21634 2524 21640 2576
rect 21692 2564 21698 2576
rect 22204 2564 22232 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 25682 2592 25688 2644
rect 25740 2632 25746 2644
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 25740 2604 25973 2632
rect 25740 2592 25746 2604
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 25961 2595 26019 2601
rect 21692 2536 22232 2564
rect 21692 2524 21698 2536
rect 6886 2468 7236 2496
rect 4341 2459 4399 2465
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 1837 2431 1895 2437
rect 1837 2428 1849 2431
rect 1728 2400 1849 2428
rect 1728 2388 1734 2400
rect 1837 2397 1849 2400
rect 1883 2397 1895 2431
rect 1837 2391 1895 2397
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 7006 2428 7012 2440
rect 5316 2400 7012 2428
rect 5316 2388 5322 2400
rect 7006 2388 7012 2400
rect 7064 2428 7070 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 7064 2400 7113 2428
rect 7064 2388 7070 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7208 2428 7236 2468
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11020 2468 11560 2496
rect 11020 2456 11026 2468
rect 7368 2431 7426 2437
rect 7208 2400 7328 2428
rect 7101 2391 7159 2397
rect 5528 2363 5586 2369
rect 5528 2329 5540 2363
rect 5574 2360 5586 2363
rect 7190 2360 7196 2372
rect 5574 2332 7196 2360
rect 5574 2329 5586 2332
rect 5528 2323 5586 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 7300 2360 7328 2400
rect 7368 2397 7380 2431
rect 7414 2428 7426 2431
rect 8202 2428 8208 2440
rect 7414 2400 8208 2428
rect 7414 2397 7426 2400
rect 7368 2391 7426 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9674 2428 9680 2440
rect 9631 2400 9680 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 10134 2428 10140 2440
rect 9732 2400 10140 2428
rect 9732 2388 9738 2400
rect 10134 2388 10140 2400
rect 10192 2428 10198 2440
rect 11238 2428 11244 2440
rect 10192 2400 11244 2428
rect 10192 2388 10198 2400
rect 11238 2388 11244 2400
rect 11296 2428 11302 2440
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 11296 2400 11437 2428
rect 11296 2388 11302 2400
rect 11425 2397 11437 2400
rect 11471 2397 11483 2431
rect 11532 2428 11560 2468
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15252 2468 15516 2496
rect 15252 2456 15258 2468
rect 15488 2440 15516 2468
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 20438 2496 20444 2508
rect 17920 2468 20444 2496
rect 17920 2456 17926 2468
rect 20438 2456 20444 2468
rect 20496 2456 20502 2508
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22554 2496 22560 2508
rect 22152 2468 22560 2496
rect 22152 2456 22158 2468
rect 22554 2456 22560 2468
rect 22612 2496 22618 2508
rect 22649 2499 22707 2505
rect 22649 2496 22661 2499
rect 22612 2468 22661 2496
rect 22612 2456 22618 2468
rect 22649 2465 22661 2468
rect 22695 2465 22707 2499
rect 22649 2459 22707 2465
rect 11681 2431 11739 2437
rect 11681 2428 11693 2431
rect 11532 2400 11693 2428
rect 11425 2391 11483 2397
rect 11681 2397 11693 2400
rect 11727 2397 11739 2431
rect 11681 2391 11739 2397
rect 13722 2388 13728 2440
rect 13780 2388 13786 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14642 2428 14648 2440
rect 14507 2400 14648 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15620 2400 15761 2428
rect 15620 2388 15626 2400
rect 15749 2397 15761 2400
rect 15795 2428 15807 2431
rect 17402 2428 17408 2440
rect 15795 2400 17408 2428
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18196 2400 18429 2428
rect 18196 2388 18202 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 18874 2428 18880 2440
rect 18656 2400 18880 2428
rect 18656 2388 18662 2400
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 20162 2428 20168 2440
rect 19760 2400 20168 2428
rect 19760 2388 19766 2400
rect 20162 2388 20168 2400
rect 20220 2428 20226 2440
rect 20530 2428 20536 2440
rect 20220 2400 20536 2428
rect 20220 2388 20226 2400
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 23382 2428 23388 2440
rect 21692 2400 23388 2428
rect 21692 2388 21698 2400
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 24394 2388 24400 2440
rect 24452 2428 24458 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24452 2400 24593 2428
rect 24452 2388 24458 2400
rect 24581 2397 24593 2400
rect 24627 2428 24639 2431
rect 26697 2431 26755 2437
rect 26697 2428 26709 2431
rect 24627 2400 26709 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 26697 2397 26709 2400
rect 26743 2397 26755 2431
rect 26697 2391 26755 2397
rect 26786 2388 26792 2440
rect 26844 2428 26850 2440
rect 26953 2431 27011 2437
rect 26953 2428 26965 2431
rect 26844 2400 26965 2428
rect 26844 2388 26850 2400
rect 26953 2397 26965 2400
rect 26999 2397 27011 2431
rect 26953 2391 27011 2397
rect 9214 2360 9220 2372
rect 7300 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9852 2363 9910 2369
rect 9852 2329 9864 2363
rect 9898 2360 9910 2363
rect 9898 2332 11744 2360
rect 9898 2329 9910 2332
rect 9852 2323 9910 2329
rect 11716 2304 11744 2332
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 15994 2363 16052 2369
rect 15994 2360 16006 2363
rect 15252 2332 16006 2360
rect 15252 2320 15258 2332
rect 15994 2329 16006 2332
rect 16040 2329 16052 2363
rect 20789 2363 20847 2369
rect 20789 2360 20801 2363
rect 15994 2323 16052 2329
rect 17604 2332 20801 2360
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 6641 2295 6699 2301
rect 6641 2261 6653 2295
rect 6687 2292 6699 2295
rect 8386 2292 8392 2304
rect 6687 2264 8392 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 15105 2295 15163 2301
rect 15105 2261 15117 2295
rect 15151 2292 15163 2295
rect 17494 2292 17500 2304
rect 15151 2264 17500 2292
rect 15151 2261 15163 2264
rect 15105 2255 15163 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 17604 2301 17632 2332
rect 20789 2329 20801 2332
rect 20835 2329 20847 2363
rect 20789 2323 20847 2329
rect 21266 2320 21272 2372
rect 21324 2360 21330 2372
rect 22894 2363 22952 2369
rect 22894 2360 22906 2363
rect 21324 2332 22906 2360
rect 21324 2320 21330 2332
rect 22894 2329 22906 2332
rect 22940 2329 22952 2363
rect 22894 2323 22952 2329
rect 24848 2363 24906 2369
rect 24848 2329 24860 2363
rect 24894 2360 24906 2363
rect 24946 2360 24952 2372
rect 24894 2332 24952 2360
rect 24894 2329 24906 2332
rect 24848 2323 24906 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 17589 2295 17647 2301
rect 17589 2261 17601 2295
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 20438 2252 20444 2304
rect 20496 2292 20502 2304
rect 21913 2295 21971 2301
rect 21913 2292 21925 2295
rect 20496 2264 21925 2292
rect 20496 2252 20502 2264
rect 21913 2261 21925 2264
rect 21959 2261 21971 2295
rect 21913 2255 21971 2261
rect 22370 2252 22376 2304
rect 22428 2292 22434 2304
rect 28077 2295 28135 2301
rect 28077 2292 28089 2295
rect 22428 2264 28089 2292
rect 22428 2252 22434 2264
rect 28077 2261 28089 2264
rect 28123 2261 28135 2295
rect 28077 2255 28135 2261
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 3510 2048 3516 2100
rect 3568 2048 3574 2100
rect 4154 2048 4160 2100
rect 4212 2048 4218 2100
rect 5813 2091 5871 2097
rect 5813 2057 5825 2091
rect 5859 2088 5871 2091
rect 7098 2088 7104 2100
rect 5859 2060 7104 2088
rect 5859 2057 5871 2060
rect 5813 2051 5871 2057
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 9122 2048 9128 2100
rect 9180 2088 9186 2100
rect 9309 2091 9367 2097
rect 9309 2088 9321 2091
rect 9180 2060 9321 2088
rect 9180 2048 9186 2060
rect 9309 2057 9321 2060
rect 9355 2057 9367 2091
rect 9309 2051 9367 2057
rect 11146 2048 11152 2100
rect 11204 2048 11210 2100
rect 11808 2060 25912 2088
rect 2400 2023 2458 2029
rect 2400 1989 2412 2023
rect 2446 2020 2458 2023
rect 2590 2020 2596 2032
rect 2446 1992 2596 2020
rect 2446 1989 2458 1992
rect 2400 1983 2458 1989
rect 2590 1980 2596 1992
rect 2648 1980 2654 2032
rect 2133 1955 2191 1961
rect 2133 1921 2145 1955
rect 2179 1952 2191 1955
rect 3973 1955 4031 1961
rect 3973 1952 3985 1955
rect 2179 1924 3985 1952
rect 2179 1921 2191 1924
rect 2133 1915 2191 1921
rect 3973 1921 3985 1924
rect 4019 1952 4031 1955
rect 4172 1952 4200 2048
rect 4240 2023 4298 2029
rect 4240 1989 4252 2023
rect 4286 2020 4298 2023
rect 6638 2020 6644 2032
rect 4286 1992 6644 2020
rect 4286 1989 4298 1992
rect 4240 1983 4298 1989
rect 6638 1980 6644 1992
rect 6696 1980 6702 2032
rect 7650 1980 7656 2032
rect 7708 2020 7714 2032
rect 8174 2023 8232 2029
rect 8174 2020 8186 2023
rect 7708 1992 8186 2020
rect 7708 1980 7714 1992
rect 8174 1989 8186 1992
rect 8220 1989 8232 2023
rect 8174 1983 8232 1989
rect 9490 1980 9496 2032
rect 9548 2020 9554 2032
rect 11808 2020 11836 2060
rect 9548 1992 11836 2020
rect 9548 1980 9554 1992
rect 12342 1980 12348 2032
rect 12400 2020 12406 2032
rect 12400 1992 12480 2020
rect 12400 1980 12406 1992
rect 5258 1952 5264 1964
rect 4019 1924 5264 1952
rect 4019 1921 4031 1924
rect 3973 1915 4031 1921
rect 5258 1912 5264 1924
rect 5316 1912 5322 1964
rect 5994 1912 6000 1964
rect 6052 1912 6058 1964
rect 6546 1912 6552 1964
rect 6604 1952 6610 1964
rect 7009 1955 7067 1961
rect 7009 1952 7021 1955
rect 6604 1924 7021 1952
rect 6604 1912 6610 1924
rect 7009 1921 7021 1924
rect 7055 1921 7067 1955
rect 7009 1915 7067 1921
rect 7098 1912 7104 1964
rect 7156 1952 7162 1964
rect 7929 1955 7987 1961
rect 7929 1952 7941 1955
rect 7156 1924 7941 1952
rect 7156 1912 7162 1924
rect 7929 1921 7941 1924
rect 7975 1921 7987 1955
rect 8938 1952 8944 1964
rect 7929 1915 7987 1921
rect 8036 1924 8944 1952
rect 8036 1884 8064 1924
rect 8938 1912 8944 1924
rect 8996 1912 9002 1964
rect 9674 1912 9680 1964
rect 9732 1952 9738 1964
rect 9769 1955 9827 1961
rect 9769 1952 9781 1955
rect 9732 1924 9781 1952
rect 9732 1912 9738 1924
rect 9769 1921 9781 1924
rect 9815 1921 9827 1955
rect 9769 1915 9827 1921
rect 10036 1955 10094 1961
rect 10036 1921 10048 1955
rect 10082 1952 10094 1955
rect 10962 1952 10968 1964
rect 10082 1924 10968 1952
rect 10082 1921 10094 1924
rect 10036 1915 10094 1921
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 11885 1955 11943 1961
rect 11885 1921 11897 1955
rect 11931 1921 11943 1955
rect 12452 1952 12480 1992
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 13510 2023 13568 2029
rect 13510 2020 13522 2023
rect 12584 1992 13522 2020
rect 12584 1980 12590 1992
rect 13510 1989 13522 1992
rect 13556 1989 13568 2023
rect 13510 1983 13568 1989
rect 14458 1980 14464 2032
rect 14516 2020 14522 2032
rect 15197 2023 15255 2029
rect 15197 2020 15209 2023
rect 14516 1992 15209 2020
rect 14516 1980 14522 1992
rect 15197 1989 15209 1992
rect 15243 2020 15255 2023
rect 15930 2020 15936 2032
rect 15243 1992 15936 2020
rect 15243 1989 15255 1992
rect 15197 1983 15255 1989
rect 15930 1980 15936 1992
rect 15988 1980 15994 2032
rect 16482 1980 16488 2032
rect 16540 2020 16546 2032
rect 17098 2023 17156 2029
rect 17098 2020 17110 2023
rect 16540 1992 17110 2020
rect 16540 1980 16546 1992
rect 17098 1989 17110 1992
rect 17144 1989 17156 2023
rect 17098 1983 17156 1989
rect 17494 1980 17500 2032
rect 17552 2020 17558 2032
rect 18938 2023 18996 2029
rect 18938 2020 18950 2023
rect 17552 1992 18950 2020
rect 17552 1980 17558 1992
rect 18938 1989 18950 1992
rect 18984 1989 18996 2023
rect 22250 2023 22308 2029
rect 22250 2020 22262 2023
rect 18938 1983 18996 1989
rect 20548 1992 22262 2020
rect 12452 1924 13124 1952
rect 11885 1915 11943 1921
rect 6886 1856 8064 1884
rect 11900 1884 11928 1915
rect 12805 1887 12863 1893
rect 12805 1884 12817 1887
rect 11900 1856 12817 1884
rect 4706 1708 4712 1760
rect 4764 1748 4770 1760
rect 5353 1751 5411 1757
rect 5353 1748 5365 1751
rect 4764 1720 5365 1748
rect 4764 1708 4770 1720
rect 5353 1717 5365 1720
rect 5399 1748 5411 1751
rect 6886 1748 6914 1856
rect 12805 1853 12817 1856
rect 12851 1853 12863 1887
rect 13096 1884 13124 1924
rect 13262 1912 13268 1964
rect 13320 1912 13326 1964
rect 14476 1952 14504 1980
rect 13372 1924 14504 1952
rect 16301 1955 16359 1961
rect 13372 1884 13400 1924
rect 16301 1921 16313 1955
rect 16347 1921 16359 1955
rect 16301 1915 16359 1921
rect 16853 1955 16911 1961
rect 16853 1921 16865 1955
rect 16899 1952 16911 1955
rect 17402 1952 17408 1964
rect 16899 1924 17408 1952
rect 16899 1921 16911 1924
rect 16853 1915 16911 1921
rect 13096 1856 13400 1884
rect 15657 1887 15715 1893
rect 12805 1847 12863 1853
rect 15657 1853 15669 1887
rect 15703 1884 15715 1887
rect 16316 1884 16344 1915
rect 17402 1912 17408 1924
rect 17460 1912 17466 1964
rect 17678 1912 17684 1964
rect 17736 1952 17742 1964
rect 17736 1924 17908 1952
rect 17736 1912 17742 1924
rect 15703 1856 16344 1884
rect 17880 1884 17908 1924
rect 18598 1912 18604 1964
rect 18656 1952 18662 1964
rect 18693 1955 18751 1961
rect 18693 1952 18705 1955
rect 18656 1924 18705 1952
rect 18656 1912 18662 1924
rect 18693 1921 18705 1924
rect 18739 1921 18751 1955
rect 18693 1915 18751 1921
rect 18800 1924 20208 1952
rect 18800 1884 18828 1924
rect 17880 1856 18828 1884
rect 15703 1853 15715 1856
rect 15657 1847 15715 1853
rect 7374 1776 7380 1828
rect 7432 1776 7438 1828
rect 12250 1816 12256 1828
rect 10704 1788 12256 1816
rect 5399 1720 6914 1748
rect 7469 1751 7527 1757
rect 5399 1717 5411 1720
rect 5353 1711 5411 1717
rect 7469 1717 7481 1751
rect 7515 1748 7527 1751
rect 10704 1748 10732 1788
rect 12250 1776 12256 1788
rect 12308 1776 12314 1828
rect 12710 1776 12716 1828
rect 12768 1776 12774 1828
rect 14274 1776 14280 1828
rect 14332 1816 14338 1828
rect 14645 1819 14703 1825
rect 14645 1816 14657 1819
rect 14332 1788 14657 1816
rect 14332 1776 14338 1788
rect 14645 1785 14657 1788
rect 14691 1785 14703 1819
rect 14645 1779 14703 1785
rect 15562 1776 15568 1828
rect 15620 1776 15626 1828
rect 17862 1776 17868 1828
rect 17920 1816 17926 1828
rect 17920 1788 18368 1816
rect 17920 1776 17926 1788
rect 7515 1720 10732 1748
rect 11701 1751 11759 1757
rect 7515 1717 7527 1720
rect 7469 1711 7527 1717
rect 11701 1717 11713 1751
rect 11747 1748 11759 1751
rect 15102 1748 15108 1760
rect 11747 1720 15108 1748
rect 11747 1717 11759 1720
rect 11701 1711 11759 1717
rect 15102 1708 15108 1720
rect 15160 1708 15166 1760
rect 16117 1751 16175 1757
rect 16117 1717 16129 1751
rect 16163 1748 16175 1751
rect 17218 1748 17224 1760
rect 16163 1720 17224 1748
rect 16163 1717 16175 1720
rect 16117 1711 16175 1717
rect 17218 1708 17224 1720
rect 17276 1708 17282 1760
rect 17954 1708 17960 1760
rect 18012 1748 18018 1760
rect 18233 1751 18291 1757
rect 18233 1748 18245 1751
rect 18012 1720 18245 1748
rect 18012 1708 18018 1720
rect 18233 1717 18245 1720
rect 18279 1717 18291 1751
rect 18340 1748 18368 1788
rect 20073 1751 20131 1757
rect 20073 1748 20085 1751
rect 18340 1720 20085 1748
rect 18233 1711 18291 1717
rect 20073 1717 20085 1720
rect 20119 1717 20131 1751
rect 20180 1748 20208 1924
rect 20548 1825 20576 1992
rect 22250 1989 22262 1992
rect 22296 1989 22308 2023
rect 22250 1983 22308 1989
rect 22554 1980 22560 2032
rect 22612 2020 22618 2032
rect 23842 2020 23848 2032
rect 22612 1992 23848 2020
rect 22612 1980 22618 1992
rect 23842 1980 23848 1992
rect 23900 1980 23906 2032
rect 20717 1955 20775 1961
rect 20717 1921 20729 1955
rect 20763 1952 20775 1955
rect 20898 1952 20904 1964
rect 20763 1924 20904 1952
rect 20763 1921 20775 1924
rect 20717 1915 20775 1921
rect 20898 1912 20904 1924
rect 20956 1912 20962 1964
rect 21358 1912 21364 1964
rect 21416 1912 21422 1964
rect 21542 1912 21548 1964
rect 21600 1952 21606 1964
rect 25884 1961 25912 2060
rect 26326 2048 26332 2100
rect 26384 2048 26390 2100
rect 24101 1955 24159 1961
rect 24101 1952 24113 1955
rect 21600 1924 24113 1952
rect 21600 1912 21606 1924
rect 24101 1921 24113 1924
rect 24147 1921 24159 1955
rect 24101 1915 24159 1921
rect 25869 1955 25927 1961
rect 25869 1921 25881 1955
rect 25915 1921 25927 1955
rect 25869 1915 25927 1921
rect 26510 1912 26516 1964
rect 26568 1912 26574 1964
rect 20622 1844 20628 1896
rect 20680 1884 20686 1896
rect 22005 1887 22063 1893
rect 22005 1884 22017 1887
rect 20680 1856 22017 1884
rect 20680 1844 20686 1856
rect 22005 1853 22017 1856
rect 22051 1853 22063 1887
rect 22005 1847 22063 1853
rect 23842 1844 23848 1896
rect 23900 1844 23906 1896
rect 20533 1819 20591 1825
rect 20533 1785 20545 1819
rect 20579 1785 20591 1819
rect 21634 1816 21640 1828
rect 20533 1779 20591 1785
rect 20640 1788 21640 1816
rect 20640 1748 20668 1788
rect 21634 1776 21640 1788
rect 21692 1776 21698 1828
rect 23382 1776 23388 1828
rect 23440 1776 23446 1828
rect 25682 1776 25688 1828
rect 25740 1776 25746 1828
rect 20180 1720 20668 1748
rect 21177 1751 21235 1757
rect 20073 1711 20131 1717
rect 21177 1717 21189 1751
rect 21223 1748 21235 1751
rect 22646 1748 22652 1760
rect 21223 1720 22652 1748
rect 21223 1717 21235 1720
rect 21177 1711 21235 1717
rect 22646 1708 22652 1720
rect 22704 1708 22710 1760
rect 23474 1708 23480 1760
rect 23532 1748 23538 1760
rect 25225 1751 25283 1757
rect 25225 1748 25237 1751
rect 23532 1720 25237 1748
rect 23532 1708 23538 1720
rect 25225 1717 25237 1720
rect 25271 1717 25283 1751
rect 25225 1711 25283 1717
rect 1104 1658 28888 1680
rect 1104 1606 4423 1658
rect 4475 1606 4487 1658
rect 4539 1606 4551 1658
rect 4603 1606 4615 1658
rect 4667 1606 4679 1658
rect 4731 1606 11369 1658
rect 11421 1606 11433 1658
rect 11485 1606 11497 1658
rect 11549 1606 11561 1658
rect 11613 1606 11625 1658
rect 11677 1606 18315 1658
rect 18367 1606 18379 1658
rect 18431 1606 18443 1658
rect 18495 1606 18507 1658
rect 18559 1606 18571 1658
rect 18623 1606 25261 1658
rect 25313 1606 25325 1658
rect 25377 1606 25389 1658
rect 25441 1606 25453 1658
rect 25505 1606 25517 1658
rect 25569 1606 28888 1658
rect 1104 1584 28888 1606
rect 5537 1547 5595 1553
rect 5537 1513 5549 1547
rect 5583 1544 5595 1547
rect 6362 1544 6368 1556
rect 5583 1516 6368 1544
rect 5583 1513 5595 1516
rect 5537 1507 5595 1513
rect 6362 1504 6368 1516
rect 6420 1504 6426 1556
rect 18138 1544 18144 1556
rect 17512 1516 18144 1544
rect 9766 1436 9772 1488
rect 9824 1436 9830 1488
rect 14550 1436 14556 1488
rect 14608 1476 14614 1488
rect 14829 1479 14887 1485
rect 14829 1476 14841 1479
rect 14608 1448 14841 1476
rect 14608 1436 14614 1448
rect 14829 1445 14841 1448
rect 14875 1476 14887 1479
rect 17310 1476 17316 1488
rect 14875 1448 17316 1476
rect 14875 1445 14887 1448
rect 14829 1439 14887 1445
rect 17310 1436 17316 1448
rect 17368 1436 17374 1488
rect 1578 1368 1584 1420
rect 1636 1368 1642 1420
rect 4154 1368 4160 1420
rect 4212 1368 4218 1420
rect 10520 1380 11192 1408
rect 1848 1343 1906 1349
rect 1848 1309 1860 1343
rect 1894 1340 1906 1343
rect 2774 1340 2780 1352
rect 1894 1312 2780 1340
rect 1894 1309 1906 1312
rect 1848 1303 1906 1309
rect 2774 1300 2780 1312
rect 2832 1300 2838 1352
rect 6641 1343 6699 1349
rect 6641 1309 6653 1343
rect 6687 1340 6699 1343
rect 6730 1340 6736 1352
rect 6687 1312 6736 1340
rect 6687 1309 6699 1312
rect 6641 1303 6699 1309
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 10318 1300 10324 1352
rect 10376 1340 10382 1352
rect 10413 1343 10471 1349
rect 10413 1340 10425 1343
rect 10376 1312 10425 1340
rect 10376 1300 10382 1312
rect 10413 1309 10425 1312
rect 10459 1309 10471 1343
rect 10413 1303 10471 1309
rect 4424 1275 4482 1281
rect 4424 1241 4436 1275
rect 4470 1272 4482 1275
rect 6908 1275 6966 1281
rect 4470 1244 5948 1272
rect 4470 1241 4482 1244
rect 4424 1235 4482 1241
rect 5920 1216 5948 1244
rect 6908 1241 6920 1275
rect 6954 1272 6966 1275
rect 8202 1272 8208 1284
rect 6954 1244 8208 1272
rect 6954 1241 6966 1244
rect 6908 1235 6966 1241
rect 8202 1232 8208 1244
rect 8260 1232 8266 1284
rect 9493 1275 9551 1281
rect 9493 1241 9505 1275
rect 9539 1272 9551 1275
rect 10520 1272 10548 1380
rect 10597 1343 10655 1349
rect 10597 1309 10609 1343
rect 10643 1340 10655 1343
rect 10686 1340 10692 1352
rect 10643 1312 10692 1340
rect 10643 1309 10655 1312
rect 10597 1303 10655 1309
rect 10686 1300 10692 1312
rect 10744 1300 10750 1352
rect 10781 1343 10839 1349
rect 10781 1309 10793 1343
rect 10827 1340 10839 1343
rect 11054 1340 11060 1352
rect 10827 1312 11060 1340
rect 10827 1309 10839 1312
rect 10781 1303 10839 1309
rect 11054 1300 11060 1312
rect 11112 1300 11118 1352
rect 11164 1340 11192 1380
rect 11238 1368 11244 1420
rect 11296 1408 11302 1420
rect 11701 1411 11759 1417
rect 11701 1408 11713 1411
rect 11296 1380 11713 1408
rect 11296 1368 11302 1380
rect 11701 1377 11713 1380
rect 11747 1377 11759 1411
rect 11701 1371 11759 1377
rect 13648 1380 13860 1408
rect 11790 1340 11796 1352
rect 11164 1312 11796 1340
rect 11790 1300 11796 1312
rect 11848 1300 11854 1352
rect 9539 1244 10548 1272
rect 9539 1241 9551 1244
rect 9493 1235 9551 1241
rect 2961 1207 3019 1213
rect 2961 1173 2973 1207
rect 3007 1204 3019 1207
rect 5810 1204 5816 1216
rect 3007 1176 5816 1204
rect 3007 1173 3019 1176
rect 2961 1167 3019 1173
rect 5810 1164 5816 1176
rect 5868 1164 5874 1216
rect 5902 1164 5908 1216
rect 5960 1164 5966 1216
rect 7742 1164 7748 1216
rect 7800 1204 7806 1216
rect 8021 1207 8079 1213
rect 8021 1204 8033 1207
rect 7800 1176 8033 1204
rect 7800 1164 7806 1176
rect 8021 1173 8033 1176
rect 8067 1173 8079 1207
rect 8021 1167 8079 1173
rect 9950 1164 9956 1216
rect 10008 1164 10014 1216
rect 10704 1204 10732 1300
rect 10870 1232 10876 1284
rect 10928 1272 10934 1284
rect 11946 1275 12004 1281
rect 11946 1272 11958 1275
rect 10928 1244 11958 1272
rect 10928 1232 10934 1244
rect 11946 1241 11958 1244
rect 11992 1241 12004 1275
rect 11946 1235 12004 1241
rect 13081 1207 13139 1213
rect 13081 1204 13093 1207
rect 10704 1176 13093 1204
rect 13081 1173 13093 1176
rect 13127 1173 13139 1207
rect 13081 1167 13139 1173
rect 13541 1207 13599 1213
rect 13541 1173 13553 1207
rect 13587 1204 13599 1207
rect 13648 1204 13676 1380
rect 13725 1343 13783 1349
rect 13725 1309 13737 1343
rect 13771 1309 13783 1343
rect 13832 1340 13860 1380
rect 14458 1368 14464 1420
rect 14516 1368 14522 1420
rect 15654 1408 15660 1420
rect 15488 1380 15660 1408
rect 15194 1340 15200 1352
rect 13832 1312 15200 1340
rect 13725 1303 13783 1309
rect 13587 1176 13676 1204
rect 13740 1204 13768 1303
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
rect 15381 1275 15439 1281
rect 15381 1241 15393 1275
rect 15427 1272 15439 1275
rect 15488 1272 15516 1380
rect 15654 1368 15660 1380
rect 15712 1368 15718 1420
rect 15749 1411 15807 1417
rect 15749 1377 15761 1411
rect 15795 1408 15807 1411
rect 17512 1408 17540 1516
rect 18138 1504 18144 1516
rect 18196 1504 18202 1556
rect 18690 1504 18696 1556
rect 18748 1544 18754 1556
rect 23474 1544 23480 1556
rect 18748 1516 23480 1544
rect 18748 1504 18754 1516
rect 23474 1504 23480 1516
rect 23532 1504 23538 1556
rect 15795 1380 15976 1408
rect 15795 1377 15807 1380
rect 15749 1371 15807 1377
rect 15565 1343 15623 1349
rect 15565 1309 15577 1343
rect 15611 1340 15623 1343
rect 15838 1340 15844 1352
rect 15611 1312 15844 1340
rect 15611 1309 15623 1312
rect 15565 1303 15623 1309
rect 15838 1300 15844 1312
rect 15896 1300 15902 1352
rect 15948 1340 15976 1380
rect 16960 1380 17540 1408
rect 19352 1380 19564 1408
rect 16960 1340 16988 1380
rect 15948 1312 16988 1340
rect 17034 1300 17040 1352
rect 17092 1300 17098 1352
rect 17402 1300 17408 1352
rect 17460 1340 17466 1352
rect 17497 1343 17555 1349
rect 17497 1340 17509 1343
rect 17460 1312 17509 1340
rect 17460 1300 17466 1312
rect 17497 1309 17509 1312
rect 17543 1309 17555 1343
rect 17497 1303 17555 1309
rect 17586 1300 17592 1352
rect 17644 1340 17650 1352
rect 19352 1340 19380 1380
rect 17644 1312 19380 1340
rect 17644 1300 17650 1312
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 19536 1340 19564 1380
rect 23842 1368 23848 1420
rect 23900 1408 23906 1420
rect 24581 1411 24639 1417
rect 24581 1408 24593 1411
rect 23900 1380 24593 1408
rect 23900 1368 23906 1380
rect 24581 1377 24593 1380
rect 24627 1377 24639 1411
rect 24581 1371 24639 1377
rect 19536 1312 19840 1340
rect 17742 1275 17800 1281
rect 17742 1272 17754 1275
rect 15427 1244 15516 1272
rect 15672 1244 17754 1272
rect 15427 1241 15439 1244
rect 15381 1235 15439 1241
rect 14921 1207 14979 1213
rect 14921 1204 14933 1207
rect 13740 1176 14933 1204
rect 13587 1173 13599 1176
rect 13541 1167 13599 1173
rect 14921 1173 14933 1176
rect 14967 1173 14979 1207
rect 14921 1167 14979 1173
rect 15102 1164 15108 1216
rect 15160 1204 15166 1216
rect 15672 1204 15700 1244
rect 17742 1241 17754 1244
rect 17788 1241 17800 1275
rect 19674 1275 19732 1281
rect 19674 1272 19686 1275
rect 17742 1235 17800 1241
rect 18248 1244 19686 1272
rect 15160 1176 15700 1204
rect 16853 1207 16911 1213
rect 15160 1164 15166 1176
rect 16853 1173 16865 1207
rect 16899 1204 16911 1207
rect 18248 1204 18276 1244
rect 19674 1241 19686 1244
rect 19720 1241 19732 1275
rect 19812 1272 19840 1312
rect 21450 1300 21456 1352
rect 21508 1300 21514 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22554 1340 22560 1352
rect 22051 1312 22560 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22554 1300 22560 1312
rect 22612 1300 22618 1352
rect 23124 1312 23980 1340
rect 22250 1275 22308 1281
rect 22250 1272 22262 1275
rect 19812 1244 22262 1272
rect 19674 1235 19732 1241
rect 22250 1241 22262 1244
rect 22296 1241 22308 1275
rect 22250 1235 22308 1241
rect 16899 1176 18276 1204
rect 16899 1173 16911 1176
rect 16853 1167 16911 1173
rect 18874 1164 18880 1216
rect 18932 1164 18938 1216
rect 20806 1164 20812 1216
rect 20864 1164 20870 1216
rect 21269 1207 21327 1213
rect 21269 1173 21281 1207
rect 21315 1204 21327 1207
rect 23124 1204 23152 1312
rect 23198 1232 23204 1284
rect 23256 1272 23262 1284
rect 23256 1244 23888 1272
rect 23256 1232 23262 1244
rect 21315 1176 23152 1204
rect 21315 1173 21327 1176
rect 21269 1167 21327 1173
rect 23382 1164 23388 1216
rect 23440 1164 23446 1216
rect 23860 1213 23888 1244
rect 23845 1207 23903 1213
rect 23845 1173 23857 1207
rect 23891 1173 23903 1207
rect 23952 1204 23980 1312
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 24854 1349 24860 1352
rect 24848 1340 24860 1349
rect 24815 1312 24860 1340
rect 24848 1303 24860 1312
rect 24854 1300 24860 1303
rect 24912 1300 24918 1352
rect 26602 1300 26608 1352
rect 26660 1300 26666 1352
rect 27338 1300 27344 1352
rect 27396 1340 27402 1352
rect 27617 1343 27675 1349
rect 27617 1340 27629 1343
rect 27396 1312 27629 1340
rect 27396 1300 27402 1312
rect 27617 1309 27629 1312
rect 27663 1309 27675 1343
rect 27617 1303 27675 1309
rect 25038 1204 25044 1216
rect 23952 1176 25044 1204
rect 23845 1167 23903 1173
rect 25038 1164 25044 1176
rect 25096 1164 25102 1216
rect 25590 1164 25596 1216
rect 25648 1204 25654 1216
rect 25961 1207 26019 1213
rect 25961 1204 25973 1207
rect 25648 1176 25973 1204
rect 25648 1164 25654 1176
rect 25961 1173 25973 1176
rect 26007 1173 26019 1207
rect 25961 1167 26019 1173
rect 26418 1164 26424 1216
rect 26476 1164 26482 1216
rect 27154 1164 27160 1216
rect 27212 1164 27218 1216
rect 1104 1114 29048 1136
rect 1104 1062 7896 1114
rect 7948 1062 7960 1114
rect 8012 1062 8024 1114
rect 8076 1062 8088 1114
rect 8140 1062 8152 1114
rect 8204 1062 14842 1114
rect 14894 1062 14906 1114
rect 14958 1062 14970 1114
rect 15022 1062 15034 1114
rect 15086 1062 15098 1114
rect 15150 1062 21788 1114
rect 21840 1062 21852 1114
rect 21904 1062 21916 1114
rect 21968 1062 21980 1114
rect 22032 1062 22044 1114
rect 22096 1062 28734 1114
rect 28786 1062 28798 1114
rect 28850 1062 28862 1114
rect 28914 1062 28926 1114
rect 28978 1062 28990 1114
rect 29042 1062 29048 1114
rect 1104 1040 29048 1062
rect 10962 960 10968 1012
rect 11020 1000 11026 1012
rect 26418 1000 26424 1012
rect 11020 972 26424 1000
rect 11020 960 11026 972
rect 26418 960 26424 972
rect 26476 960 26482 1012
rect 9950 892 9956 944
rect 10008 932 10014 944
rect 26602 932 26608 944
rect 10008 904 26608 932
rect 10008 892 10014 904
rect 26602 892 26608 904
rect 26660 892 26666 944
rect 4062 824 4068 876
rect 4120 864 4126 876
rect 27154 864 27160 876
rect 4120 836 27160 864
rect 4120 824 4126 836
rect 27154 824 27160 836
rect 27212 824 27218 876
rect 5902 756 5908 808
rect 5960 796 5966 808
rect 26694 796 26700 808
rect 5960 768 26700 796
rect 5960 756 5966 768
rect 26694 756 26700 768
rect 26752 756 26758 808
rect 16758 688 16764 740
rect 16816 728 16822 740
rect 20806 728 20812 740
rect 16816 700 20812 728
rect 16816 688 16822 700
rect 20806 688 20812 700
rect 20864 688 20870 740
rect 23382 728 23388 740
rect 21008 700 23388 728
rect 3970 620 3976 672
rect 4028 660 4034 672
rect 4028 632 12434 660
rect 4028 620 4034 632
rect 12406 524 12434 632
rect 15562 552 15568 604
rect 15620 592 15626 604
rect 18874 592 18880 604
rect 15620 564 18880 592
rect 15620 552 15626 564
rect 18874 552 18880 564
rect 18932 552 18938 604
rect 19058 552 19064 604
rect 19116 592 19122 604
rect 21008 592 21036 700
rect 23382 688 23388 700
rect 23440 688 23446 740
rect 27338 660 27344 672
rect 19116 564 21036 592
rect 22066 632 27344 660
rect 19116 552 19122 564
rect 22066 524 22094 632
rect 27338 620 27344 632
rect 27396 620 27402 672
rect 12406 496 22094 524
<< via1 >>
rect 14004 33600 14056 33652
rect 21180 33600 21232 33652
rect 12808 33532 12860 33584
rect 19156 33532 19208 33584
rect 9220 33464 9272 33516
rect 16764 33464 16816 33516
rect 17132 33464 17184 33516
rect 25596 33464 25648 33516
rect 14464 33396 14516 33448
rect 24952 33396 25004 33448
rect 7656 33328 7708 33380
rect 16488 33328 16540 33380
rect 16856 33328 16908 33380
rect 23388 33328 23440 33380
rect 4804 33260 4856 33312
rect 6920 33260 6972 33312
rect 27344 33260 27396 33312
rect 10048 33192 10100 33244
rect 10416 33124 10468 33176
rect 17132 33124 17184 33176
rect 17316 33192 17368 33244
rect 27896 33192 27948 33244
rect 26792 33124 26844 33176
rect 8484 33056 8536 33108
rect 13820 33056 13872 33108
rect 14096 33056 14148 33108
rect 19064 33056 19116 33108
rect 19156 33056 19208 33108
rect 23480 33056 23532 33108
rect 13728 32988 13780 33040
rect 23664 32988 23716 33040
rect 12532 32920 12584 32972
rect 16396 32920 16448 32972
rect 16764 32920 16816 32972
rect 27712 32920 27764 32972
rect 2320 32852 2372 32904
rect 9496 32852 9548 32904
rect 13176 32852 13228 32904
rect 16948 32852 17000 32904
rect 17132 32852 17184 32904
rect 8300 32784 8352 32836
rect 17316 32784 17368 32836
rect 19248 32852 19300 32904
rect 22928 32852 22980 32904
rect 21272 32784 21324 32836
rect 11704 32716 11756 32768
rect 14648 32716 14700 32768
rect 16488 32716 16540 32768
rect 26424 32784 26476 32836
rect 22192 32716 22244 32768
rect 25780 32716 25832 32768
rect 7896 32614 7948 32666
rect 7960 32614 8012 32666
rect 8024 32614 8076 32666
rect 8088 32614 8140 32666
rect 8152 32614 8204 32666
rect 14842 32614 14894 32666
rect 14906 32614 14958 32666
rect 14970 32614 15022 32666
rect 15034 32614 15086 32666
rect 15098 32614 15150 32666
rect 21788 32614 21840 32666
rect 21852 32614 21904 32666
rect 21916 32614 21968 32666
rect 21980 32614 22032 32666
rect 22044 32614 22096 32666
rect 28734 32614 28786 32666
rect 28798 32614 28850 32666
rect 28862 32614 28914 32666
rect 28926 32614 28978 32666
rect 28990 32614 29042 32666
rect 2320 32555 2372 32564
rect 2320 32521 2329 32555
rect 2329 32521 2363 32555
rect 2363 32521 2372 32555
rect 2320 32512 2372 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 3332 32444 3384 32496
rect 8392 32444 8444 32496
rect 2872 32376 2924 32428
rect 2412 32351 2464 32360
rect 2412 32317 2421 32351
rect 2421 32317 2455 32351
rect 2455 32317 2464 32351
rect 2412 32308 2464 32317
rect 2688 32308 2740 32360
rect 7012 32376 7064 32428
rect 9956 32512 10008 32564
rect 9588 32444 9640 32496
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 3240 32308 3292 32360
rect 4804 32351 4856 32360
rect 4804 32317 4813 32351
rect 4813 32317 4847 32351
rect 4847 32317 4856 32351
rect 4804 32308 4856 32317
rect 6644 32308 6696 32360
rect 7472 32308 7524 32360
rect 2872 32215 2924 32224
rect 2872 32181 2881 32215
rect 2881 32181 2915 32215
rect 2915 32181 2924 32215
rect 2872 32172 2924 32181
rect 3148 32172 3200 32224
rect 4252 32240 4304 32292
rect 5172 32283 5224 32292
rect 5172 32249 5181 32283
rect 5181 32249 5215 32283
rect 5215 32249 5224 32283
rect 5172 32240 5224 32249
rect 7196 32240 7248 32292
rect 7748 32240 7800 32292
rect 11152 32376 11204 32428
rect 9036 32308 9088 32360
rect 11612 32444 11664 32496
rect 14372 32512 14424 32564
rect 22100 32512 22152 32564
rect 13268 32351 13320 32360
rect 13268 32317 13277 32351
rect 13277 32317 13311 32351
rect 13311 32317 13320 32351
rect 13268 32308 13320 32317
rect 13636 32376 13688 32428
rect 14372 32376 14424 32428
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 14648 32376 14700 32428
rect 16028 32376 16080 32428
rect 17316 32376 17368 32428
rect 18052 32376 18104 32428
rect 20444 32444 20496 32496
rect 14188 32308 14240 32360
rect 14556 32308 14608 32360
rect 16672 32308 16724 32360
rect 19432 32308 19484 32360
rect 10140 32240 10192 32292
rect 12440 32240 12492 32292
rect 12532 32240 12584 32292
rect 11612 32172 11664 32224
rect 12808 32215 12860 32224
rect 12808 32181 12817 32215
rect 12817 32181 12851 32215
rect 12851 32181 12860 32215
rect 12808 32172 12860 32181
rect 13544 32283 13596 32292
rect 13544 32249 13553 32283
rect 13553 32249 13587 32283
rect 13587 32249 13596 32283
rect 13544 32240 13596 32249
rect 14832 32240 14884 32292
rect 16212 32240 16264 32292
rect 13728 32215 13780 32224
rect 13728 32181 13737 32215
rect 13737 32181 13771 32215
rect 13771 32181 13780 32215
rect 13728 32172 13780 32181
rect 13912 32172 13964 32224
rect 17408 32240 17460 32292
rect 22100 32376 22152 32428
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 25872 32512 25924 32564
rect 25136 32444 25188 32496
rect 23480 32419 23532 32428
rect 23480 32385 23489 32419
rect 23489 32385 23523 32419
rect 23523 32385 23532 32419
rect 23480 32376 23532 32385
rect 25964 32376 26016 32428
rect 23572 32308 23624 32360
rect 19616 32172 19668 32224
rect 20444 32172 20496 32224
rect 21180 32215 21232 32224
rect 21180 32181 21189 32215
rect 21189 32181 21223 32215
rect 21223 32181 21232 32215
rect 21180 32172 21232 32181
rect 21272 32172 21324 32224
rect 28080 32240 28132 32292
rect 27988 32215 28040 32224
rect 27988 32181 27997 32215
rect 27997 32181 28031 32215
rect 28031 32181 28040 32215
rect 27988 32172 28040 32181
rect 4423 32070 4475 32122
rect 4487 32070 4539 32122
rect 4551 32070 4603 32122
rect 4615 32070 4667 32122
rect 4679 32070 4731 32122
rect 11369 32070 11421 32122
rect 11433 32070 11485 32122
rect 11497 32070 11549 32122
rect 11561 32070 11613 32122
rect 11625 32070 11677 32122
rect 18315 32070 18367 32122
rect 18379 32070 18431 32122
rect 18443 32070 18495 32122
rect 18507 32070 18559 32122
rect 18571 32070 18623 32122
rect 25261 32070 25313 32122
rect 25325 32070 25377 32122
rect 25389 32070 25441 32122
rect 25453 32070 25505 32122
rect 25517 32070 25569 32122
rect 3332 32011 3384 32020
rect 3332 31977 3341 32011
rect 3341 31977 3375 32011
rect 3375 31977 3384 32011
rect 3332 31968 3384 31977
rect 3424 31968 3476 32020
rect 27988 31968 28040 32020
rect 4252 31900 4304 31952
rect 4344 31900 4396 31952
rect 5264 31943 5316 31952
rect 5264 31909 5273 31943
rect 5273 31909 5307 31943
rect 5307 31909 5316 31943
rect 5264 31900 5316 31909
rect 7748 31943 7800 31952
rect 7748 31909 7757 31943
rect 7757 31909 7791 31943
rect 7791 31909 7800 31943
rect 7748 31900 7800 31909
rect 8300 31900 8352 31952
rect 8484 31943 8536 31952
rect 8484 31909 8493 31943
rect 8493 31909 8527 31943
rect 8527 31909 8536 31943
rect 8484 31900 8536 31909
rect 10600 31900 10652 31952
rect 13176 31900 13228 31952
rect 2596 31875 2648 31884
rect 2596 31841 2605 31875
rect 2605 31841 2639 31875
rect 2639 31841 2648 31875
rect 2596 31832 2648 31841
rect 2688 31875 2740 31884
rect 2688 31841 2697 31875
rect 2697 31841 2731 31875
rect 2731 31841 2740 31875
rect 2688 31832 2740 31841
rect 2872 31832 2924 31884
rect 10508 31832 10560 31884
rect 3976 31764 4028 31816
rect 3056 31696 3108 31748
rect 4160 31764 4212 31816
rect 5724 31807 5776 31816
rect 5724 31773 5733 31807
rect 5733 31773 5767 31807
rect 5767 31773 5776 31807
rect 5724 31764 5776 31773
rect 6092 31807 6144 31816
rect 6092 31773 6101 31807
rect 6101 31773 6135 31807
rect 6135 31773 6144 31807
rect 6092 31764 6144 31773
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 7564 31764 7616 31816
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 10048 31764 10100 31816
rect 10416 31807 10468 31816
rect 10416 31773 10425 31807
rect 10425 31773 10459 31807
rect 10459 31773 10468 31807
rect 10416 31764 10468 31773
rect 9588 31739 9640 31748
rect 9588 31705 9597 31739
rect 9597 31705 9631 31739
rect 9631 31705 9640 31739
rect 9588 31696 9640 31705
rect 4344 31628 4396 31680
rect 4528 31628 4580 31680
rect 5172 31628 5224 31680
rect 10692 31807 10744 31816
rect 10692 31773 10701 31807
rect 10701 31773 10735 31807
rect 10735 31773 10744 31807
rect 10692 31764 10744 31773
rect 13452 31764 13504 31816
rect 13268 31739 13320 31748
rect 13268 31705 13277 31739
rect 13277 31705 13311 31739
rect 13311 31705 13320 31739
rect 13268 31696 13320 31705
rect 17592 31900 17644 31952
rect 18236 31900 18288 31952
rect 20812 31943 20864 31952
rect 20812 31909 20821 31943
rect 20821 31909 20855 31943
rect 20855 31909 20864 31943
rect 20812 31900 20864 31909
rect 22928 31943 22980 31952
rect 22928 31909 22937 31943
rect 22937 31909 22971 31943
rect 22971 31909 22980 31943
rect 22928 31900 22980 31909
rect 14096 31832 14148 31884
rect 15752 31764 15804 31816
rect 14188 31696 14240 31748
rect 16304 31696 16356 31748
rect 17132 31764 17184 31816
rect 16580 31696 16632 31748
rect 16856 31696 16908 31748
rect 17684 31696 17736 31748
rect 18420 31764 18472 31816
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 10508 31628 10560 31680
rect 13544 31628 13596 31680
rect 15292 31628 15344 31680
rect 15568 31671 15620 31680
rect 15568 31637 15577 31671
rect 15577 31637 15611 31671
rect 15611 31637 15620 31671
rect 15568 31628 15620 31637
rect 17776 31628 17828 31680
rect 18788 31628 18840 31680
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 23664 31832 23716 31884
rect 25872 31900 25924 31952
rect 26424 31943 26476 31952
rect 26424 31909 26433 31943
rect 26433 31909 26467 31943
rect 26467 31909 26476 31943
rect 26424 31900 26476 31909
rect 26516 31900 26568 31952
rect 27712 31943 27764 31952
rect 27712 31909 27721 31943
rect 27721 31909 27755 31943
rect 27755 31909 27764 31943
rect 27712 31900 27764 31909
rect 26332 31764 26384 31816
rect 26424 31807 26476 31816
rect 26424 31773 26433 31807
rect 26433 31773 26467 31807
rect 26467 31773 26476 31807
rect 26424 31764 26476 31773
rect 26608 31807 26660 31816
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 21548 31628 21600 31680
rect 23940 31696 23992 31748
rect 27344 31764 27396 31816
rect 23388 31671 23440 31680
rect 23388 31637 23397 31671
rect 23397 31637 23431 31671
rect 23431 31637 23440 31671
rect 23388 31628 23440 31637
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 3148 31424 3200 31476
rect 4528 31424 4580 31476
rect 5172 31467 5224 31476
rect 5172 31433 5181 31467
rect 5181 31433 5215 31467
rect 5215 31433 5224 31467
rect 5172 31424 5224 31433
rect 7840 31467 7892 31476
rect 7840 31433 7849 31467
rect 7849 31433 7883 31467
rect 7883 31433 7892 31467
rect 7840 31424 7892 31433
rect 9036 31424 9088 31476
rect 2504 31331 2556 31340
rect 2504 31297 2513 31331
rect 2513 31297 2547 31331
rect 2547 31297 2556 31331
rect 2504 31288 2556 31297
rect 4804 31331 4856 31340
rect 4804 31297 4813 31331
rect 4813 31297 4847 31331
rect 4847 31297 4856 31331
rect 4804 31288 4856 31297
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 6092 31288 6144 31340
rect 7196 31356 7248 31408
rect 10140 31356 10192 31408
rect 3056 31220 3108 31272
rect 5724 31220 5776 31272
rect 6460 31220 6512 31272
rect 6644 31263 6696 31272
rect 6644 31229 6653 31263
rect 6653 31229 6687 31263
rect 6687 31229 6696 31263
rect 9036 31288 9088 31340
rect 9404 31331 9456 31340
rect 9404 31297 9438 31331
rect 9438 31297 9456 31331
rect 9404 31288 9456 31297
rect 6644 31220 6696 31229
rect 7472 31263 7524 31272
rect 7472 31229 7481 31263
rect 7481 31229 7515 31263
rect 7515 31229 7524 31263
rect 7472 31220 7524 31229
rect 9128 31263 9180 31272
rect 9128 31229 9137 31263
rect 9137 31229 9171 31263
rect 9171 31229 9180 31263
rect 9128 31220 9180 31229
rect 11704 31424 11756 31476
rect 13820 31424 13872 31476
rect 16488 31424 16540 31476
rect 17408 31424 17460 31476
rect 19064 31424 19116 31476
rect 14740 31356 14792 31408
rect 12440 31288 12492 31340
rect 13360 31331 13412 31340
rect 13360 31297 13394 31331
rect 13394 31297 13412 31331
rect 13360 31288 13412 31297
rect 15476 31288 15528 31340
rect 13084 31263 13136 31272
rect 13084 31229 13093 31263
rect 13093 31229 13127 31263
rect 13127 31229 13136 31263
rect 13084 31220 13136 31229
rect 14556 31220 14608 31272
rect 16580 31288 16632 31340
rect 17500 31263 17552 31272
rect 17500 31229 17509 31263
rect 17509 31229 17543 31263
rect 17543 31229 17552 31263
rect 17500 31220 17552 31229
rect 3240 31152 3292 31204
rect 7840 31195 7892 31204
rect 7840 31161 7849 31195
rect 7849 31161 7883 31195
rect 7883 31161 7892 31195
rect 7840 31152 7892 31161
rect 16672 31152 16724 31204
rect 1584 31084 1636 31136
rect 2504 31084 2556 31136
rect 4344 31084 4396 31136
rect 10232 31084 10284 31136
rect 10416 31084 10468 31136
rect 10600 31084 10652 31136
rect 13728 31084 13780 31136
rect 14464 31127 14516 31136
rect 14464 31093 14473 31127
rect 14473 31093 14507 31127
rect 14507 31093 14516 31127
rect 14464 31084 14516 31093
rect 15200 31084 15252 31136
rect 17224 31084 17276 31136
rect 19340 31263 19392 31272
rect 19340 31229 19349 31263
rect 19349 31229 19383 31263
rect 19383 31229 19392 31263
rect 19340 31220 19392 31229
rect 21732 31424 21784 31476
rect 21640 31288 21692 31340
rect 23664 31288 23716 31340
rect 21548 31220 21600 31272
rect 24676 31331 24728 31340
rect 24676 31297 24685 31331
rect 24685 31297 24719 31331
rect 24719 31297 24728 31331
rect 24676 31288 24728 31297
rect 24952 31288 25004 31340
rect 25964 31288 26016 31340
rect 26240 31220 26292 31272
rect 26792 31288 26844 31340
rect 20720 31195 20772 31204
rect 20720 31161 20729 31195
rect 20729 31161 20763 31195
rect 20763 31161 20772 31195
rect 20720 31152 20772 31161
rect 20996 31152 21048 31204
rect 18696 31084 18748 31136
rect 21456 31084 21508 31136
rect 25780 31152 25832 31204
rect 26516 31084 26568 31136
rect 26792 31084 26844 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 9956 30923 10008 30932
rect 9956 30889 9965 30923
rect 9965 30889 9999 30923
rect 9999 30889 10008 30923
rect 9956 30880 10008 30889
rect 13728 30923 13780 30932
rect 13728 30889 13737 30923
rect 13737 30889 13771 30923
rect 13771 30889 13780 30923
rect 13728 30880 13780 30889
rect 13820 30880 13872 30932
rect 3884 30812 3936 30864
rect 6092 30855 6144 30864
rect 6092 30821 6101 30855
rect 6101 30821 6135 30855
rect 6135 30821 6144 30855
rect 6092 30812 6144 30821
rect 3332 30787 3384 30796
rect 3332 30753 3341 30787
rect 3341 30753 3375 30787
rect 3375 30753 3384 30787
rect 3332 30744 3384 30753
rect 13084 30812 13136 30864
rect 9036 30744 9088 30796
rect 13636 30744 13688 30796
rect 13728 30787 13780 30796
rect 13728 30753 13737 30787
rect 13737 30753 13771 30787
rect 13771 30753 13780 30787
rect 13728 30744 13780 30753
rect 16488 30855 16540 30864
rect 16488 30821 16497 30855
rect 16497 30821 16531 30855
rect 16531 30821 16540 30855
rect 18236 30880 18288 30932
rect 18788 30880 18840 30932
rect 18880 30880 18932 30932
rect 16488 30812 16540 30821
rect 19524 30812 19576 30864
rect 15384 30744 15436 30796
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 2412 30676 2464 30728
rect 4344 30651 4396 30660
rect 4344 30617 4353 30651
rect 4353 30617 4387 30651
rect 4387 30617 4396 30651
rect 4344 30608 4396 30617
rect 5724 30719 5776 30728
rect 5724 30685 5733 30719
rect 5733 30685 5767 30719
rect 5767 30685 5776 30719
rect 6552 30719 6604 30728
rect 5724 30676 5776 30685
rect 6552 30685 6561 30719
rect 6561 30685 6595 30719
rect 6595 30685 6604 30719
rect 6552 30676 6604 30685
rect 6828 30676 6880 30728
rect 8300 30676 8352 30728
rect 9680 30676 9732 30728
rect 10140 30676 10192 30728
rect 10600 30676 10652 30728
rect 6736 30608 6788 30660
rect 12716 30608 12768 30660
rect 4252 30540 4304 30592
rect 5172 30540 5224 30592
rect 7472 30540 7524 30592
rect 11704 30540 11756 30592
rect 12900 30608 12952 30660
rect 15568 30676 15620 30728
rect 17684 30744 17736 30796
rect 18052 30744 18104 30796
rect 21548 30880 21600 30932
rect 22284 30880 22336 30932
rect 23940 30880 23992 30932
rect 25136 30880 25188 30932
rect 26240 30880 26292 30932
rect 27804 30855 27856 30864
rect 27804 30821 27813 30855
rect 27813 30821 27847 30855
rect 27847 30821 27856 30855
rect 27804 30812 27856 30821
rect 15936 30608 15988 30660
rect 14648 30540 14700 30592
rect 15292 30540 15344 30592
rect 15476 30540 15528 30592
rect 15660 30540 15712 30592
rect 17776 30676 17828 30728
rect 17960 30719 18012 30728
rect 17960 30685 17969 30719
rect 17969 30685 18003 30719
rect 18003 30685 18012 30719
rect 17960 30676 18012 30685
rect 17868 30608 17920 30660
rect 19432 30676 19484 30728
rect 20720 30608 20772 30660
rect 21456 30676 21508 30728
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23572 30676 23624 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 25964 30744 26016 30796
rect 24952 30676 25004 30728
rect 27068 30744 27120 30796
rect 17408 30540 17460 30592
rect 21732 30608 21784 30660
rect 22376 30540 22428 30592
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 3976 30336 4028 30388
rect 5540 30336 5592 30388
rect 7564 30336 7616 30388
rect 9956 30336 10008 30388
rect 12072 30379 12124 30388
rect 12072 30345 12081 30379
rect 12081 30345 12115 30379
rect 12115 30345 12124 30379
rect 12072 30336 12124 30345
rect 12164 30336 12216 30388
rect 2136 30311 2188 30320
rect 2136 30277 2145 30311
rect 2145 30277 2179 30311
rect 2179 30277 2188 30311
rect 2136 30268 2188 30277
rect 7012 30268 7064 30320
rect 7656 30268 7708 30320
rect 1952 30243 2004 30252
rect 1952 30209 1961 30243
rect 1961 30209 1995 30243
rect 1995 30209 2004 30243
rect 1952 30200 2004 30209
rect 2044 30243 2096 30252
rect 2044 30209 2053 30243
rect 2053 30209 2087 30243
rect 2087 30209 2096 30243
rect 2044 30200 2096 30209
rect 1860 29996 1912 30048
rect 2320 30200 2372 30252
rect 2872 30243 2924 30252
rect 2872 30209 2881 30243
rect 2881 30209 2915 30243
rect 2915 30209 2924 30243
rect 2872 30200 2924 30209
rect 4896 30200 4948 30252
rect 4804 30132 4856 30184
rect 6000 30132 6052 30184
rect 6828 30200 6880 30252
rect 10140 30268 10192 30320
rect 10692 30268 10744 30320
rect 7104 30132 7156 30184
rect 7656 30175 7708 30184
rect 7656 30141 7665 30175
rect 7665 30141 7699 30175
rect 7699 30141 7708 30175
rect 7656 30132 7708 30141
rect 12072 30243 12124 30252
rect 12072 30209 12081 30243
rect 12081 30209 12115 30243
rect 12115 30209 12124 30243
rect 12072 30200 12124 30209
rect 13084 30268 13136 30320
rect 13452 30336 13504 30388
rect 14188 30336 14240 30388
rect 14464 30336 14516 30388
rect 14832 30336 14884 30388
rect 15752 30336 15804 30388
rect 15384 30268 15436 30320
rect 15936 30268 15988 30320
rect 17132 30311 17184 30320
rect 17132 30277 17166 30311
rect 17166 30277 17184 30311
rect 17132 30268 17184 30277
rect 17684 30336 17736 30388
rect 18696 30336 18748 30388
rect 20720 30379 20772 30388
rect 20720 30345 20729 30379
rect 20729 30345 20763 30379
rect 20763 30345 20772 30379
rect 20720 30336 20772 30345
rect 18144 30268 18196 30320
rect 13728 30200 13780 30252
rect 15292 30200 15344 30252
rect 20904 30243 20956 30252
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 22192 30336 22244 30388
rect 23204 30336 23256 30388
rect 23480 30268 23532 30320
rect 9772 30175 9824 30184
rect 9772 30141 9781 30175
rect 9781 30141 9815 30175
rect 9815 30141 9824 30175
rect 9772 30132 9824 30141
rect 11704 30175 11756 30184
rect 11704 30141 11713 30175
rect 11713 30141 11747 30175
rect 11747 30141 11756 30175
rect 11704 30132 11756 30141
rect 14464 30132 14516 30184
rect 14740 30132 14792 30184
rect 15476 30175 15528 30184
rect 15476 30141 15485 30175
rect 15485 30141 15519 30175
rect 15519 30141 15528 30175
rect 15476 30132 15528 30141
rect 5816 30064 5868 30116
rect 7380 30064 7432 30116
rect 9588 29996 9640 30048
rect 11980 30064 12032 30116
rect 10692 29996 10744 30048
rect 11152 30039 11204 30048
rect 11152 30005 11161 30039
rect 11161 30005 11195 30039
rect 11195 30005 11204 30039
rect 11152 29996 11204 30005
rect 11796 29996 11848 30048
rect 12532 29996 12584 30048
rect 15844 30107 15896 30116
rect 15844 30073 15853 30107
rect 15853 30073 15887 30107
rect 15887 30073 15896 30107
rect 15844 30064 15896 30073
rect 15568 29996 15620 30048
rect 15936 29996 15988 30048
rect 16120 29996 16172 30048
rect 18236 30132 18288 30184
rect 19432 30132 19484 30184
rect 20720 30132 20772 30184
rect 23664 30200 23716 30252
rect 24584 30200 24636 30252
rect 22560 30132 22612 30184
rect 24860 30243 24912 30252
rect 24860 30209 24869 30243
rect 24869 30209 24903 30243
rect 24903 30209 24912 30243
rect 24860 30200 24912 30209
rect 26240 30268 26292 30320
rect 25964 30243 26016 30252
rect 25964 30209 25997 30243
rect 25997 30209 26016 30243
rect 25964 30200 26016 30209
rect 26056 30200 26108 30252
rect 27068 30200 27120 30252
rect 27988 30243 28040 30252
rect 27988 30209 27997 30243
rect 27997 30209 28031 30243
rect 28031 30209 28040 30243
rect 27988 30200 28040 30209
rect 26792 30132 26844 30184
rect 17132 29996 17184 30048
rect 17500 29996 17552 30048
rect 17592 29996 17644 30048
rect 22744 30064 22796 30116
rect 18144 29996 18196 30048
rect 21916 29996 21968 30048
rect 23020 29996 23072 30048
rect 27804 30039 27856 30048
rect 27804 30005 27813 30039
rect 27813 30005 27847 30039
rect 27847 30005 27856 30039
rect 27804 29996 27856 30005
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 2780 29835 2832 29844
rect 2780 29801 2789 29835
rect 2789 29801 2823 29835
rect 2823 29801 2832 29835
rect 2780 29792 2832 29801
rect 4068 29792 4120 29844
rect 11060 29792 11112 29844
rect 11980 29792 12032 29844
rect 3240 29724 3292 29776
rect 5264 29767 5316 29776
rect 5264 29733 5273 29767
rect 5273 29733 5307 29767
rect 5307 29733 5316 29767
rect 5264 29724 5316 29733
rect 6092 29767 6144 29776
rect 6092 29733 6101 29767
rect 6101 29733 6135 29767
rect 6135 29733 6144 29767
rect 6092 29724 6144 29733
rect 8576 29724 8628 29776
rect 14556 29767 14608 29776
rect 14556 29733 14565 29767
rect 14565 29733 14599 29767
rect 14599 29733 14608 29767
rect 14556 29724 14608 29733
rect 14924 29724 14976 29776
rect 16488 29792 16540 29844
rect 17868 29792 17920 29844
rect 18052 29792 18104 29844
rect 21548 29792 21600 29844
rect 16764 29724 16816 29776
rect 3148 29656 3200 29708
rect 5724 29699 5776 29708
rect 5724 29665 5733 29699
rect 5733 29665 5767 29699
rect 5767 29665 5776 29699
rect 5724 29656 5776 29665
rect 2412 29631 2464 29640
rect 2412 29597 2421 29631
rect 2421 29597 2455 29631
rect 2455 29597 2464 29631
rect 2412 29588 2464 29597
rect 1952 29520 2004 29572
rect 4160 29588 4212 29640
rect 4988 29588 5040 29640
rect 5356 29588 5408 29640
rect 8300 29656 8352 29708
rect 14096 29656 14148 29708
rect 22560 29792 22612 29844
rect 22744 29792 22796 29844
rect 26148 29792 26200 29844
rect 5724 29520 5776 29572
rect 1492 29452 1544 29504
rect 2044 29452 2096 29504
rect 5172 29452 5224 29504
rect 7472 29588 7524 29640
rect 8484 29452 8536 29504
rect 9128 29588 9180 29640
rect 11244 29588 11296 29640
rect 13728 29631 13780 29640
rect 13728 29597 13737 29631
rect 13737 29597 13771 29631
rect 13771 29597 13780 29631
rect 13728 29588 13780 29597
rect 14280 29588 14332 29640
rect 14556 29588 14608 29640
rect 15016 29631 15068 29640
rect 15016 29597 15025 29631
rect 15025 29597 15059 29631
rect 15059 29597 15068 29631
rect 15016 29588 15068 29597
rect 16396 29588 16448 29640
rect 17132 29631 17184 29640
rect 17132 29597 17141 29631
rect 17141 29597 17175 29631
rect 17175 29597 17184 29631
rect 17132 29588 17184 29597
rect 17224 29588 17276 29640
rect 12256 29520 12308 29572
rect 15936 29520 15988 29572
rect 16120 29520 16172 29572
rect 10140 29452 10192 29504
rect 11888 29452 11940 29504
rect 15476 29452 15528 29504
rect 16948 29520 17000 29572
rect 19432 29631 19484 29640
rect 19432 29597 19441 29631
rect 19441 29597 19475 29631
rect 19475 29597 19484 29631
rect 19432 29588 19484 29597
rect 19524 29588 19576 29640
rect 21916 29588 21968 29640
rect 26516 29724 26568 29776
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 23848 29631 23900 29640
rect 23848 29597 23857 29631
rect 23857 29597 23891 29631
rect 23891 29597 23900 29631
rect 23848 29588 23900 29597
rect 24584 29588 24636 29640
rect 26608 29588 26660 29640
rect 27620 29588 27672 29640
rect 19340 29452 19392 29504
rect 20536 29452 20588 29504
rect 20628 29452 20680 29504
rect 24492 29520 24544 29572
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 2596 29248 2648 29300
rect 3792 29223 3844 29232
rect 3792 29189 3801 29223
rect 3801 29189 3835 29223
rect 3835 29189 3844 29223
rect 3792 29180 3844 29189
rect 3976 29223 4028 29232
rect 3976 29189 3985 29223
rect 3985 29189 4019 29223
rect 4019 29189 4028 29223
rect 3976 29180 4028 29189
rect 4804 29112 4856 29164
rect 5172 29248 5224 29300
rect 8484 29248 8536 29300
rect 9128 29248 9180 29300
rect 5264 29112 5316 29164
rect 4712 29087 4764 29096
rect 4712 29053 4721 29087
rect 4721 29053 4755 29087
rect 4755 29053 4764 29087
rect 4712 29044 4764 29053
rect 4988 29044 5040 29096
rect 12072 29180 12124 29232
rect 13636 29248 13688 29300
rect 14372 29248 14424 29300
rect 15384 29248 15436 29300
rect 14096 29180 14148 29232
rect 14832 29180 14884 29232
rect 15200 29180 15252 29232
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 7196 29112 7248 29164
rect 7564 29112 7616 29164
rect 8300 29112 8352 29164
rect 8760 29112 8812 29164
rect 9220 29112 9272 29164
rect 12164 29112 12216 29164
rect 13636 29112 13688 29164
rect 13728 29112 13780 29164
rect 15384 29112 15436 29164
rect 6552 29087 6604 29096
rect 6552 29053 6561 29087
rect 6561 29053 6595 29087
rect 6595 29053 6604 29087
rect 6552 29044 6604 29053
rect 4160 29019 4212 29028
rect 4160 28985 4169 29019
rect 4169 28985 4203 29019
rect 4203 28985 4212 29019
rect 4160 28976 4212 28985
rect 5540 28976 5592 29028
rect 6736 28976 6788 29028
rect 8576 29019 8628 29028
rect 8576 28985 8585 29019
rect 8585 28985 8619 29019
rect 8619 28985 8628 29019
rect 8576 28976 8628 28985
rect 9036 28976 9088 29028
rect 10508 29019 10560 29028
rect 10508 28985 10517 29019
rect 10517 28985 10551 29019
rect 10551 28985 10560 29019
rect 10508 28976 10560 28985
rect 10692 29019 10744 29028
rect 10692 28985 10701 29019
rect 10701 28985 10735 29019
rect 10735 28985 10744 29019
rect 10692 28976 10744 28985
rect 12348 29087 12400 29096
rect 12348 29053 12357 29087
rect 12357 29053 12391 29087
rect 12391 29053 12400 29087
rect 12348 29044 12400 29053
rect 14464 29044 14516 29096
rect 15476 29044 15528 29096
rect 5448 28908 5500 28960
rect 7012 28908 7064 28960
rect 14832 28976 14884 29028
rect 15200 28976 15252 29028
rect 16488 29248 16540 29300
rect 16672 29248 16724 29300
rect 19340 29248 19392 29300
rect 20904 29248 20956 29300
rect 16764 29180 16816 29232
rect 18144 29180 18196 29232
rect 18604 29180 18656 29232
rect 18972 29180 19024 29232
rect 22284 29248 22336 29300
rect 22836 29248 22888 29300
rect 24952 29248 25004 29300
rect 17040 29112 17092 29164
rect 17132 29112 17184 29164
rect 21548 29180 21600 29232
rect 25872 29223 25924 29232
rect 25872 29189 25881 29223
rect 25881 29189 25915 29223
rect 25915 29189 25924 29223
rect 25872 29180 25924 29189
rect 27160 29248 27212 29300
rect 17224 29044 17276 29096
rect 14280 28908 14332 28960
rect 14372 28908 14424 28960
rect 16212 28976 16264 29028
rect 15936 28908 15988 28960
rect 18236 28908 18288 28960
rect 18604 28908 18656 28960
rect 19432 29112 19484 29164
rect 21456 29112 21508 29164
rect 22100 29112 22152 29164
rect 21088 29044 21140 29096
rect 22836 29155 22888 29164
rect 22836 29121 22845 29155
rect 22845 29121 22879 29155
rect 22879 29121 22888 29155
rect 22836 29112 22888 29121
rect 23664 29044 23716 29096
rect 19156 28976 19208 29028
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 26516 29112 26568 29164
rect 26700 29180 26752 29232
rect 19708 28908 19760 28960
rect 20444 28908 20496 28960
rect 23480 28951 23532 28960
rect 23480 28917 23489 28951
rect 23489 28917 23523 28951
rect 23523 28917 23532 28951
rect 23480 28908 23532 28917
rect 23664 28908 23716 28960
rect 26240 29044 26292 29096
rect 27068 29112 27120 29164
rect 27896 29112 27948 29164
rect 24952 28976 25004 29028
rect 25596 28976 25648 29028
rect 25688 28908 25740 28960
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 7196 28704 7248 28756
rect 7748 28636 7800 28688
rect 3884 28568 3936 28620
rect 9680 28636 9732 28688
rect 10968 28636 11020 28688
rect 1860 28500 1912 28552
rect 3240 28500 3292 28552
rect 4804 28500 4856 28552
rect 6828 28543 6880 28552
rect 6828 28509 6837 28543
rect 6837 28509 6871 28543
rect 6871 28509 6880 28543
rect 6828 28500 6880 28509
rect 7472 28543 7524 28552
rect 7472 28509 7481 28543
rect 7481 28509 7515 28543
rect 7515 28509 7524 28543
rect 7472 28500 7524 28509
rect 11152 28568 11204 28620
rect 12164 28568 12216 28620
rect 4988 28432 5040 28484
rect 5080 28432 5132 28484
rect 9864 28543 9916 28552
rect 9864 28509 9873 28543
rect 9873 28509 9907 28543
rect 9907 28509 9916 28543
rect 9864 28500 9916 28509
rect 1952 28364 2004 28416
rect 3148 28407 3200 28416
rect 3148 28373 3157 28407
rect 3157 28373 3191 28407
rect 3191 28373 3200 28407
rect 3148 28364 3200 28373
rect 4252 28407 4304 28416
rect 4252 28373 4261 28407
rect 4261 28373 4295 28407
rect 4295 28373 4304 28407
rect 4252 28364 4304 28373
rect 4344 28364 4396 28416
rect 9680 28432 9732 28484
rect 9128 28364 9180 28416
rect 11888 28500 11940 28552
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 10968 28364 11020 28416
rect 12624 28364 12676 28416
rect 13636 28500 13688 28552
rect 14004 28636 14056 28688
rect 14648 28636 14700 28688
rect 16028 28704 16080 28756
rect 21088 28704 21140 28756
rect 21456 28747 21508 28756
rect 21456 28713 21465 28747
rect 21465 28713 21499 28747
rect 21499 28713 21508 28747
rect 21456 28704 21508 28713
rect 23848 28704 23900 28756
rect 17408 28636 17460 28688
rect 17960 28636 18012 28688
rect 18696 28636 18748 28688
rect 18972 28636 19024 28688
rect 26056 28704 26108 28756
rect 26240 28636 26292 28688
rect 14096 28568 14148 28620
rect 15660 28543 15712 28552
rect 15660 28509 15669 28543
rect 15669 28509 15703 28543
rect 15703 28509 15712 28543
rect 15660 28500 15712 28509
rect 17040 28500 17092 28552
rect 17868 28500 17920 28552
rect 19524 28500 19576 28552
rect 13728 28364 13780 28416
rect 14832 28364 14884 28416
rect 18236 28432 18288 28484
rect 18328 28432 18380 28484
rect 20352 28500 20404 28552
rect 21272 28500 21324 28552
rect 19708 28432 19760 28484
rect 18696 28364 18748 28416
rect 22100 28432 22152 28484
rect 23664 28500 23716 28552
rect 24584 28543 24636 28552
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 25596 28568 25648 28620
rect 25780 28500 25832 28552
rect 25872 28432 25924 28484
rect 20628 28364 20680 28416
rect 25044 28364 25096 28416
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 2320 28160 2372 28212
rect 3148 28160 3200 28212
rect 1768 28067 1820 28076
rect 1768 28033 1777 28067
rect 1777 28033 1811 28067
rect 1811 28033 1820 28067
rect 1768 28024 1820 28033
rect 3884 28092 3936 28144
rect 5172 28160 5224 28212
rect 7196 28203 7248 28212
rect 7196 28169 7205 28203
rect 7205 28169 7239 28203
rect 7239 28169 7248 28203
rect 7196 28160 7248 28169
rect 7380 28160 7432 28212
rect 9128 28203 9180 28212
rect 9128 28169 9137 28203
rect 9137 28169 9171 28203
rect 9171 28169 9180 28203
rect 9128 28160 9180 28169
rect 11888 28203 11940 28212
rect 11888 28169 11897 28203
rect 11897 28169 11931 28203
rect 11931 28169 11940 28203
rect 11888 28160 11940 28169
rect 14188 28160 14240 28212
rect 15752 28160 15804 28212
rect 16212 28160 16264 28212
rect 1952 28024 2004 28076
rect 4068 28024 4120 28076
rect 5172 28024 5224 28076
rect 2044 27999 2096 28008
rect 2044 27965 2053 27999
rect 2053 27965 2087 27999
rect 2087 27965 2096 27999
rect 2044 27956 2096 27965
rect 5264 27956 5316 28008
rect 3700 27888 3752 27940
rect 5724 28024 5776 28076
rect 6828 28024 6880 28076
rect 7012 28024 7064 28076
rect 7380 28024 7432 28076
rect 8484 28092 8536 28144
rect 6000 27999 6052 28008
rect 6000 27965 6009 27999
rect 6009 27965 6043 27999
rect 6043 27965 6052 27999
rect 6000 27956 6052 27965
rect 5908 27931 5960 27940
rect 5908 27897 5917 27931
rect 5917 27897 5951 27931
rect 5951 27897 5960 27931
rect 5908 27888 5960 27897
rect 7472 27956 7524 28008
rect 8760 27999 8812 28008
rect 8760 27965 8769 27999
rect 8769 27965 8803 27999
rect 8803 27965 8812 27999
rect 8760 27956 8812 27965
rect 7012 27888 7064 27940
rect 11704 28092 11756 28144
rect 9220 28024 9272 28076
rect 14372 28092 14424 28144
rect 14096 28067 14148 28076
rect 14096 28033 14105 28067
rect 14105 28033 14139 28067
rect 14139 28033 14148 28067
rect 14096 28024 14148 28033
rect 14464 28024 14516 28076
rect 15108 28067 15160 28076
rect 15108 28033 15117 28067
rect 15117 28033 15151 28067
rect 15151 28033 15160 28067
rect 15108 28024 15160 28033
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 17408 28092 17460 28144
rect 18512 28092 18564 28144
rect 16764 28024 16816 28076
rect 18972 28160 19024 28212
rect 19984 28160 20036 28212
rect 20628 28160 20680 28212
rect 21456 28160 21508 28212
rect 24676 28160 24728 28212
rect 24768 28203 24820 28212
rect 24768 28169 24777 28203
rect 24777 28169 24811 28203
rect 24811 28169 24820 28203
rect 24768 28160 24820 28169
rect 25136 28160 25188 28212
rect 26056 28160 26108 28212
rect 26332 28160 26384 28212
rect 22376 28092 22428 28144
rect 7196 27820 7248 27872
rect 9036 27820 9088 27872
rect 10968 27956 11020 28008
rect 11244 27956 11296 28008
rect 14372 27956 14424 28008
rect 13268 27888 13320 27940
rect 15476 27956 15528 28008
rect 16212 27956 16264 28008
rect 15108 27888 15160 27940
rect 9772 27820 9824 27872
rect 9956 27820 10008 27872
rect 15660 27820 15712 27872
rect 16028 27888 16080 27940
rect 16488 27888 16540 27940
rect 18328 27888 18380 27940
rect 17592 27820 17644 27872
rect 19064 28067 19116 28076
rect 19064 28033 19073 28067
rect 19073 28033 19107 28067
rect 19107 28033 19116 28067
rect 19064 28024 19116 28033
rect 19432 28024 19484 28076
rect 20628 28024 20680 28076
rect 24860 28024 24912 28076
rect 25136 28024 25188 28076
rect 25596 28067 25648 28076
rect 25596 28033 25605 28067
rect 25605 28033 25639 28067
rect 25639 28033 25648 28067
rect 25596 28024 25648 28033
rect 26056 28067 26108 28076
rect 26056 28033 26065 28067
rect 26065 28033 26099 28067
rect 26099 28033 26108 28067
rect 26056 28024 26108 28033
rect 26424 28024 26476 28076
rect 27620 28024 27672 28076
rect 19248 27956 19300 28008
rect 19524 27956 19576 28008
rect 19800 27956 19852 28008
rect 19064 27820 19116 27872
rect 19892 27820 19944 27872
rect 22652 27820 22704 27872
rect 24032 27820 24084 27872
rect 24124 27820 24176 27872
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 480 27616 532 27668
rect 3608 27616 3660 27668
rect 9772 27616 9824 27668
rect 10048 27616 10100 27668
rect 11704 27616 11756 27668
rect 12072 27616 12124 27668
rect 13820 27616 13872 27668
rect 14372 27616 14424 27668
rect 18052 27616 18104 27668
rect 3976 27548 4028 27600
rect 4068 27591 4120 27600
rect 4068 27557 4077 27591
rect 4077 27557 4111 27591
rect 4111 27557 4120 27591
rect 4068 27548 4120 27557
rect 5172 27548 5224 27600
rect 5724 27548 5776 27600
rect 7472 27548 7524 27600
rect 6920 27523 6972 27532
rect 6920 27489 6929 27523
rect 6929 27489 6963 27523
rect 6963 27489 6972 27523
rect 6920 27480 6972 27489
rect 1952 27412 2004 27464
rect 1768 27344 1820 27396
rect 4252 27455 4304 27464
rect 4252 27421 4261 27455
rect 4261 27421 4295 27455
rect 4295 27421 4304 27455
rect 4252 27412 4304 27421
rect 2412 27344 2464 27396
rect 4988 27412 5040 27464
rect 5264 27455 5316 27464
rect 5264 27421 5273 27455
rect 5273 27421 5307 27455
rect 5307 27421 5316 27455
rect 5264 27412 5316 27421
rect 5540 27412 5592 27464
rect 5632 27412 5684 27464
rect 6000 27412 6052 27464
rect 4896 27344 4948 27396
rect 6276 27455 6328 27464
rect 6276 27421 6285 27455
rect 6285 27421 6319 27455
rect 6319 27421 6328 27455
rect 6276 27412 6328 27421
rect 9864 27480 9916 27532
rect 12624 27548 12676 27600
rect 15292 27548 15344 27600
rect 19248 27548 19300 27600
rect 20720 27548 20772 27600
rect 20904 27616 20956 27668
rect 26240 27616 26292 27668
rect 21548 27548 21600 27600
rect 22008 27548 22060 27600
rect 9128 27412 9180 27464
rect 7012 27344 7064 27396
rect 3332 27276 3384 27328
rect 5724 27276 5776 27328
rect 6368 27276 6420 27328
rect 6644 27276 6696 27328
rect 7472 27276 7524 27328
rect 8392 27276 8444 27328
rect 9220 27276 9272 27328
rect 10048 27412 10100 27464
rect 11244 27412 11296 27464
rect 9588 27344 9640 27396
rect 10784 27344 10836 27396
rect 15752 27523 15804 27532
rect 15752 27489 15761 27523
rect 15761 27489 15795 27523
rect 15795 27489 15804 27523
rect 15752 27480 15804 27489
rect 12348 27455 12400 27464
rect 12348 27421 12357 27455
rect 12357 27421 12391 27455
rect 12391 27421 12400 27455
rect 12348 27412 12400 27421
rect 12624 27412 12676 27464
rect 13176 27455 13228 27464
rect 13176 27421 13185 27455
rect 13185 27421 13219 27455
rect 13219 27421 13228 27455
rect 13176 27412 13228 27421
rect 11704 27276 11756 27328
rect 12808 27276 12860 27328
rect 13912 27412 13964 27464
rect 14372 27412 14424 27464
rect 15476 27412 15528 27464
rect 20168 27480 20220 27532
rect 14556 27387 14608 27396
rect 14556 27353 14565 27387
rect 14565 27353 14599 27387
rect 14599 27353 14608 27387
rect 14556 27344 14608 27353
rect 15200 27344 15252 27396
rect 15752 27319 15804 27328
rect 15752 27285 15761 27319
rect 15761 27285 15795 27319
rect 15795 27285 15804 27319
rect 15752 27276 15804 27285
rect 17316 27276 17368 27328
rect 17868 27412 17920 27464
rect 18420 27344 18472 27396
rect 20812 27412 20864 27464
rect 20904 27455 20956 27464
rect 20904 27421 20913 27455
rect 20913 27421 20947 27455
rect 20947 27421 20956 27455
rect 20904 27412 20956 27421
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 22008 27455 22060 27464
rect 22008 27421 22017 27455
rect 22017 27421 22051 27455
rect 22051 27421 22060 27455
rect 22008 27412 22060 27421
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 22652 27412 22704 27421
rect 19340 27276 19392 27328
rect 19616 27276 19668 27328
rect 20076 27276 20128 27328
rect 20628 27276 20680 27328
rect 21640 27344 21692 27396
rect 22376 27344 22428 27396
rect 24676 27412 24728 27464
rect 21548 27319 21600 27328
rect 21548 27285 21557 27319
rect 21557 27285 21591 27319
rect 21591 27285 21600 27319
rect 21548 27276 21600 27285
rect 22192 27276 22244 27328
rect 22284 27276 22336 27328
rect 24124 27276 24176 27328
rect 25136 27276 25188 27328
rect 27620 27276 27672 27328
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 2872 27072 2924 27124
rect 2504 27004 2556 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 2136 26911 2188 26920
rect 2136 26877 2145 26911
rect 2145 26877 2179 26911
rect 2179 26877 2188 26911
rect 2136 26868 2188 26877
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 6092 27004 6144 27056
rect 9128 27072 9180 27124
rect 9312 27115 9364 27124
rect 9312 27081 9321 27115
rect 9321 27081 9355 27115
rect 9355 27081 9364 27115
rect 9312 27072 9364 27081
rect 10232 27072 10284 27124
rect 12624 27072 12676 27124
rect 12808 27072 12860 27124
rect 14096 27072 14148 27124
rect 14556 27072 14608 27124
rect 14740 27004 14792 27056
rect 15384 27072 15436 27124
rect 16580 27072 16632 27124
rect 16856 27072 16908 27124
rect 17960 27072 18012 27124
rect 19064 27072 19116 27124
rect 19340 27072 19392 27124
rect 19432 27115 19484 27124
rect 19432 27081 19441 27115
rect 19441 27081 19475 27115
rect 19475 27081 19484 27115
rect 19432 27072 19484 27081
rect 19524 27072 19576 27124
rect 20996 27072 21048 27124
rect 15476 27004 15528 27056
rect 15844 27004 15896 27056
rect 3516 26868 3568 26920
rect 6644 26936 6696 26988
rect 7012 26936 7064 26988
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 6184 26868 6236 26920
rect 6828 26868 6880 26920
rect 7656 26868 7708 26920
rect 8484 26936 8536 26988
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 9404 26868 9456 26920
rect 10324 26911 10376 26920
rect 10324 26877 10333 26911
rect 10333 26877 10367 26911
rect 10367 26877 10376 26911
rect 10324 26868 10376 26877
rect 11152 26979 11204 26988
rect 11152 26945 11161 26979
rect 11161 26945 11195 26979
rect 11195 26945 11204 26979
rect 11152 26936 11204 26945
rect 12348 26979 12400 26988
rect 12348 26945 12357 26979
rect 12357 26945 12391 26979
rect 12391 26945 12400 26979
rect 13176 26979 13228 26988
rect 12348 26936 12400 26945
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 14096 26936 14148 26945
rect 14188 26936 14240 26988
rect 15108 26979 15160 26988
rect 15108 26945 15117 26979
rect 15117 26945 15151 26979
rect 15151 26945 15160 26979
rect 15108 26936 15160 26945
rect 15384 26936 15436 26988
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 21640 27004 21692 27056
rect 22376 27004 22428 27056
rect 23204 27004 23256 27056
rect 17960 26936 18012 26988
rect 18052 26979 18104 26988
rect 18052 26945 18061 26979
rect 18061 26945 18095 26979
rect 18095 26945 18104 26979
rect 18052 26936 18104 26945
rect 4068 26843 4120 26852
rect 4068 26809 4077 26843
rect 4077 26809 4111 26843
rect 4111 26809 4120 26843
rect 4068 26800 4120 26809
rect 4160 26800 4212 26852
rect 5908 26843 5960 26852
rect 5908 26809 5917 26843
rect 5917 26809 5951 26843
rect 5951 26809 5960 26843
rect 5908 26800 5960 26809
rect 7012 26843 7064 26852
rect 7012 26809 7021 26843
rect 7021 26809 7055 26843
rect 7055 26809 7064 26843
rect 7012 26800 7064 26809
rect 17868 26868 17920 26920
rect 11980 26800 12032 26852
rect 12808 26800 12860 26852
rect 13636 26800 13688 26852
rect 16304 26800 16356 26852
rect 16580 26800 16632 26852
rect 17224 26800 17276 26852
rect 19432 26936 19484 26988
rect 19616 26979 19668 26988
rect 19616 26945 19617 26979
rect 19617 26945 19651 26979
rect 19651 26945 19668 26979
rect 19616 26936 19668 26945
rect 18420 26868 18472 26920
rect 18696 26868 18748 26920
rect 20720 26936 20772 26988
rect 21180 26936 21232 26988
rect 24308 26936 24360 26988
rect 21548 26868 21600 26920
rect 24768 26936 24820 26988
rect 25872 26936 25924 26988
rect 24952 26868 25004 26920
rect 28080 26936 28132 26988
rect 9220 26732 9272 26784
rect 15108 26732 15160 26784
rect 17684 26732 17736 26784
rect 17868 26732 17920 26784
rect 19340 26732 19392 26784
rect 19616 26732 19668 26784
rect 20444 26732 20496 26784
rect 20536 26732 20588 26784
rect 23388 26775 23440 26784
rect 23388 26741 23397 26775
rect 23397 26741 23431 26775
rect 23431 26741 23440 26775
rect 23388 26732 23440 26741
rect 23756 26732 23808 26784
rect 23940 26732 23992 26784
rect 25964 26732 26016 26784
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 3792 26528 3844 26580
rect 6000 26528 6052 26580
rect 8392 26528 8444 26580
rect 4160 26435 4212 26444
rect 4160 26401 4169 26435
rect 4169 26401 4203 26435
rect 4203 26401 4212 26435
rect 4160 26392 4212 26401
rect 4988 26460 5040 26512
rect 5816 26460 5868 26512
rect 6460 26392 6512 26444
rect 7288 26460 7340 26512
rect 1768 26324 1820 26376
rect 5080 26324 5132 26376
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 5356 26324 5408 26376
rect 6368 26324 6420 26376
rect 6920 26324 6972 26376
rect 1676 26299 1728 26308
rect 1676 26265 1685 26299
rect 1685 26265 1719 26299
rect 1719 26265 1728 26299
rect 1676 26256 1728 26265
rect 4068 26299 4120 26308
rect 4068 26265 4077 26299
rect 4077 26265 4111 26299
rect 4111 26265 4120 26299
rect 4068 26256 4120 26265
rect 4988 26256 5040 26308
rect 6644 26299 6696 26308
rect 6644 26265 6653 26299
rect 6653 26265 6687 26299
rect 6687 26265 6696 26299
rect 6644 26256 6696 26265
rect 5724 26188 5776 26240
rect 8668 26460 8720 26512
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 7748 26367 7800 26376
rect 7748 26333 7757 26367
rect 7757 26333 7791 26367
rect 7791 26333 7800 26367
rect 7748 26324 7800 26333
rect 9588 26528 9640 26580
rect 10784 26528 10836 26580
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 11888 26460 11940 26512
rect 8576 26231 8628 26240
rect 8576 26197 8585 26231
rect 8585 26197 8619 26231
rect 8619 26197 8628 26231
rect 8576 26188 8628 26197
rect 9312 26188 9364 26240
rect 9864 26392 9916 26444
rect 9956 26324 10008 26376
rect 10416 26367 10468 26376
rect 10416 26333 10425 26367
rect 10425 26333 10459 26367
rect 10459 26333 10468 26367
rect 10416 26324 10468 26333
rect 10692 26324 10744 26376
rect 12348 26392 12400 26444
rect 13268 26435 13320 26444
rect 13268 26401 13277 26435
rect 13277 26401 13311 26435
rect 13311 26401 13320 26435
rect 13268 26392 13320 26401
rect 14004 26528 14056 26580
rect 20904 26528 20956 26580
rect 21088 26528 21140 26580
rect 13636 26503 13688 26512
rect 13636 26469 13645 26503
rect 13645 26469 13679 26503
rect 13679 26469 13688 26503
rect 13636 26460 13688 26469
rect 14464 26460 14516 26512
rect 15108 26460 15160 26512
rect 14648 26392 14700 26444
rect 14832 26367 14884 26376
rect 14832 26333 14841 26367
rect 14841 26333 14875 26367
rect 14875 26333 14884 26367
rect 14832 26324 14884 26333
rect 16120 26460 16172 26512
rect 17960 26460 18012 26512
rect 19248 26460 19300 26512
rect 22928 26460 22980 26512
rect 23388 26460 23440 26512
rect 17684 26392 17736 26444
rect 16120 26324 16172 26376
rect 16488 26367 16540 26376
rect 16488 26333 16497 26367
rect 16497 26333 16531 26367
rect 16531 26333 16540 26367
rect 16488 26324 16540 26333
rect 17316 26324 17368 26376
rect 10324 26299 10376 26308
rect 10324 26265 10333 26299
rect 10333 26265 10367 26299
rect 10367 26265 10376 26299
rect 10324 26256 10376 26265
rect 11060 26256 11112 26308
rect 12992 26256 13044 26308
rect 15936 26256 15988 26308
rect 16028 26256 16080 26308
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 10784 26188 10836 26240
rect 11428 26188 11480 26240
rect 13636 26231 13688 26240
rect 13636 26197 13645 26231
rect 13645 26197 13679 26231
rect 13679 26197 13688 26231
rect 13636 26188 13688 26197
rect 14648 26188 14700 26240
rect 15292 26188 15344 26240
rect 15476 26231 15528 26240
rect 15476 26197 15485 26231
rect 15485 26197 15519 26231
rect 15519 26197 15528 26231
rect 15476 26188 15528 26197
rect 19800 26256 19852 26308
rect 22284 26324 22336 26376
rect 20904 26256 20956 26308
rect 21640 26256 21692 26308
rect 22468 26324 22520 26376
rect 22744 26324 22796 26376
rect 23112 26367 23164 26376
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23296 26324 23348 26333
rect 24676 26392 24728 26444
rect 18788 26188 18840 26240
rect 19432 26188 19484 26240
rect 20352 26188 20404 26240
rect 20812 26231 20864 26240
rect 20812 26197 20821 26231
rect 20821 26197 20855 26231
rect 20855 26197 20864 26231
rect 20812 26188 20864 26197
rect 20996 26188 21048 26240
rect 22652 26231 22704 26240
rect 22652 26197 22661 26231
rect 22661 26197 22695 26231
rect 22695 26197 22704 26231
rect 22652 26188 22704 26197
rect 23204 26299 23256 26308
rect 23204 26265 23213 26299
rect 23213 26265 23247 26299
rect 23247 26265 23256 26299
rect 23204 26256 23256 26265
rect 26148 26324 26200 26376
rect 23848 26299 23900 26308
rect 23848 26265 23857 26299
rect 23857 26265 23891 26299
rect 23891 26265 23900 26299
rect 23848 26256 23900 26265
rect 24860 26256 24912 26308
rect 26516 26231 26568 26240
rect 26516 26197 26525 26231
rect 26525 26197 26559 26231
rect 26559 26197 26568 26231
rect 26516 26188 26568 26197
rect 28356 26231 28408 26240
rect 28356 26197 28365 26231
rect 28365 26197 28399 26231
rect 28399 26197 28408 26231
rect 28356 26188 28408 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 2412 26027 2464 26036
rect 2412 25993 2421 26027
rect 2421 25993 2455 26027
rect 2455 25993 2464 26027
rect 2412 25984 2464 25993
rect 5908 25984 5960 26036
rect 7472 25984 7524 26036
rect 8576 25984 8628 26036
rect 9496 25984 9548 26036
rect 9772 26027 9824 26036
rect 9772 25993 9781 26027
rect 9781 25993 9815 26027
rect 9815 25993 9824 26027
rect 9772 25984 9824 25993
rect 9864 26027 9916 26036
rect 9864 25993 9873 26027
rect 9873 25993 9907 26027
rect 9907 25993 9916 26027
rect 9864 25984 9916 25993
rect 11152 25984 11204 26036
rect 11428 25984 11480 26036
rect 3424 25959 3476 25968
rect 3424 25925 3433 25959
rect 3433 25925 3467 25959
rect 3467 25925 3476 25959
rect 3424 25916 3476 25925
rect 9128 25916 9180 25968
rect 1400 25780 1452 25832
rect 1860 25780 1912 25832
rect 2320 25780 2372 25832
rect 3700 25848 3752 25900
rect 4804 25848 4856 25900
rect 5632 25891 5684 25900
rect 5632 25857 5641 25891
rect 5641 25857 5675 25891
rect 5675 25857 5684 25891
rect 5632 25848 5684 25857
rect 6460 25848 6512 25900
rect 2964 25823 3016 25832
rect 2964 25789 2973 25823
rect 2973 25789 3007 25823
rect 3007 25789 3016 25823
rect 2964 25780 3016 25789
rect 8208 25848 8260 25900
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 9312 25916 9364 25968
rect 16948 25916 17000 25968
rect 18604 25916 18656 25968
rect 20076 25984 20128 26036
rect 25044 25984 25096 26036
rect 20996 25916 21048 25968
rect 22284 25959 22336 25968
rect 22284 25925 22307 25959
rect 22307 25925 22336 25959
rect 22284 25916 22336 25925
rect 10508 25848 10560 25900
rect 1676 25712 1728 25764
rect 2596 25712 2648 25764
rect 5908 25755 5960 25764
rect 5908 25721 5917 25755
rect 5917 25721 5951 25755
rect 5951 25721 5960 25755
rect 5908 25712 5960 25721
rect 6920 25712 6972 25764
rect 7840 25712 7892 25764
rect 8116 25755 8168 25764
rect 8116 25721 8125 25755
rect 8125 25721 8159 25755
rect 8159 25721 8168 25755
rect 8116 25712 8168 25721
rect 8576 25823 8628 25832
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 9036 25780 9088 25832
rect 9496 25780 9548 25832
rect 9588 25780 9640 25832
rect 10968 25848 11020 25900
rect 12532 25848 12584 25900
rect 12716 25891 12768 25900
rect 12716 25857 12750 25891
rect 12750 25857 12768 25891
rect 12716 25848 12768 25857
rect 13452 25848 13504 25900
rect 16212 25848 16264 25900
rect 16488 25848 16540 25900
rect 16672 25848 16724 25900
rect 17500 25848 17552 25900
rect 17868 25848 17920 25900
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 20076 25848 20128 25900
rect 20536 25848 20588 25900
rect 23020 25916 23072 25968
rect 23204 25916 23256 25968
rect 24952 25916 25004 25968
rect 25596 25916 25648 25968
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 12440 25780 12492 25789
rect 17776 25780 17828 25832
rect 18236 25780 18288 25832
rect 18604 25780 18656 25832
rect 19248 25780 19300 25832
rect 11152 25712 11204 25764
rect 12256 25712 12308 25764
rect 18144 25712 18196 25764
rect 21180 25780 21232 25832
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 7288 25644 7340 25653
rect 7656 25644 7708 25696
rect 7932 25644 7984 25696
rect 9680 25644 9732 25696
rect 10968 25644 11020 25696
rect 12808 25644 12860 25696
rect 14464 25644 14516 25696
rect 16304 25687 16356 25696
rect 16304 25653 16313 25687
rect 16313 25653 16347 25687
rect 16347 25653 16356 25687
rect 16304 25644 16356 25653
rect 19340 25644 19392 25696
rect 22744 25848 22796 25900
rect 21548 25780 21600 25832
rect 23480 25848 23532 25900
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 22008 25644 22060 25696
rect 22376 25644 22428 25696
rect 22744 25644 22796 25696
rect 25872 25755 25924 25764
rect 25872 25721 25881 25755
rect 25881 25721 25915 25755
rect 25915 25721 25924 25755
rect 25872 25712 25924 25721
rect 24584 25644 24636 25696
rect 24952 25644 25004 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 7472 25440 7524 25492
rect 8208 25440 8260 25492
rect 8760 25440 8812 25492
rect 10600 25440 10652 25492
rect 12532 25440 12584 25492
rect 13084 25440 13136 25492
rect 15016 25483 15068 25492
rect 15016 25449 15025 25483
rect 15025 25449 15059 25483
rect 15059 25449 15068 25483
rect 15016 25440 15068 25449
rect 17868 25483 17920 25492
rect 17868 25449 17877 25483
rect 17877 25449 17911 25483
rect 17911 25449 17920 25483
rect 17868 25440 17920 25449
rect 19248 25440 19300 25492
rect 19800 25483 19852 25492
rect 19800 25449 19809 25483
rect 19809 25449 19843 25483
rect 19843 25449 19852 25483
rect 19800 25440 19852 25449
rect 20904 25440 20956 25492
rect 5540 25372 5592 25424
rect 5908 25304 5960 25356
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 2044 25236 2096 25288
rect 2504 25236 2556 25288
rect 6828 25372 6880 25424
rect 6368 25304 6420 25356
rect 8576 25304 8628 25356
rect 9772 25304 9824 25356
rect 10416 25372 10468 25424
rect 10968 25372 11020 25424
rect 13820 25372 13872 25424
rect 16028 25372 16080 25424
rect 16120 25372 16172 25424
rect 21272 25372 21324 25424
rect 22008 25483 22060 25492
rect 22008 25449 22017 25483
rect 22017 25449 22051 25483
rect 22051 25449 22060 25483
rect 22008 25440 22060 25449
rect 22560 25440 22612 25492
rect 23204 25440 23256 25492
rect 24124 25440 24176 25492
rect 25688 25440 25740 25492
rect 27620 25440 27672 25492
rect 24768 25372 24820 25424
rect 6460 25279 6512 25288
rect 6460 25245 6495 25279
rect 6495 25245 6512 25279
rect 6460 25236 6512 25245
rect 6736 25236 6788 25288
rect 7932 25236 7984 25288
rect 9220 25279 9272 25288
rect 9220 25245 9229 25279
rect 9229 25245 9263 25279
rect 9263 25245 9272 25279
rect 9220 25236 9272 25245
rect 9496 25236 9548 25288
rect 18052 25304 18104 25356
rect 10048 25236 10100 25288
rect 12440 25236 12492 25288
rect 12624 25236 12676 25288
rect 14004 25236 14056 25288
rect 14188 25236 14240 25288
rect 1860 25168 1912 25220
rect 5356 25143 5408 25152
rect 5356 25109 5365 25143
rect 5365 25109 5399 25143
rect 5399 25109 5408 25143
rect 5356 25100 5408 25109
rect 7288 25168 7340 25220
rect 7840 25168 7892 25220
rect 6552 25100 6604 25152
rect 6828 25100 6880 25152
rect 6920 25100 6972 25152
rect 8208 25100 8260 25152
rect 8392 25143 8444 25152
rect 8392 25109 8401 25143
rect 8401 25109 8435 25143
rect 8435 25109 8444 25143
rect 8392 25100 8444 25109
rect 8484 25100 8536 25152
rect 8760 25168 8812 25220
rect 9680 25168 9732 25220
rect 10968 25168 11020 25220
rect 11060 25168 11112 25220
rect 10416 25100 10468 25152
rect 10508 25100 10560 25152
rect 12440 25100 12492 25152
rect 13176 25100 13228 25152
rect 13728 25168 13780 25220
rect 15384 25236 15436 25288
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 16856 25236 16908 25288
rect 15292 25168 15344 25220
rect 17684 25211 17736 25220
rect 17684 25177 17693 25211
rect 17693 25177 17727 25211
rect 17727 25177 17736 25211
rect 17684 25168 17736 25177
rect 14096 25100 14148 25152
rect 14188 25100 14240 25152
rect 16488 25100 16540 25152
rect 17224 25100 17276 25152
rect 18052 25168 18104 25220
rect 19248 25304 19300 25356
rect 20628 25304 20680 25356
rect 19340 25236 19392 25288
rect 21088 25236 21140 25288
rect 22468 25236 22520 25288
rect 18972 25168 19024 25220
rect 19892 25168 19944 25220
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 23572 25168 23624 25220
rect 26056 25279 26108 25288
rect 26056 25245 26065 25279
rect 26065 25245 26099 25279
rect 26099 25245 26108 25279
rect 26056 25236 26108 25245
rect 26424 25168 26476 25220
rect 23664 25100 23716 25152
rect 24676 25143 24728 25152
rect 24676 25109 24685 25143
rect 24685 25109 24719 25143
rect 24719 25109 24728 25143
rect 24676 25100 24728 25109
rect 27436 25143 27488 25152
rect 27436 25109 27445 25143
rect 27445 25109 27479 25143
rect 27479 25109 27488 25143
rect 27436 25100 27488 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 1860 24939 1912 24948
rect 1860 24905 1869 24939
rect 1869 24905 1903 24939
rect 1903 24905 1912 24939
rect 1860 24896 1912 24905
rect 5264 24896 5316 24948
rect 6092 24896 6144 24948
rect 6460 24896 6512 24948
rect 2964 24828 3016 24880
rect 1400 24760 1452 24812
rect 1860 24803 1912 24812
rect 1860 24769 1869 24803
rect 1869 24769 1903 24803
rect 1903 24769 1912 24803
rect 1860 24760 1912 24769
rect 4068 24760 4120 24812
rect 5448 24828 5500 24880
rect 5356 24760 5408 24812
rect 6000 24828 6052 24880
rect 6368 24828 6420 24880
rect 6552 24871 6604 24880
rect 6552 24837 6561 24871
rect 6561 24837 6595 24871
rect 6595 24837 6604 24871
rect 6552 24828 6604 24837
rect 7380 24896 7432 24948
rect 7840 24896 7892 24948
rect 8760 24896 8812 24948
rect 9312 24896 9364 24948
rect 10416 24896 10468 24948
rect 10784 24896 10836 24948
rect 11336 24896 11388 24948
rect 12164 24896 12216 24948
rect 12440 24896 12492 24948
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 6920 24760 6972 24812
rect 8484 24828 8536 24880
rect 8852 24828 8904 24880
rect 2044 24692 2096 24744
rect 2504 24692 2556 24744
rect 3332 24556 3384 24608
rect 7288 24692 7340 24744
rect 7380 24692 7432 24744
rect 9312 24760 9364 24812
rect 9496 24760 9548 24812
rect 11060 24828 11112 24880
rect 10048 24692 10100 24744
rect 10508 24760 10560 24812
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 10968 24760 11020 24812
rect 12900 24828 12952 24880
rect 15292 24828 15344 24880
rect 20076 24896 20128 24948
rect 23388 24896 23440 24948
rect 26608 24896 26660 24948
rect 10784 24692 10836 24744
rect 12624 24760 12676 24812
rect 13544 24760 13596 24812
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 15752 24803 15804 24812
rect 15752 24769 15762 24803
rect 15762 24769 15796 24803
rect 15796 24769 15804 24803
rect 15752 24760 15804 24769
rect 15936 24803 15988 24812
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 16028 24803 16080 24812
rect 16028 24769 16037 24803
rect 16037 24769 16071 24803
rect 16071 24769 16080 24803
rect 16028 24760 16080 24769
rect 16120 24803 16172 24812
rect 16120 24769 16134 24803
rect 16134 24769 16168 24803
rect 16168 24769 16172 24803
rect 24584 24828 24636 24880
rect 25044 24828 25096 24880
rect 25596 24828 25648 24880
rect 16120 24760 16172 24769
rect 17684 24760 17736 24812
rect 16396 24692 16448 24744
rect 17776 24692 17828 24744
rect 6368 24624 6420 24676
rect 7932 24624 7984 24676
rect 8852 24624 8904 24676
rect 12808 24624 12860 24676
rect 14556 24624 14608 24676
rect 16948 24624 17000 24676
rect 4068 24556 4120 24608
rect 4896 24556 4948 24608
rect 6000 24556 6052 24608
rect 8668 24556 8720 24608
rect 8760 24599 8812 24608
rect 8760 24565 8769 24599
rect 8769 24565 8803 24599
rect 8803 24565 8812 24599
rect 8760 24556 8812 24565
rect 9036 24556 9088 24608
rect 11336 24556 11388 24608
rect 11520 24556 11572 24608
rect 12900 24556 12952 24608
rect 15568 24556 15620 24608
rect 17960 24624 18012 24676
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 19064 24760 19116 24812
rect 20076 24760 20128 24812
rect 21364 24760 21416 24812
rect 19340 24692 19392 24744
rect 18788 24624 18840 24676
rect 19524 24692 19576 24744
rect 23020 24760 23072 24812
rect 21548 24692 21600 24744
rect 22008 24735 22060 24744
rect 22008 24701 22017 24735
rect 22017 24701 22051 24735
rect 22051 24701 22060 24735
rect 22008 24692 22060 24701
rect 23756 24692 23808 24744
rect 18972 24556 19024 24608
rect 19616 24624 19668 24676
rect 20904 24556 20956 24608
rect 20996 24599 21048 24608
rect 20996 24565 21005 24599
rect 21005 24565 21039 24599
rect 21039 24565 21048 24599
rect 20996 24556 21048 24565
rect 23480 24624 23532 24676
rect 24860 24624 24912 24676
rect 23388 24599 23440 24608
rect 23388 24565 23397 24599
rect 23397 24565 23431 24599
rect 23431 24565 23440 24599
rect 23388 24556 23440 24565
rect 24492 24599 24544 24608
rect 24492 24565 24501 24599
rect 24501 24565 24535 24599
rect 24535 24565 24544 24599
rect 24492 24556 24544 24565
rect 25872 24556 25924 24608
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 3516 24352 3568 24404
rect 5448 24352 5500 24404
rect 5632 24352 5684 24404
rect 7656 24352 7708 24404
rect 7840 24352 7892 24404
rect 8576 24352 8628 24404
rect 9588 24352 9640 24404
rect 10508 24284 10560 24336
rect 10600 24284 10652 24336
rect 10968 24352 11020 24404
rect 17316 24352 17368 24404
rect 17776 24395 17828 24404
rect 17776 24361 17785 24395
rect 17785 24361 17819 24395
rect 17819 24361 17828 24395
rect 17776 24352 17828 24361
rect 19524 24352 19576 24404
rect 2044 24191 2096 24200
rect 2044 24157 2053 24191
rect 2053 24157 2087 24191
rect 2087 24157 2096 24191
rect 2044 24148 2096 24157
rect 2136 24148 2188 24200
rect 3884 24148 3936 24200
rect 4712 24148 4764 24200
rect 4988 24148 5040 24200
rect 5264 24148 5316 24200
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 5908 24216 5960 24268
rect 7656 24216 7708 24268
rect 8852 24216 8904 24268
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 9036 24148 9088 24200
rect 9128 24148 9180 24200
rect 4344 24123 4396 24132
rect 4344 24089 4353 24123
rect 4353 24089 4387 24123
rect 4387 24089 4396 24123
rect 4344 24080 4396 24089
rect 6000 24080 6052 24132
rect 6092 24080 6144 24132
rect 6552 24123 6604 24132
rect 6552 24089 6561 24123
rect 6561 24089 6595 24123
rect 6595 24089 6604 24123
rect 6552 24080 6604 24089
rect 3056 24012 3108 24064
rect 4804 24012 4856 24064
rect 6460 24012 6512 24064
rect 8300 24123 8352 24132
rect 8300 24089 8309 24123
rect 8309 24089 8343 24123
rect 8343 24089 8352 24123
rect 8300 24080 8352 24089
rect 9588 24123 9640 24132
rect 9588 24089 9597 24123
rect 9597 24089 9631 24123
rect 9631 24089 9640 24123
rect 9588 24080 9640 24089
rect 10508 24148 10560 24200
rect 10784 24148 10836 24200
rect 11336 24148 11388 24200
rect 11612 24080 11664 24132
rect 8392 24012 8444 24064
rect 8484 24012 8536 24064
rect 12072 24216 12124 24268
rect 15200 24284 15252 24336
rect 17408 24284 17460 24336
rect 18236 24284 18288 24336
rect 18328 24284 18380 24336
rect 18880 24284 18932 24336
rect 19064 24284 19116 24336
rect 19800 24284 19852 24336
rect 20628 24352 20680 24404
rect 24952 24352 25004 24404
rect 11888 24148 11940 24200
rect 12256 24191 12308 24200
rect 12256 24157 12266 24191
rect 12266 24157 12300 24191
rect 12300 24157 12308 24191
rect 12256 24148 12308 24157
rect 12624 24191 12676 24200
rect 12624 24157 12638 24191
rect 12638 24157 12672 24191
rect 12672 24157 12676 24191
rect 12624 24148 12676 24157
rect 13912 24148 13964 24200
rect 11796 24012 11848 24064
rect 13268 24080 13320 24132
rect 13728 24080 13780 24132
rect 14096 24012 14148 24064
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 15384 24216 15436 24268
rect 16948 24216 17000 24268
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 15016 24191 15068 24200
rect 15016 24157 15025 24191
rect 15025 24157 15059 24191
rect 15059 24157 15068 24191
rect 15016 24148 15068 24157
rect 16212 24148 16264 24200
rect 16488 24148 16540 24200
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 18144 24148 18196 24200
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 14464 24080 14516 24132
rect 16120 24080 16172 24132
rect 18972 24216 19024 24268
rect 19432 24216 19484 24268
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 20996 24284 21048 24336
rect 21456 24284 21508 24336
rect 23664 24327 23716 24336
rect 23664 24293 23673 24327
rect 23673 24293 23707 24327
rect 23707 24293 23716 24327
rect 23664 24284 23716 24293
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24216 21600 24268
rect 22008 24216 22060 24268
rect 26056 24216 26108 24268
rect 22836 24148 22888 24200
rect 23296 24148 23348 24200
rect 25136 24148 25188 24200
rect 16948 24012 17000 24064
rect 17408 24012 17460 24064
rect 19524 24080 19576 24132
rect 22376 24080 22428 24132
rect 22560 24123 22612 24132
rect 22560 24089 22594 24123
rect 22594 24089 22612 24123
rect 22560 24080 22612 24089
rect 23204 24080 23256 24132
rect 23940 24080 23992 24132
rect 24860 24123 24912 24132
rect 24860 24089 24894 24123
rect 24894 24089 24912 24123
rect 24860 24080 24912 24089
rect 26516 24148 26568 24200
rect 21272 24012 21324 24064
rect 21364 24055 21416 24064
rect 21364 24021 21373 24055
rect 21373 24021 21407 24055
rect 21407 24021 21416 24055
rect 21364 24012 21416 24021
rect 23112 24012 23164 24064
rect 26240 24080 26292 24132
rect 25596 24012 25648 24064
rect 27804 24055 27856 24064
rect 27804 24021 27813 24055
rect 27813 24021 27847 24055
rect 27847 24021 27856 24055
rect 27804 24012 27856 24021
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 1768 23783 1820 23792
rect 1768 23749 1777 23783
rect 1777 23749 1811 23783
rect 1811 23749 1820 23783
rect 1768 23740 1820 23749
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 2596 23783 2648 23792
rect 2596 23749 2605 23783
rect 2605 23749 2639 23783
rect 2639 23749 2648 23783
rect 2596 23740 2648 23749
rect 2964 23808 3016 23860
rect 3884 23851 3936 23860
rect 3884 23817 3893 23851
rect 3893 23817 3927 23851
rect 3927 23817 3936 23851
rect 3884 23808 3936 23817
rect 4436 23808 4488 23860
rect 4620 23808 4672 23860
rect 3424 23672 3476 23724
rect 3976 23740 4028 23792
rect 6276 23808 6328 23860
rect 6368 23808 6420 23860
rect 6736 23808 6788 23860
rect 7288 23808 7340 23860
rect 9864 23808 9916 23860
rect 10600 23808 10652 23860
rect 11244 23808 11296 23860
rect 3884 23672 3936 23724
rect 5724 23740 5776 23792
rect 4712 23604 4764 23656
rect 480 23536 532 23588
rect 4068 23536 4120 23588
rect 6460 23672 6512 23724
rect 6368 23604 6420 23656
rect 7012 23672 7064 23724
rect 7380 23672 7432 23724
rect 8852 23715 8904 23724
rect 8852 23681 8879 23715
rect 8879 23681 8904 23715
rect 8852 23672 8904 23681
rect 9772 23672 9824 23724
rect 10784 23783 10836 23792
rect 10784 23749 10793 23783
rect 10793 23749 10827 23783
rect 10827 23749 10836 23783
rect 10784 23740 10836 23749
rect 11980 23740 12032 23792
rect 13452 23808 13504 23860
rect 13820 23851 13872 23860
rect 13820 23817 13829 23851
rect 13829 23817 13863 23851
rect 13863 23817 13872 23851
rect 13820 23808 13872 23817
rect 14740 23808 14792 23860
rect 7840 23604 7892 23656
rect 8392 23647 8444 23656
rect 8392 23613 8401 23647
rect 8401 23613 8435 23647
rect 8435 23613 8444 23647
rect 8392 23604 8444 23613
rect 8576 23647 8628 23656
rect 8576 23613 8585 23647
rect 8585 23613 8619 23647
rect 8619 23613 8628 23647
rect 8576 23604 8628 23613
rect 6920 23579 6972 23588
rect 6920 23545 6929 23579
rect 6929 23545 6963 23579
rect 6963 23545 6972 23579
rect 6920 23536 6972 23545
rect 4160 23468 4212 23520
rect 4896 23468 4948 23520
rect 7932 23468 7984 23520
rect 9312 23604 9364 23656
rect 9864 23604 9916 23656
rect 10048 23647 10100 23656
rect 10048 23613 10057 23647
rect 10057 23613 10091 23647
rect 10091 23613 10100 23647
rect 10048 23604 10100 23613
rect 10232 23647 10284 23656
rect 10232 23613 10241 23647
rect 10241 23613 10275 23647
rect 10275 23613 10284 23647
rect 10232 23604 10284 23613
rect 13544 23740 13596 23792
rect 12900 23672 12952 23724
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 9772 23536 9824 23588
rect 9588 23468 9640 23520
rect 11060 23604 11112 23656
rect 11888 23604 11940 23656
rect 12440 23604 12492 23656
rect 13268 23672 13320 23724
rect 15200 23740 15252 23792
rect 17960 23808 18012 23860
rect 18144 23808 18196 23860
rect 18696 23808 18748 23860
rect 15016 23672 15068 23724
rect 14464 23604 14516 23656
rect 14740 23604 14792 23656
rect 16304 23740 16356 23792
rect 16856 23740 16908 23792
rect 17316 23740 17368 23792
rect 18052 23740 18104 23792
rect 15936 23672 15988 23724
rect 17316 23604 17368 23656
rect 17776 23715 17828 23724
rect 17776 23681 17785 23715
rect 17785 23681 17819 23715
rect 17819 23681 17828 23715
rect 17776 23672 17828 23681
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 19984 23808 20036 23860
rect 20168 23808 20220 23860
rect 22284 23808 22336 23860
rect 22376 23808 22428 23860
rect 24768 23808 24820 23860
rect 28356 23808 28408 23860
rect 18972 23715 19024 23724
rect 18972 23681 18981 23715
rect 18981 23681 19015 23715
rect 19015 23681 19024 23715
rect 18972 23672 19024 23681
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 20260 23672 20312 23724
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 23020 23604 23072 23656
rect 12532 23536 12584 23588
rect 12900 23536 12952 23588
rect 10508 23468 10560 23520
rect 14832 23511 14884 23520
rect 14832 23477 14841 23511
rect 14841 23477 14875 23511
rect 14875 23477 14884 23511
rect 14832 23468 14884 23477
rect 15660 23511 15712 23520
rect 15660 23477 15669 23511
rect 15669 23477 15703 23511
rect 15703 23477 15712 23511
rect 15660 23468 15712 23477
rect 16212 23468 16264 23520
rect 20444 23536 20496 23588
rect 21272 23536 21324 23588
rect 23572 23740 23624 23792
rect 23296 23672 23348 23724
rect 23480 23715 23532 23724
rect 23480 23681 23514 23715
rect 23514 23681 23532 23715
rect 23480 23672 23532 23681
rect 24216 23672 24268 23724
rect 20720 23468 20772 23520
rect 23940 23468 23992 23520
rect 24124 23468 24176 23520
rect 24492 23468 24544 23520
rect 26148 23468 26200 23520
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 1860 23264 1912 23316
rect 4068 23307 4120 23316
rect 4068 23273 4077 23307
rect 4077 23273 4111 23307
rect 4111 23273 4120 23307
rect 4068 23264 4120 23273
rect 2412 23196 2464 23248
rect 2964 23128 3016 23180
rect 3700 23128 3752 23180
rect 5816 23264 5868 23316
rect 1860 23060 1912 23112
rect 1308 22992 1360 23044
rect 2964 23035 3016 23044
rect 2964 23001 2973 23035
rect 2973 23001 3007 23035
rect 3007 23001 3016 23035
rect 2964 22992 3016 23001
rect 4436 23103 4488 23112
rect 4436 23069 4445 23103
rect 4445 23069 4479 23103
rect 4479 23069 4488 23103
rect 4436 23060 4488 23069
rect 4620 23060 4672 23112
rect 4988 23060 5040 23112
rect 6552 23196 6604 23248
rect 7380 23264 7432 23316
rect 8392 23264 8444 23316
rect 9680 23264 9732 23316
rect 10876 23264 10928 23316
rect 11796 23264 11848 23316
rect 12164 23264 12216 23316
rect 12808 23264 12860 23316
rect 10784 23196 10836 23248
rect 11244 23196 11296 23248
rect 12900 23196 12952 23248
rect 14556 23264 14608 23316
rect 15016 23264 15068 23316
rect 15752 23264 15804 23316
rect 16028 23307 16080 23316
rect 16028 23273 16037 23307
rect 16037 23273 16071 23307
rect 16071 23273 16080 23307
rect 16028 23264 16080 23273
rect 16396 23264 16448 23316
rect 17592 23264 17644 23316
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 20076 23264 20128 23316
rect 14372 23196 14424 23248
rect 14648 23239 14700 23248
rect 14648 23205 14657 23239
rect 14657 23205 14691 23239
rect 14691 23205 14700 23239
rect 14648 23196 14700 23205
rect 6644 23128 6696 23180
rect 5540 23103 5592 23112
rect 5540 23069 5549 23103
rect 5549 23069 5583 23103
rect 5583 23069 5592 23103
rect 5540 23060 5592 23069
rect 5724 23060 5776 23112
rect 6000 23060 6052 23112
rect 5816 22992 5868 23044
rect 6828 23060 6880 23112
rect 7932 23128 7984 23180
rect 9312 23128 9364 23180
rect 7840 23103 7892 23112
rect 7840 23069 7849 23103
rect 7849 23069 7883 23103
rect 7883 23069 7892 23103
rect 7840 23060 7892 23069
rect 11060 23128 11112 23180
rect 7196 22992 7248 23044
rect 10416 23060 10468 23112
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 12348 23128 12400 23180
rect 14004 23128 14056 23180
rect 14556 23128 14608 23180
rect 15384 23196 15436 23248
rect 18512 23196 18564 23248
rect 19156 23196 19208 23248
rect 19708 23239 19760 23248
rect 19708 23205 19717 23239
rect 19717 23205 19751 23239
rect 19751 23205 19760 23239
rect 19708 23196 19760 23205
rect 19984 23196 20036 23248
rect 22836 23264 22888 23316
rect 23296 23264 23348 23316
rect 24860 23264 24912 23316
rect 22468 23196 22520 23248
rect 12164 23103 12216 23112
rect 12164 23069 12171 23103
rect 12171 23069 12216 23103
rect 12164 23060 12216 23069
rect 12440 23103 12492 23112
rect 12440 23069 12454 23103
rect 12454 23069 12488 23103
rect 12488 23069 12492 23103
rect 12440 23060 12492 23069
rect 12624 23060 12676 23112
rect 16764 23128 16816 23180
rect 18696 23128 18748 23180
rect 2504 22924 2556 22976
rect 3056 22924 3108 22976
rect 4068 22924 4120 22976
rect 4252 22924 4304 22976
rect 6092 22967 6144 22976
rect 6092 22933 6101 22967
rect 6101 22933 6135 22967
rect 6135 22933 6144 22967
rect 6092 22924 6144 22933
rect 6184 22924 6236 22976
rect 9128 22967 9180 22976
rect 9128 22933 9137 22967
rect 9137 22933 9171 22967
rect 9171 22933 9180 22967
rect 9128 22924 9180 22933
rect 9588 22967 9640 22976
rect 9588 22933 9597 22967
rect 9597 22933 9631 22967
rect 9631 22933 9640 22967
rect 9588 22924 9640 22933
rect 10324 22924 10376 22976
rect 10508 22924 10560 22976
rect 11888 22924 11940 22976
rect 12072 22924 12124 22976
rect 12348 23035 12400 23044
rect 12348 23001 12357 23035
rect 12357 23001 12391 23035
rect 12391 23001 12400 23035
rect 12348 22992 12400 23001
rect 13176 22992 13228 23044
rect 14280 23035 14332 23044
rect 14280 23001 14289 23035
rect 14289 23001 14323 23035
rect 14323 23001 14332 23035
rect 14280 22992 14332 23001
rect 16212 23060 16264 23112
rect 15752 22992 15804 23044
rect 16580 22992 16632 23044
rect 17132 23060 17184 23112
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 17868 23060 17920 23112
rect 19340 23060 19392 23112
rect 20168 23060 20220 23112
rect 22376 23128 22428 23180
rect 13452 22924 13504 22976
rect 13544 22967 13596 22976
rect 13544 22933 13569 22967
rect 13569 22933 13596 22967
rect 13544 22924 13596 22933
rect 15292 22924 15344 22976
rect 16856 22924 16908 22976
rect 18604 22992 18656 23044
rect 19432 23035 19484 23044
rect 19432 23001 19441 23035
rect 19441 23001 19475 23035
rect 19475 23001 19484 23035
rect 19432 22992 19484 23001
rect 20076 22992 20128 23044
rect 18788 22924 18840 22976
rect 19156 22924 19208 22976
rect 19340 22924 19392 22976
rect 19892 22924 19944 22976
rect 23020 23060 23072 23112
rect 23296 22992 23348 23044
rect 24400 22992 24452 23044
rect 24032 22924 24084 22976
rect 25780 22924 25832 22976
rect 26148 23060 26200 23112
rect 26516 22992 26568 23044
rect 26424 22924 26476 22976
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 1768 22720 1820 22772
rect 2688 22720 2740 22772
rect 2136 22584 2188 22636
rect 3240 22584 3292 22636
rect 3700 22720 3752 22772
rect 3700 22627 3752 22636
rect 3700 22593 3709 22627
rect 3709 22593 3743 22627
rect 3743 22593 3752 22627
rect 3700 22584 3752 22593
rect 4988 22720 5040 22772
rect 5540 22720 5592 22772
rect 7748 22720 7800 22772
rect 6184 22652 6236 22704
rect 6460 22652 6512 22704
rect 10324 22720 10376 22772
rect 11796 22720 11848 22772
rect 12348 22720 12400 22772
rect 13728 22720 13780 22772
rect 14096 22720 14148 22772
rect 15384 22720 15436 22772
rect 17776 22720 17828 22772
rect 17960 22720 18012 22772
rect 2044 22516 2096 22568
rect 3976 22516 4028 22568
rect 4068 22516 4120 22568
rect 9036 22584 9088 22636
rect 4988 22516 5040 22568
rect 4344 22448 4396 22500
rect 2412 22380 2464 22432
rect 2872 22380 2924 22432
rect 3240 22423 3292 22432
rect 3240 22389 3249 22423
rect 3249 22389 3283 22423
rect 3283 22389 3292 22423
rect 3240 22380 3292 22389
rect 3516 22380 3568 22432
rect 5448 22448 5500 22500
rect 6000 22516 6052 22568
rect 7380 22516 7432 22568
rect 7748 22559 7800 22568
rect 7748 22525 7757 22559
rect 7757 22525 7791 22559
rect 7791 22525 7800 22559
rect 7748 22516 7800 22525
rect 10140 22652 10192 22704
rect 10692 22652 10744 22704
rect 9680 22584 9732 22636
rect 10876 22584 10928 22636
rect 12532 22584 12584 22636
rect 13360 22652 13412 22704
rect 13636 22695 13688 22704
rect 13636 22661 13645 22695
rect 13645 22661 13679 22695
rect 13679 22661 13688 22695
rect 13636 22652 13688 22661
rect 14188 22652 14240 22704
rect 16580 22652 16632 22704
rect 17500 22652 17552 22704
rect 14464 22584 14516 22636
rect 15660 22584 15712 22636
rect 7196 22491 7248 22500
rect 7196 22457 7205 22491
rect 7205 22457 7239 22491
rect 7239 22457 7248 22491
rect 7196 22448 7248 22457
rect 13360 22516 13412 22568
rect 13820 22516 13872 22568
rect 16028 22584 16080 22636
rect 16396 22584 16448 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17776 22584 17828 22636
rect 18052 22652 18104 22704
rect 18696 22695 18748 22704
rect 18696 22661 18705 22695
rect 18705 22661 18739 22695
rect 18739 22661 18748 22695
rect 18696 22652 18748 22661
rect 18236 22584 18288 22636
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 6736 22380 6788 22432
rect 7104 22380 7156 22432
rect 10692 22448 10744 22500
rect 17408 22516 17460 22568
rect 19340 22720 19392 22772
rect 20628 22720 20680 22772
rect 22560 22720 22612 22772
rect 22836 22720 22888 22772
rect 23112 22720 23164 22772
rect 19156 22584 19208 22636
rect 17592 22448 17644 22500
rect 9956 22380 10008 22432
rect 12532 22423 12584 22432
rect 12532 22389 12541 22423
rect 12541 22389 12575 22423
rect 12575 22389 12584 22423
rect 12532 22380 12584 22389
rect 13912 22380 13964 22432
rect 15016 22423 15068 22432
rect 15016 22389 15025 22423
rect 15025 22389 15059 22423
rect 15059 22389 15068 22423
rect 15016 22380 15068 22389
rect 15660 22380 15712 22432
rect 18512 22448 18564 22500
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 18144 22380 18196 22432
rect 19156 22448 19208 22500
rect 19616 22652 19668 22704
rect 20444 22652 20496 22704
rect 20536 22695 20588 22704
rect 20536 22661 20545 22695
rect 20545 22661 20579 22695
rect 20579 22661 20588 22695
rect 20536 22652 20588 22661
rect 21640 22652 21692 22704
rect 23572 22652 23624 22704
rect 19708 22584 19760 22636
rect 20720 22584 20772 22636
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22560 22584 22612 22636
rect 24584 22627 24636 22636
rect 24584 22593 24593 22627
rect 24593 22593 24627 22627
rect 24627 22593 24636 22627
rect 24584 22584 24636 22593
rect 25136 22584 25188 22636
rect 22744 22559 22796 22568
rect 22744 22525 22753 22559
rect 22753 22525 22787 22559
rect 22787 22525 22796 22559
rect 22744 22516 22796 22525
rect 24860 22516 24912 22568
rect 25964 22584 26016 22636
rect 19064 22380 19116 22432
rect 22376 22380 22428 22432
rect 24676 22491 24728 22500
rect 24676 22457 24685 22491
rect 24685 22457 24719 22491
rect 24719 22457 24728 22491
rect 24676 22448 24728 22457
rect 23388 22380 23440 22432
rect 24308 22380 24360 22432
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 2872 22176 2924 22228
rect 3700 22176 3752 22228
rect 4712 22176 4764 22228
rect 5080 22176 5132 22228
rect 5356 22176 5408 22228
rect 6920 22176 6972 22228
rect 7656 22176 7708 22228
rect 8392 22176 8444 22228
rect 1492 22040 1544 22092
rect 1768 22015 1820 22024
rect 1768 21981 1777 22015
rect 1777 21981 1811 22015
rect 1811 21981 1820 22015
rect 1768 21972 1820 21981
rect 1860 21972 1912 22024
rect 2136 22015 2188 22024
rect 2136 21981 2145 22015
rect 2145 21981 2179 22015
rect 2179 21981 2188 22015
rect 2136 21972 2188 21981
rect 572 21904 624 21956
rect 2688 22015 2740 22024
rect 2688 21981 2698 22015
rect 2698 21981 2732 22015
rect 2732 21981 2740 22015
rect 2688 21972 2740 21981
rect 7380 22108 7432 22160
rect 10784 22176 10836 22228
rect 11336 22176 11388 22228
rect 13084 22176 13136 22228
rect 17224 22176 17276 22228
rect 17592 22219 17644 22228
rect 17592 22185 17601 22219
rect 17601 22185 17635 22219
rect 17635 22185 17644 22219
rect 17592 22176 17644 22185
rect 3792 22040 3844 22092
rect 5356 22040 5408 22092
rect 5908 22040 5960 22092
rect 6920 22040 6972 22092
rect 4804 21972 4856 22024
rect 5080 21972 5132 22024
rect 3240 21904 3292 21956
rect 4344 21904 4396 21956
rect 4896 21904 4948 21956
rect 2228 21836 2280 21888
rect 3056 21836 3108 21888
rect 5356 21879 5408 21888
rect 5356 21845 5365 21879
rect 5365 21845 5399 21879
rect 5399 21845 5408 21879
rect 5356 21836 5408 21845
rect 5540 21836 5592 21888
rect 5816 22015 5868 22024
rect 5816 21981 5825 22015
rect 5825 21981 5859 22015
rect 5859 21981 5868 22015
rect 5816 21972 5868 21981
rect 7104 21972 7156 22024
rect 8392 21972 8444 22024
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 6460 21904 6512 21956
rect 6644 21904 6696 21956
rect 10324 22108 10376 22160
rect 10968 22108 11020 22160
rect 14740 22151 14792 22160
rect 14740 22117 14749 22151
rect 14749 22117 14783 22151
rect 14783 22117 14792 22151
rect 14740 22108 14792 22117
rect 15108 22108 15160 22160
rect 18144 22176 18196 22228
rect 18604 22176 18656 22228
rect 18972 22176 19024 22228
rect 19432 22219 19484 22228
rect 19432 22185 19441 22219
rect 19441 22185 19475 22219
rect 19475 22185 19484 22219
rect 19432 22176 19484 22185
rect 19524 22176 19576 22228
rect 19708 22176 19760 22228
rect 24860 22176 24912 22228
rect 25136 22176 25188 22228
rect 21640 22108 21692 22160
rect 8852 22040 8904 22092
rect 13268 22040 13320 22092
rect 16028 22040 16080 22092
rect 9864 21972 9916 22024
rect 10140 21972 10192 22024
rect 9772 21904 9824 21956
rect 10968 21972 11020 22024
rect 12164 21904 12216 21956
rect 12992 21972 13044 22024
rect 13544 21972 13596 22024
rect 14648 21972 14700 22024
rect 18972 22040 19024 22092
rect 20812 22040 20864 22092
rect 21088 22083 21140 22092
rect 21088 22049 21097 22083
rect 21097 22049 21131 22083
rect 21131 22049 21140 22083
rect 21088 22040 21140 22049
rect 12808 21904 12860 21956
rect 15752 21904 15804 21956
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 17132 21904 17184 21956
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 19340 21972 19392 22024
rect 19708 21972 19760 22024
rect 18604 21904 18656 21956
rect 22652 22015 22704 22024
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 24124 22040 24176 22092
rect 6552 21836 6604 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9496 21836 9548 21888
rect 13360 21879 13412 21888
rect 13360 21845 13385 21879
rect 13385 21845 13412 21879
rect 13360 21836 13412 21845
rect 13820 21836 13872 21888
rect 14648 21836 14700 21888
rect 15108 21836 15160 21888
rect 15200 21836 15252 21888
rect 16028 21836 16080 21888
rect 16764 21879 16816 21888
rect 16764 21845 16773 21879
rect 16773 21845 16807 21879
rect 16807 21845 16816 21879
rect 16764 21836 16816 21845
rect 17408 21879 17460 21888
rect 17408 21845 17433 21879
rect 17433 21845 17460 21879
rect 17408 21836 17460 21845
rect 18328 21836 18380 21888
rect 20444 21904 20496 21956
rect 20904 21947 20956 21956
rect 20904 21913 20913 21947
rect 20913 21913 20947 21947
rect 20947 21913 20956 21947
rect 20904 21904 20956 21913
rect 21456 21904 21508 21956
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 23756 21836 23808 21888
rect 23848 21836 23900 21888
rect 24676 21836 24728 21888
rect 28172 21879 28224 21888
rect 28172 21845 28181 21879
rect 28181 21845 28215 21879
rect 28215 21845 28224 21879
rect 28172 21836 28224 21845
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 3608 21632 3660 21684
rect 5264 21632 5316 21684
rect 6276 21632 6328 21684
rect 7656 21632 7708 21684
rect 1768 21564 1820 21616
rect 4896 21564 4948 21616
rect 6644 21564 6696 21616
rect 6736 21564 6788 21616
rect 2228 21539 2280 21548
rect 2228 21505 2237 21539
rect 2237 21505 2271 21539
rect 2271 21505 2280 21539
rect 2228 21496 2280 21505
rect 2504 21539 2556 21548
rect 2504 21505 2513 21539
rect 2513 21505 2547 21539
rect 2547 21505 2556 21539
rect 2504 21496 2556 21505
rect 3056 21539 3108 21548
rect 3056 21505 3065 21539
rect 3065 21505 3099 21539
rect 3099 21505 3108 21539
rect 3056 21496 3108 21505
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 5172 21496 5224 21548
rect 480 21428 532 21480
rect 1768 21428 1820 21480
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 5816 21496 5868 21548
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7104 21539 7156 21548
rect 7104 21505 7113 21539
rect 7113 21505 7147 21539
rect 7147 21505 7156 21539
rect 7104 21496 7156 21505
rect 7748 21496 7800 21548
rect 8760 21496 8812 21548
rect 9956 21632 10008 21684
rect 10692 21632 10744 21684
rect 10784 21632 10836 21684
rect 11060 21564 11112 21616
rect 11152 21564 11204 21616
rect 12716 21675 12768 21684
rect 12716 21641 12725 21675
rect 12725 21641 12759 21675
rect 12759 21641 12768 21675
rect 12716 21632 12768 21641
rect 12900 21632 12952 21684
rect 15844 21675 15896 21684
rect 15844 21641 15853 21675
rect 15853 21641 15887 21675
rect 15887 21641 15896 21675
rect 15844 21632 15896 21641
rect 16212 21632 16264 21684
rect 14280 21564 14332 21616
rect 15752 21564 15804 21616
rect 16948 21564 17000 21616
rect 17224 21564 17276 21616
rect 18420 21632 18472 21684
rect 19708 21675 19760 21684
rect 19708 21641 19717 21675
rect 19717 21641 19751 21675
rect 19751 21641 19760 21675
rect 19708 21632 19760 21641
rect 22192 21632 22244 21684
rect 22284 21632 22336 21684
rect 26240 21632 26292 21684
rect 18144 21564 18196 21616
rect 10692 21496 10744 21548
rect 10784 21496 10836 21548
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 11796 21496 11848 21548
rect 12440 21496 12492 21548
rect 12624 21496 12676 21548
rect 5540 21428 5592 21480
rect 12992 21496 13044 21548
rect 16488 21496 16540 21548
rect 17316 21496 17368 21548
rect 19892 21564 19944 21616
rect 23940 21607 23992 21616
rect 23940 21573 23974 21607
rect 23974 21573 23992 21607
rect 23940 21564 23992 21573
rect 24032 21564 24084 21616
rect 25044 21564 25096 21616
rect 20352 21496 20404 21548
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 21272 21539 21324 21548
rect 21272 21505 21281 21539
rect 21281 21505 21315 21539
rect 21315 21505 21324 21539
rect 21272 21496 21324 21505
rect 21732 21496 21784 21548
rect 23296 21496 23348 21548
rect 1952 21360 2004 21412
rect 9404 21403 9456 21412
rect 9404 21369 9413 21403
rect 9413 21369 9447 21403
rect 9447 21369 9456 21403
rect 9404 21360 9456 21369
rect 9680 21360 9732 21412
rect 9956 21360 10008 21412
rect 1676 21292 1728 21344
rect 6092 21292 6144 21344
rect 6920 21292 6972 21344
rect 8300 21292 8352 21344
rect 8944 21292 8996 21344
rect 9496 21292 9548 21344
rect 10232 21335 10284 21344
rect 10232 21301 10241 21335
rect 10241 21301 10275 21335
rect 10275 21301 10284 21335
rect 10232 21292 10284 21301
rect 10692 21292 10744 21344
rect 10968 21292 11020 21344
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 12072 21292 12124 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 13728 21292 13780 21344
rect 15200 21335 15252 21344
rect 15200 21301 15209 21335
rect 15209 21301 15243 21335
rect 15243 21301 15252 21335
rect 15200 21292 15252 21301
rect 17040 21335 17092 21344
rect 17040 21301 17049 21335
rect 17049 21301 17083 21335
rect 17083 21301 17092 21335
rect 17040 21292 17092 21301
rect 20996 21428 21048 21480
rect 22100 21428 22152 21480
rect 19156 21360 19208 21412
rect 22284 21403 22336 21412
rect 22284 21369 22293 21403
rect 22293 21369 22327 21403
rect 22327 21369 22336 21403
rect 22284 21360 22336 21369
rect 22652 21428 22704 21480
rect 23480 21360 23532 21412
rect 18788 21292 18840 21344
rect 20444 21292 20496 21344
rect 22836 21292 22888 21344
rect 23112 21292 23164 21344
rect 25596 21360 25648 21412
rect 25044 21335 25096 21344
rect 25044 21301 25053 21335
rect 25053 21301 25087 21335
rect 25087 21301 25096 21335
rect 25044 21292 25096 21301
rect 25136 21292 25188 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 2596 21088 2648 21140
rect 3424 21131 3476 21140
rect 3424 21097 3433 21131
rect 3433 21097 3467 21131
rect 3467 21097 3476 21131
rect 3424 21088 3476 21097
rect 2044 21020 2096 21072
rect 3240 21020 3292 21072
rect 4160 21020 4212 21072
rect 5264 21020 5316 21072
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 7012 21088 7064 21140
rect 7564 21088 7616 21140
rect 10048 21088 10100 21140
rect 12992 21088 13044 21140
rect 13084 21088 13136 21140
rect 13636 21088 13688 21140
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 15292 21088 15344 21140
rect 15660 21088 15712 21140
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 17960 21088 18012 21140
rect 18880 21088 18932 21140
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 5540 21020 5592 21072
rect 6552 21063 6604 21072
rect 6552 21029 6561 21063
rect 6561 21029 6595 21063
rect 6595 21029 6604 21063
rect 6552 21020 6604 21029
rect 9496 21020 9548 21072
rect 9680 21020 9732 21072
rect 12624 21063 12676 21072
rect 12624 21029 12633 21063
rect 12633 21029 12667 21063
rect 12667 21029 12676 21063
rect 12624 21020 12676 21029
rect 12808 21020 12860 21072
rect 1676 20927 1728 20936
rect 1676 20893 1686 20927
rect 1686 20893 1720 20927
rect 1720 20893 1728 20927
rect 3056 20952 3108 21004
rect 1676 20884 1728 20893
rect 2044 20927 2096 20936
rect 2044 20893 2058 20927
rect 2058 20893 2092 20927
rect 2092 20893 2096 20927
rect 2044 20884 2096 20893
rect 2228 20816 2280 20868
rect 3240 20927 3292 20936
rect 3240 20893 3254 20927
rect 3254 20893 3288 20927
rect 3288 20893 3292 20927
rect 3240 20884 3292 20893
rect 3516 20884 3568 20936
rect 6644 20995 6696 21004
rect 6644 20961 6653 20995
rect 6653 20961 6687 20995
rect 6687 20961 6696 20995
rect 6644 20952 6696 20961
rect 9312 20952 9364 21004
rect 10324 20952 10376 21004
rect 10784 20952 10836 21004
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 5080 20884 5132 20936
rect 5264 20927 5316 20936
rect 5264 20893 5273 20927
rect 5273 20893 5307 20927
rect 5307 20893 5316 20927
rect 5264 20884 5316 20893
rect 5448 20884 5500 20936
rect 2320 20748 2372 20800
rect 2872 20748 2924 20800
rect 3700 20816 3752 20868
rect 8392 20884 8444 20936
rect 8576 20927 8628 20936
rect 8576 20893 8585 20927
rect 8585 20893 8619 20927
rect 8619 20893 8628 20927
rect 8576 20884 8628 20893
rect 9680 20884 9732 20936
rect 13912 20952 13964 21004
rect 17776 21020 17828 21072
rect 23112 21063 23164 21072
rect 23112 21029 23121 21063
rect 23121 21029 23155 21063
rect 23155 21029 23164 21063
rect 23112 21020 23164 21029
rect 23296 21131 23348 21140
rect 23296 21097 23305 21131
rect 23305 21097 23339 21131
rect 23339 21097 23348 21131
rect 23296 21088 23348 21097
rect 23572 21020 23624 21072
rect 8300 20816 8352 20868
rect 8668 20816 8720 20868
rect 9312 20816 9364 20868
rect 11428 20859 11480 20868
rect 11428 20825 11437 20859
rect 11437 20825 11471 20859
rect 11471 20825 11480 20859
rect 11428 20816 11480 20825
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 13360 20884 13412 20936
rect 13176 20816 13228 20868
rect 4068 20748 4120 20800
rect 4344 20748 4396 20800
rect 9588 20748 9640 20800
rect 10048 20791 10100 20800
rect 10048 20757 10057 20791
rect 10057 20757 10091 20791
rect 10091 20757 10100 20791
rect 10048 20748 10100 20757
rect 10784 20748 10836 20800
rect 14004 20816 14056 20868
rect 15752 20884 15804 20936
rect 17040 20884 17092 20936
rect 17868 20884 17920 20936
rect 13912 20748 13964 20800
rect 15108 20816 15160 20868
rect 15936 20816 15988 20868
rect 16028 20816 16080 20868
rect 17500 20816 17552 20868
rect 17684 20816 17736 20868
rect 18328 20816 18380 20868
rect 16304 20748 16356 20800
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 17960 20748 18012 20800
rect 19248 20884 19300 20936
rect 19708 20952 19760 21004
rect 24400 20952 24452 21004
rect 19616 20927 19668 20936
rect 19616 20893 19623 20927
rect 19623 20893 19668 20927
rect 19616 20884 19668 20893
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 19892 20927 19944 20936
rect 19892 20893 19906 20927
rect 19906 20893 19940 20927
rect 19940 20893 19944 20927
rect 19892 20884 19944 20893
rect 19156 20816 19208 20868
rect 20444 20816 20496 20868
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 20812 20816 20864 20868
rect 21548 20859 21600 20868
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 22100 20816 22152 20868
rect 23020 20816 23072 20868
rect 19616 20748 19668 20800
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 27804 21088 27856 21140
rect 24584 20995 24636 21004
rect 24584 20961 24593 20995
rect 24593 20961 24627 20995
rect 24627 20961 24636 20995
rect 24584 20952 24636 20961
rect 25136 20884 25188 20936
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 24952 20816 25004 20868
rect 25872 20748 25924 20800
rect 26332 20748 26384 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 1308 20544 1360 20596
rect 2412 20544 2464 20596
rect 2872 20476 2924 20528
rect 1676 20408 1728 20460
rect 2136 20408 2188 20460
rect 3516 20544 3568 20596
rect 1124 20340 1176 20392
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 3516 20408 3568 20460
rect 4252 20476 4304 20528
rect 4712 20519 4764 20528
rect 4712 20485 4721 20519
rect 4721 20485 4755 20519
rect 4755 20485 4764 20519
rect 4712 20476 4764 20485
rect 4988 20587 5040 20596
rect 4988 20553 4997 20587
rect 4997 20553 5031 20587
rect 5031 20553 5040 20587
rect 4988 20544 5040 20553
rect 5080 20544 5132 20596
rect 5908 20476 5960 20528
rect 4436 20451 4488 20460
rect 4436 20417 4445 20451
rect 4445 20417 4479 20451
rect 4479 20417 4488 20451
rect 4436 20408 4488 20417
rect 4988 20408 5040 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 6736 20476 6788 20528
rect 7380 20408 7432 20460
rect 7564 20408 7616 20460
rect 10232 20476 10284 20528
rect 9864 20408 9916 20460
rect 4160 20340 4212 20392
rect 5448 20383 5500 20392
rect 5448 20349 5457 20383
rect 5457 20349 5491 20383
rect 5491 20349 5500 20383
rect 5448 20340 5500 20349
rect 1492 20204 1544 20256
rect 4804 20272 4856 20324
rect 8852 20383 8904 20392
rect 8852 20349 8861 20383
rect 8861 20349 8895 20383
rect 8895 20349 8904 20383
rect 8852 20340 8904 20349
rect 6092 20272 6144 20324
rect 9772 20272 9824 20324
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 11888 20476 11940 20528
rect 11152 20408 11204 20460
rect 13544 20544 13596 20596
rect 14464 20544 14516 20596
rect 18236 20544 18288 20596
rect 13452 20476 13504 20528
rect 20076 20544 20128 20596
rect 24216 20544 24268 20596
rect 25688 20544 25740 20596
rect 13268 20408 13320 20460
rect 14832 20408 14884 20460
rect 16488 20408 16540 20460
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17500 20408 17552 20460
rect 17868 20451 17920 20460
rect 17868 20417 17877 20451
rect 17877 20417 17911 20451
rect 17911 20417 17920 20451
rect 17868 20408 17920 20417
rect 18880 20451 18932 20460
rect 18880 20417 18889 20451
rect 18889 20417 18923 20451
rect 18923 20417 18932 20451
rect 18880 20408 18932 20417
rect 21548 20476 21600 20528
rect 21732 20476 21784 20528
rect 24768 20476 24820 20528
rect 19156 20451 19208 20460
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 11060 20340 11112 20392
rect 12440 20340 12492 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 15292 20340 15344 20392
rect 15752 20340 15804 20392
rect 17592 20340 17644 20392
rect 17960 20340 18012 20392
rect 19892 20408 19944 20460
rect 20444 20451 20496 20460
rect 20444 20417 20453 20451
rect 20453 20417 20487 20451
rect 20487 20417 20496 20451
rect 20444 20408 20496 20417
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 19524 20340 19576 20392
rect 19800 20340 19852 20392
rect 19984 20340 20036 20392
rect 22744 20408 22796 20460
rect 24584 20408 24636 20460
rect 25136 20408 25188 20460
rect 26240 20408 26292 20460
rect 10692 20272 10744 20324
rect 10784 20272 10836 20324
rect 3148 20204 3200 20256
rect 3792 20247 3844 20256
rect 3792 20213 3801 20247
rect 3801 20213 3835 20247
rect 3835 20213 3844 20247
rect 3792 20204 3844 20213
rect 4712 20204 4764 20256
rect 5540 20204 5592 20256
rect 6276 20204 6328 20256
rect 7380 20204 7432 20256
rect 7840 20204 7892 20256
rect 8852 20204 8904 20256
rect 10232 20204 10284 20256
rect 14004 20204 14056 20256
rect 14188 20204 14240 20256
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 16028 20204 16080 20256
rect 19892 20272 19944 20324
rect 20628 20272 20680 20324
rect 21732 20272 21784 20324
rect 19524 20247 19576 20256
rect 19524 20213 19533 20247
rect 19533 20213 19567 20247
rect 19567 20213 19576 20247
rect 19524 20204 19576 20213
rect 22836 20204 22888 20256
rect 23572 20247 23624 20256
rect 23572 20213 23581 20247
rect 23581 20213 23615 20247
rect 23615 20213 23624 20247
rect 23572 20204 23624 20213
rect 26516 20204 26568 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 3976 20000 4028 20052
rect 4896 20000 4948 20052
rect 7840 20000 7892 20052
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 8392 20000 8444 20052
rect 2596 19932 2648 19984
rect 5448 19932 5500 19984
rect 5172 19907 5224 19916
rect 5172 19873 5181 19907
rect 5181 19873 5215 19907
rect 5215 19873 5224 19907
rect 5172 19864 5224 19873
rect 5632 19864 5684 19916
rect 1952 19839 2004 19848
rect 1952 19805 1961 19839
rect 1961 19805 1995 19839
rect 1995 19805 2004 19839
rect 1952 19796 2004 19805
rect 1860 19728 1912 19780
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 2872 19796 2924 19805
rect 3332 19796 3384 19848
rect 3608 19796 3660 19848
rect 3976 19796 4028 19848
rect 4160 19796 4212 19848
rect 4712 19796 4764 19848
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 5908 19796 5960 19848
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 11704 20000 11756 20052
rect 11980 20000 12032 20052
rect 12532 20000 12584 20052
rect 13084 20000 13136 20052
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 12624 19932 12676 19984
rect 12900 19932 12952 19984
rect 15476 20000 15528 20052
rect 16212 20000 16264 20052
rect 17776 20000 17828 20052
rect 17868 20000 17920 20052
rect 18972 20000 19024 20052
rect 16672 19932 16724 19984
rect 18052 19932 18104 19984
rect 19432 19932 19484 19984
rect 20720 20000 20772 20052
rect 21272 20000 21324 20052
rect 24952 20000 25004 20052
rect 22192 19932 22244 19984
rect 26424 19932 26476 19984
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 11336 19864 11388 19916
rect 11888 19864 11940 19916
rect 12348 19864 12400 19916
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 848 19660 900 19712
rect 2228 19660 2280 19712
rect 2780 19728 2832 19780
rect 4804 19728 4856 19780
rect 6184 19728 6236 19780
rect 9220 19796 9272 19848
rect 8668 19728 8720 19780
rect 12532 19796 12584 19848
rect 12624 19796 12676 19848
rect 13176 19796 13228 19848
rect 13452 19796 13504 19848
rect 19524 19864 19576 19916
rect 21088 19864 21140 19916
rect 23572 19864 23624 19916
rect 26792 19864 26844 19916
rect 14372 19796 14424 19848
rect 14924 19796 14976 19848
rect 15384 19796 15436 19848
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 15936 19796 15988 19848
rect 16304 19796 16356 19848
rect 17408 19796 17460 19848
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17500 19796 17552 19805
rect 5632 19703 5684 19712
rect 5632 19669 5641 19703
rect 5641 19669 5675 19703
rect 5675 19669 5684 19703
rect 5632 19660 5684 19669
rect 9496 19660 9548 19712
rect 11244 19728 11296 19780
rect 14280 19728 14332 19780
rect 11796 19660 11848 19712
rect 12072 19703 12124 19712
rect 12072 19669 12097 19703
rect 12097 19669 12124 19703
rect 12072 19660 12124 19669
rect 12992 19660 13044 19712
rect 14464 19660 14516 19712
rect 15660 19728 15712 19780
rect 15752 19728 15804 19780
rect 17316 19728 17368 19780
rect 14924 19703 14976 19712
rect 14924 19669 14949 19703
rect 14949 19669 14976 19703
rect 14924 19660 14976 19669
rect 15108 19703 15160 19712
rect 15108 19669 15117 19703
rect 15117 19669 15151 19703
rect 15151 19669 15160 19703
rect 15108 19660 15160 19669
rect 19800 19796 19852 19848
rect 20720 19796 20772 19848
rect 22284 19796 22336 19848
rect 19524 19728 19576 19780
rect 20444 19728 20496 19780
rect 21180 19728 21232 19780
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 24216 19728 24268 19780
rect 21548 19660 21600 19712
rect 22560 19660 22612 19712
rect 26056 19660 26108 19712
rect 28356 19703 28408 19712
rect 28356 19669 28365 19703
rect 28365 19669 28399 19703
rect 28399 19669 28408 19703
rect 28356 19660 28408 19669
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 2504 19456 2556 19508
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 3148 19456 3200 19508
rect 3240 19456 3292 19508
rect 4436 19456 4488 19508
rect 4804 19456 4856 19508
rect 5172 19456 5224 19508
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 10784 19456 10836 19508
rect 11244 19456 11296 19508
rect 14464 19456 14516 19508
rect 14556 19456 14608 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 16672 19456 16724 19508
rect 17960 19456 18012 19508
rect 22376 19456 22428 19508
rect 22744 19456 22796 19508
rect 23388 19499 23440 19508
rect 23388 19465 23397 19499
rect 23397 19465 23431 19499
rect 23431 19465 23440 19499
rect 23388 19456 23440 19465
rect 3792 19388 3844 19440
rect 3976 19388 4028 19440
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 2688 19320 2740 19372
rect 4160 19320 4212 19372
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2596 19252 2648 19304
rect 2044 19184 2096 19236
rect 5080 19388 5132 19440
rect 6092 19388 6144 19440
rect 7380 19388 7432 19440
rect 9772 19388 9824 19440
rect 4988 19363 5040 19372
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 5448 19320 5500 19372
rect 5540 19320 5592 19372
rect 6184 19320 6236 19372
rect 7472 19320 7524 19372
rect 7656 19320 7708 19372
rect 8944 19363 8996 19372
rect 8944 19329 8953 19363
rect 8953 19329 8987 19363
rect 8987 19329 8996 19363
rect 8944 19320 8996 19329
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 9404 19320 9456 19372
rect 10692 19363 10744 19372
rect 6552 19252 6604 19304
rect 10324 19252 10376 19304
rect 2964 19116 3016 19168
rect 3608 19116 3660 19168
rect 3700 19116 3752 19168
rect 5080 19116 5132 19168
rect 7472 19184 7524 19236
rect 5540 19116 5592 19168
rect 6092 19116 6144 19168
rect 8208 19116 8260 19168
rect 9404 19184 9456 19236
rect 10692 19329 10701 19363
rect 10701 19329 10735 19363
rect 10735 19329 10744 19363
rect 10692 19320 10744 19329
rect 10784 19295 10836 19304
rect 10784 19261 10793 19295
rect 10793 19261 10827 19295
rect 10827 19261 10836 19295
rect 10784 19252 10836 19261
rect 11612 19320 11664 19372
rect 13176 19388 13228 19440
rect 13268 19431 13320 19440
rect 13268 19397 13293 19431
rect 13293 19397 13320 19431
rect 13268 19388 13320 19397
rect 13544 19388 13596 19440
rect 13912 19431 13964 19440
rect 13912 19397 13921 19431
rect 13921 19397 13955 19431
rect 13955 19397 13964 19431
rect 13912 19388 13964 19397
rect 14004 19388 14056 19440
rect 14648 19388 14700 19440
rect 14832 19388 14884 19440
rect 15476 19388 15528 19440
rect 16396 19388 16448 19440
rect 17132 19388 17184 19440
rect 17868 19388 17920 19440
rect 18144 19388 18196 19440
rect 18972 19388 19024 19440
rect 19892 19431 19944 19440
rect 19892 19397 19901 19431
rect 19901 19397 19935 19431
rect 19935 19397 19944 19431
rect 19892 19388 19944 19397
rect 21456 19388 21508 19440
rect 23020 19388 23072 19440
rect 23756 19388 23808 19440
rect 15660 19320 15712 19372
rect 11152 19252 11204 19304
rect 11244 19252 11296 19304
rect 12348 19295 12400 19304
rect 12348 19261 12382 19295
rect 12382 19261 12400 19295
rect 16212 19320 16264 19372
rect 17592 19320 17644 19372
rect 17776 19320 17828 19372
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 12348 19252 12400 19261
rect 12900 19184 12952 19236
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 18144 19252 18196 19304
rect 18604 19320 18656 19372
rect 21088 19320 21140 19372
rect 19340 19252 19392 19304
rect 20628 19252 20680 19304
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 21272 19252 21324 19304
rect 26792 19388 26844 19440
rect 24308 19363 24360 19372
rect 24308 19329 24331 19363
rect 24331 19329 24360 19363
rect 24308 19320 24360 19329
rect 20168 19227 20220 19236
rect 20168 19193 20177 19227
rect 20177 19193 20211 19227
rect 20211 19193 20220 19227
rect 20168 19184 20220 19193
rect 9496 19116 9548 19168
rect 10692 19116 10744 19168
rect 11336 19116 11388 19168
rect 13268 19159 13320 19168
rect 13268 19125 13277 19159
rect 13277 19125 13311 19159
rect 13311 19125 13320 19159
rect 13268 19116 13320 19125
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 14096 19159 14148 19168
rect 14096 19125 14105 19159
rect 14105 19125 14139 19159
rect 14139 19125 14148 19159
rect 14096 19116 14148 19125
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 15844 19159 15896 19168
rect 15844 19125 15853 19159
rect 15853 19125 15887 19159
rect 15887 19125 15896 19159
rect 15844 19116 15896 19125
rect 17500 19116 17552 19168
rect 18052 19116 18104 19168
rect 18604 19116 18656 19168
rect 20904 19116 20956 19168
rect 20996 19116 21048 19168
rect 23296 19227 23348 19236
rect 23296 19193 23305 19227
rect 23305 19193 23339 19227
rect 23339 19193 23348 19227
rect 23296 19184 23348 19193
rect 23572 19184 23624 19236
rect 23848 19116 23900 19168
rect 28172 19184 28224 19236
rect 25044 19116 25096 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 4160 18912 4212 18964
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 2228 18776 2280 18828
rect 1860 18572 1912 18624
rect 2596 18708 2648 18760
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 4252 18844 4304 18896
rect 4344 18887 4396 18896
rect 4344 18853 4353 18887
rect 4353 18853 4387 18887
rect 4387 18853 4396 18887
rect 4344 18844 4396 18853
rect 4436 18844 4488 18896
rect 4988 18844 5040 18896
rect 7472 18912 7524 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 10324 18912 10376 18964
rect 13820 18912 13872 18964
rect 16764 18912 16816 18964
rect 19248 18912 19300 18964
rect 21180 18912 21232 18964
rect 21640 18955 21692 18964
rect 21640 18921 21649 18955
rect 21649 18921 21683 18955
rect 21683 18921 21692 18955
rect 21640 18912 21692 18921
rect 6828 18844 6880 18896
rect 7840 18844 7892 18896
rect 8852 18844 8904 18896
rect 11612 18844 11664 18896
rect 11980 18844 12032 18896
rect 16212 18844 16264 18896
rect 16856 18844 16908 18896
rect 18604 18844 18656 18896
rect 24952 18912 25004 18964
rect 4160 18776 4212 18828
rect 6736 18776 6788 18828
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3792 18708 3844 18760
rect 4252 18708 4304 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4896 18708 4948 18760
rect 2780 18640 2832 18692
rect 6184 18708 6236 18760
rect 6644 18708 6696 18760
rect 7472 18708 7524 18760
rect 5632 18640 5684 18692
rect 6092 18640 6144 18692
rect 7196 18640 7248 18692
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 9220 18708 9272 18760
rect 9864 18776 9916 18828
rect 10600 18776 10652 18828
rect 11060 18776 11112 18828
rect 10508 18708 10560 18760
rect 11520 18776 11572 18828
rect 11888 18776 11940 18828
rect 12256 18776 12308 18828
rect 23296 18844 23348 18896
rect 8944 18640 8996 18692
rect 2872 18572 2924 18624
rect 5264 18572 5316 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 6184 18572 6236 18624
rect 7748 18572 7800 18624
rect 10784 18640 10836 18692
rect 11612 18708 11664 18760
rect 14004 18708 14056 18760
rect 12348 18640 12400 18692
rect 12992 18640 13044 18692
rect 10140 18572 10192 18624
rect 10692 18572 10744 18624
rect 11152 18572 11204 18624
rect 11428 18572 11480 18624
rect 12808 18572 12860 18624
rect 13084 18615 13136 18624
rect 14280 18640 14332 18692
rect 14464 18640 14516 18692
rect 15384 18708 15436 18760
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 17868 18708 17920 18760
rect 18052 18708 18104 18760
rect 20720 18776 20772 18828
rect 19340 18708 19392 18760
rect 15200 18640 15252 18692
rect 19892 18751 19944 18760
rect 19892 18717 19901 18751
rect 19901 18717 19935 18751
rect 19935 18717 19944 18751
rect 19892 18708 19944 18717
rect 20168 18751 20220 18760
rect 20168 18717 20177 18751
rect 20177 18717 20211 18751
rect 20211 18717 20220 18751
rect 20168 18708 20220 18717
rect 20352 18708 20404 18760
rect 20904 18708 20956 18760
rect 21364 18708 21416 18760
rect 13084 18581 13109 18615
rect 13109 18581 13136 18615
rect 13084 18572 13136 18581
rect 13636 18572 13688 18624
rect 15292 18572 15344 18624
rect 17132 18572 17184 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 20260 18640 20312 18692
rect 21180 18640 21232 18692
rect 18696 18572 18748 18624
rect 19432 18615 19484 18624
rect 19432 18581 19441 18615
rect 19441 18581 19475 18615
rect 19475 18581 19484 18615
rect 19432 18572 19484 18581
rect 20812 18572 20864 18624
rect 21364 18572 21416 18624
rect 21916 18640 21968 18692
rect 24400 18776 24452 18828
rect 25136 18776 25188 18828
rect 22836 18708 22888 18760
rect 23480 18708 23532 18760
rect 22560 18683 22612 18692
rect 22100 18572 22152 18624
rect 22560 18649 22572 18683
rect 22572 18649 22612 18683
rect 22560 18640 22612 18649
rect 23572 18572 23624 18624
rect 23664 18615 23716 18624
rect 23664 18581 23673 18615
rect 23673 18581 23707 18615
rect 23707 18581 23716 18615
rect 23664 18572 23716 18581
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 2136 18411 2188 18420
rect 2136 18377 2145 18411
rect 2145 18377 2179 18411
rect 2179 18377 2188 18411
rect 2136 18368 2188 18377
rect 4528 18368 4580 18420
rect 3700 18300 3752 18352
rect 4988 18368 5040 18420
rect 5356 18368 5408 18420
rect 2412 18232 2464 18284
rect 2688 18275 2740 18284
rect 2688 18241 2697 18275
rect 2697 18241 2731 18275
rect 2731 18241 2740 18275
rect 2688 18232 2740 18241
rect 2872 18275 2924 18284
rect 2872 18241 2879 18275
rect 2879 18241 2924 18275
rect 2872 18232 2924 18241
rect 2964 18275 3016 18284
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 4344 18275 4396 18284
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 4528 18275 4580 18284
rect 4528 18241 4535 18275
rect 4535 18241 4580 18275
rect 4528 18232 4580 18241
rect 4896 18232 4948 18284
rect 7196 18368 7248 18420
rect 8116 18368 8168 18420
rect 8576 18368 8628 18420
rect 10600 18368 10652 18420
rect 13636 18368 13688 18420
rect 14832 18368 14884 18420
rect 16948 18368 17000 18420
rect 17040 18368 17092 18420
rect 18328 18368 18380 18420
rect 20628 18368 20680 18420
rect 23664 18368 23716 18420
rect 11980 18300 12032 18352
rect 12256 18343 12308 18352
rect 12256 18309 12265 18343
rect 12265 18309 12299 18343
rect 12299 18309 12308 18343
rect 12256 18300 12308 18309
rect 12348 18343 12400 18352
rect 12348 18309 12357 18343
rect 12357 18309 12391 18343
rect 12391 18309 12400 18343
rect 12348 18300 12400 18309
rect 12440 18343 12492 18352
rect 12440 18309 12449 18343
rect 12449 18309 12483 18343
rect 12483 18309 12492 18343
rect 12440 18300 12492 18309
rect 13360 18300 13412 18352
rect 3608 18164 3660 18216
rect 4620 18164 4672 18216
rect 1308 18028 1360 18080
rect 7288 18232 7340 18284
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 9496 18232 9548 18284
rect 9772 18232 9824 18284
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 11428 18232 11480 18284
rect 12072 18232 12124 18284
rect 13268 18232 13320 18284
rect 7104 18207 7156 18216
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 13544 18232 13596 18284
rect 14188 18232 14240 18284
rect 19432 18300 19484 18352
rect 5908 18096 5960 18148
rect 6368 18096 6420 18148
rect 3148 18028 3200 18080
rect 4068 18028 4120 18080
rect 7748 18028 7800 18080
rect 7840 18028 7892 18080
rect 8852 18028 8904 18080
rect 11612 18164 11664 18216
rect 12900 18164 12952 18216
rect 13360 18164 13412 18216
rect 14096 18164 14148 18216
rect 10692 18028 10744 18080
rect 15016 18096 15068 18148
rect 15384 18164 15436 18216
rect 15660 18232 15712 18284
rect 16396 18232 16448 18284
rect 17500 18232 17552 18284
rect 19340 18232 19392 18284
rect 20168 18300 20220 18352
rect 21456 18300 21508 18352
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 19800 18232 19852 18284
rect 13544 18028 13596 18080
rect 13636 18028 13688 18080
rect 14832 18028 14884 18080
rect 16120 18096 16172 18148
rect 16212 18028 16264 18080
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 18604 18164 18656 18216
rect 20076 18164 20128 18216
rect 20812 18096 20864 18148
rect 19340 18028 19392 18080
rect 22468 18096 22520 18148
rect 23756 18232 23808 18284
rect 24124 18232 24176 18284
rect 23664 18164 23716 18216
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 27436 18164 27488 18216
rect 22560 18028 22612 18080
rect 23940 18096 23992 18148
rect 22744 18028 22796 18080
rect 25044 18028 25096 18080
rect 25780 18071 25832 18080
rect 25780 18037 25789 18071
rect 25789 18037 25823 18071
rect 25823 18037 25832 18071
rect 25780 18028 25832 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 1032 17824 1084 17876
rect 2780 17824 2832 17876
rect 4160 17824 4212 17876
rect 4344 17824 4396 17876
rect 5540 17824 5592 17876
rect 5632 17867 5684 17876
rect 5632 17833 5641 17867
rect 5641 17833 5675 17867
rect 5675 17833 5684 17867
rect 5632 17824 5684 17833
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 3976 17756 4028 17808
rect 2596 17620 2648 17672
rect 1860 17552 1912 17604
rect 2412 17595 2464 17604
rect 2412 17561 2421 17595
rect 2421 17561 2455 17595
rect 2455 17561 2464 17595
rect 2412 17552 2464 17561
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 3424 17731 3476 17740
rect 3424 17697 3433 17731
rect 3433 17697 3467 17731
rect 3467 17697 3476 17731
rect 5724 17756 5776 17808
rect 8300 17824 8352 17876
rect 8392 17824 8444 17876
rect 7012 17756 7064 17808
rect 7840 17756 7892 17808
rect 3424 17688 3476 17697
rect 4344 17688 4396 17740
rect 3424 17552 3476 17604
rect 4896 17620 4948 17672
rect 5172 17620 5224 17672
rect 5632 17620 5684 17672
rect 7472 17688 7524 17740
rect 9864 17756 9916 17808
rect 10508 17756 10560 17808
rect 10692 17756 10744 17808
rect 12808 17867 12860 17876
rect 12808 17833 12817 17867
rect 12817 17833 12851 17867
rect 12851 17833 12860 17867
rect 12808 17824 12860 17833
rect 13636 17824 13688 17876
rect 13820 17824 13872 17876
rect 15384 17824 15436 17876
rect 6736 17663 6788 17672
rect 6736 17629 6745 17663
rect 6745 17629 6779 17663
rect 6779 17629 6788 17663
rect 6736 17620 6788 17629
rect 4068 17552 4120 17604
rect 6552 17552 6604 17604
rect 7196 17552 7248 17604
rect 7748 17620 7800 17672
rect 7840 17663 7892 17672
rect 7840 17629 7849 17663
rect 7849 17629 7883 17663
rect 7883 17629 7892 17663
rect 7840 17620 7892 17629
rect 8484 17620 8536 17672
rect 10324 17688 10376 17740
rect 10416 17688 10468 17740
rect 11428 17688 11480 17740
rect 8300 17552 8352 17604
rect 9680 17620 9732 17672
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 9956 17552 10008 17604
rect 10968 17620 11020 17672
rect 11060 17620 11112 17672
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12256 17620 12308 17672
rect 12532 17688 12584 17740
rect 15200 17688 15252 17740
rect 15660 17799 15712 17808
rect 15660 17765 15669 17799
rect 15669 17765 15703 17799
rect 15703 17765 15712 17799
rect 15660 17756 15712 17765
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 17776 17824 17828 17876
rect 18788 17824 18840 17876
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 16764 17756 16816 17808
rect 19984 17756 20036 17808
rect 20168 17688 20220 17740
rect 22560 17756 22612 17808
rect 23020 17756 23072 17808
rect 23848 17824 23900 17876
rect 26332 17824 26384 17876
rect 24308 17756 24360 17808
rect 23940 17688 23992 17740
rect 26792 17824 26844 17876
rect 27804 17799 27856 17808
rect 27804 17765 27813 17799
rect 27813 17765 27847 17799
rect 27847 17765 27856 17799
rect 27804 17756 27856 17765
rect 13268 17620 13320 17672
rect 11152 17552 11204 17604
rect 11428 17552 11480 17604
rect 4988 17484 5040 17536
rect 5356 17484 5408 17536
rect 6092 17484 6144 17536
rect 8852 17484 8904 17536
rect 9864 17484 9916 17536
rect 11704 17484 11756 17536
rect 12348 17552 12400 17604
rect 13912 17552 13964 17604
rect 15016 17620 15068 17672
rect 15936 17620 15988 17672
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 12808 17484 12860 17536
rect 16028 17552 16080 17604
rect 16304 17552 16356 17604
rect 17132 17595 17184 17604
rect 17132 17561 17141 17595
rect 17141 17561 17175 17595
rect 17175 17561 17184 17595
rect 17132 17552 17184 17561
rect 17592 17552 17644 17604
rect 15384 17484 15436 17536
rect 15660 17484 15712 17536
rect 16396 17527 16448 17536
rect 16396 17493 16421 17527
rect 16421 17493 16448 17527
rect 16396 17484 16448 17493
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 16856 17484 16908 17536
rect 18052 17552 18104 17604
rect 19248 17620 19300 17672
rect 19524 17620 19576 17672
rect 19984 17620 20036 17672
rect 18604 17552 18656 17604
rect 18972 17484 19024 17536
rect 19616 17595 19668 17604
rect 19616 17561 19625 17595
rect 19625 17561 19659 17595
rect 19659 17561 19668 17595
rect 19616 17552 19668 17561
rect 20076 17552 20128 17604
rect 19248 17484 19300 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 22468 17620 22520 17672
rect 21548 17552 21600 17604
rect 22560 17552 22612 17604
rect 21456 17484 21508 17536
rect 22836 17527 22888 17536
rect 22836 17493 22845 17527
rect 22845 17493 22879 17527
rect 22879 17493 22888 17527
rect 22836 17484 22888 17493
rect 23020 17552 23072 17604
rect 23572 17527 23624 17536
rect 23572 17493 23581 17527
rect 23581 17493 23615 17527
rect 23615 17493 23624 17527
rect 23572 17484 23624 17493
rect 26516 17620 26568 17672
rect 24308 17552 24360 17604
rect 26148 17484 26200 17536
rect 28356 17484 28408 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 2228 17280 2280 17332
rect 2688 17280 2740 17332
rect 3240 17212 3292 17264
rect 2044 17144 2096 17196
rect 2136 17144 2188 17196
rect 2320 17144 2372 17196
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 5816 17280 5868 17332
rect 6000 17280 6052 17332
rect 6552 17280 6604 17332
rect 7380 17280 7432 17332
rect 9220 17280 9272 17332
rect 9772 17280 9824 17332
rect 10324 17280 10376 17332
rect 12072 17280 12124 17332
rect 7564 17212 7616 17264
rect 2504 17144 2556 17153
rect 1952 17076 2004 17128
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4712 17144 4764 17196
rect 4804 17144 4856 17196
rect 1584 16940 1636 16992
rect 4436 17076 4488 17128
rect 5080 17144 5132 17196
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6460 17144 6512 17196
rect 7288 17144 7340 17196
rect 10968 17212 11020 17264
rect 11152 17212 11204 17264
rect 12532 17280 12584 17332
rect 13728 17280 13780 17332
rect 16304 17280 16356 17332
rect 16488 17280 16540 17332
rect 13176 17212 13228 17264
rect 13360 17212 13412 17264
rect 13544 17212 13596 17264
rect 13820 17212 13872 17264
rect 13912 17212 13964 17264
rect 17316 17212 17368 17264
rect 8116 17144 8168 17196
rect 8392 17144 8444 17196
rect 8944 17144 8996 17196
rect 9128 17144 9180 17196
rect 9772 17144 9824 17196
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 5080 17008 5132 17060
rect 5172 17051 5224 17060
rect 5172 17017 5181 17051
rect 5181 17017 5215 17051
rect 5215 17017 5224 17051
rect 5172 17008 5224 17017
rect 3332 16940 3384 16992
rect 5816 16940 5868 16992
rect 6736 16940 6788 16992
rect 10048 17076 10100 17128
rect 7196 17008 7248 17060
rect 7656 17008 7708 17060
rect 9680 17008 9732 17060
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 11428 17144 11480 17196
rect 12256 17076 12308 17128
rect 12992 17076 13044 17128
rect 13268 17076 13320 17128
rect 10784 17008 10836 17060
rect 8300 16940 8352 16992
rect 10140 16940 10192 16992
rect 12072 16940 12124 16992
rect 13820 17008 13872 17060
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 17040 17144 17092 17196
rect 18236 17212 18288 17264
rect 20444 17323 20496 17332
rect 20444 17289 20453 17323
rect 20453 17289 20487 17323
rect 20487 17289 20496 17323
rect 20444 17280 20496 17289
rect 22284 17280 22336 17332
rect 22376 17212 22428 17264
rect 18696 17187 18748 17196
rect 18696 17153 18703 17187
rect 18703 17153 18748 17187
rect 14648 17076 14700 17128
rect 16672 17076 16724 17128
rect 17592 17076 17644 17128
rect 15476 17008 15528 17060
rect 18696 17144 18748 17153
rect 12900 16940 12952 16992
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 14372 16940 14424 16992
rect 14740 16940 14792 16992
rect 16764 16940 16816 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18788 17008 18840 17060
rect 18972 17187 19024 17196
rect 18972 17153 18986 17187
rect 18986 17153 19020 17187
rect 19020 17153 19024 17187
rect 18972 17144 19024 17153
rect 19984 17187 20036 17196
rect 19984 17153 19991 17187
rect 19991 17153 20036 17187
rect 19984 17144 20036 17153
rect 20720 17144 20772 17196
rect 21180 17144 21232 17196
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 20536 17076 20588 17128
rect 21916 17076 21968 17128
rect 26148 17280 26200 17332
rect 22560 17212 22612 17264
rect 23112 17144 23164 17196
rect 25044 17144 25096 17196
rect 26240 17144 26292 17196
rect 22836 17076 22888 17128
rect 22376 17051 22428 17060
rect 22376 17017 22385 17051
rect 22385 17017 22419 17051
rect 22419 17017 22428 17051
rect 22376 17008 22428 17017
rect 22468 17051 22520 17060
rect 22468 17017 22477 17051
rect 22477 17017 22511 17051
rect 22511 17017 22520 17051
rect 22468 17008 22520 17017
rect 21088 16940 21140 16992
rect 24584 17051 24636 17060
rect 24584 17017 24593 17051
rect 24593 17017 24627 17051
rect 24627 17017 24636 17051
rect 24584 17008 24636 17017
rect 27620 17076 27672 17128
rect 27804 17008 27856 17060
rect 26792 16940 26844 16992
rect 27068 16940 27120 16992
rect 27528 16940 27580 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 5356 16736 5408 16788
rect 5540 16736 5592 16788
rect 7012 16736 7064 16788
rect 7196 16736 7248 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 10324 16736 10376 16788
rect 12716 16736 12768 16788
rect 14004 16736 14056 16788
rect 14188 16736 14240 16788
rect 15476 16736 15528 16788
rect 15936 16736 15988 16788
rect 16948 16736 17000 16788
rect 17776 16736 17828 16788
rect 18788 16736 18840 16788
rect 1952 16668 2004 16720
rect 2780 16668 2832 16720
rect 5264 16668 5316 16720
rect 8300 16668 8352 16720
rect 1584 16532 1636 16584
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 3148 16532 3200 16584
rect 3792 16532 3844 16584
rect 6552 16600 6604 16652
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 6644 16600 6696 16609
rect 6736 16600 6788 16652
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 6368 16532 6420 16584
rect 7656 16532 7708 16584
rect 7932 16532 7984 16584
rect 8852 16600 8904 16652
rect 11980 16668 12032 16720
rect 12164 16668 12216 16720
rect 12992 16668 13044 16720
rect 15384 16668 15436 16720
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 10692 16600 10744 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 2504 16464 2556 16516
rect 2596 16464 2648 16516
rect 4160 16464 4212 16516
rect 4252 16439 4304 16448
rect 4252 16405 4261 16439
rect 4261 16405 4295 16439
rect 4295 16405 4304 16439
rect 4252 16396 4304 16405
rect 4712 16507 4764 16516
rect 4712 16473 4721 16507
rect 4721 16473 4755 16507
rect 4755 16473 4764 16507
rect 4712 16464 4764 16473
rect 5172 16396 5224 16448
rect 5724 16396 5776 16448
rect 6460 16396 6512 16448
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7564 16507 7616 16516
rect 7564 16473 7573 16507
rect 7573 16473 7607 16507
rect 7607 16473 7616 16507
rect 7564 16464 7616 16473
rect 7748 16507 7800 16516
rect 7748 16473 7757 16507
rect 7757 16473 7791 16507
rect 7791 16473 7800 16507
rect 7748 16464 7800 16473
rect 9956 16464 10008 16516
rect 10232 16464 10284 16516
rect 12348 16532 12400 16584
rect 12440 16532 12492 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 13084 16532 13136 16584
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 16672 16532 16724 16584
rect 16948 16600 17000 16652
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17592 16600 17644 16652
rect 17776 16600 17828 16652
rect 18052 16600 18104 16652
rect 18972 16668 19024 16720
rect 20720 16668 20772 16720
rect 22284 16711 22336 16720
rect 22284 16677 22293 16711
rect 22293 16677 22327 16711
rect 22327 16677 22336 16711
rect 25688 16736 25740 16788
rect 22284 16668 22336 16677
rect 18696 16532 18748 16584
rect 11060 16464 11112 16516
rect 11428 16507 11480 16516
rect 11428 16473 11437 16507
rect 11437 16473 11471 16507
rect 11471 16473 11480 16507
rect 11428 16464 11480 16473
rect 11520 16507 11572 16516
rect 11520 16473 11529 16507
rect 11529 16473 11563 16507
rect 11563 16473 11572 16507
rect 11520 16464 11572 16473
rect 12164 16464 12216 16516
rect 9404 16396 9456 16448
rect 10048 16396 10100 16448
rect 10692 16396 10744 16448
rect 13360 16507 13412 16516
rect 13360 16473 13369 16507
rect 13369 16473 13403 16507
rect 13403 16473 13412 16507
rect 13360 16464 13412 16473
rect 12992 16396 13044 16448
rect 17868 16464 17920 16516
rect 19248 16600 19300 16652
rect 19892 16600 19944 16652
rect 21180 16600 21232 16652
rect 23848 16668 23900 16720
rect 24584 16600 24636 16652
rect 20904 16532 20956 16584
rect 23388 16532 23440 16584
rect 26792 16736 26844 16788
rect 21180 16507 21232 16516
rect 21180 16473 21189 16507
rect 21189 16473 21223 16507
rect 21223 16473 21232 16507
rect 21180 16464 21232 16473
rect 13544 16439 13596 16448
rect 13544 16405 13569 16439
rect 13569 16405 13596 16439
rect 13544 16396 13596 16405
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 13820 16396 13872 16448
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 16672 16396 16724 16405
rect 16948 16396 17000 16448
rect 20352 16396 20404 16448
rect 20444 16396 20496 16448
rect 20996 16396 21048 16448
rect 21640 16464 21692 16516
rect 21916 16507 21968 16516
rect 21916 16473 21925 16507
rect 21925 16473 21959 16507
rect 21959 16473 21968 16507
rect 21916 16464 21968 16473
rect 22008 16464 22060 16516
rect 23296 16464 23348 16516
rect 24860 16464 24912 16516
rect 26056 16464 26108 16516
rect 23480 16396 23532 16448
rect 24032 16396 24084 16448
rect 24124 16396 24176 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 3792 16192 3844 16244
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 7012 16192 7064 16244
rect 8852 16235 8904 16244
rect 8852 16201 8861 16235
rect 8861 16201 8895 16235
rect 8895 16201 8904 16235
rect 8852 16192 8904 16201
rect 10232 16192 10284 16244
rect 10416 16235 10468 16244
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 10876 16192 10928 16244
rect 11060 16192 11112 16244
rect 11980 16192 12032 16244
rect 12716 16192 12768 16244
rect 14648 16192 14700 16244
rect 14924 16192 14976 16244
rect 5356 16124 5408 16176
rect 1768 16056 1820 16108
rect 2504 16056 2556 16108
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 4068 16056 4120 16108
rect 4712 16056 4764 16108
rect 5264 16056 5316 16108
rect 6276 16124 6328 16176
rect 6460 16124 6512 16176
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 8392 16124 8444 16176
rect 6000 16056 6052 16065
rect 2136 15988 2188 16040
rect 6000 15920 6052 15972
rect 3056 15852 3108 15904
rect 5540 15852 5592 15904
rect 5632 15852 5684 15904
rect 7104 16056 7156 16108
rect 7288 16056 7340 16108
rect 7564 16031 7616 16040
rect 7564 15997 7573 16031
rect 7573 15997 7607 16031
rect 7607 15997 7616 16031
rect 7564 15988 7616 15997
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 13268 16124 13320 16176
rect 9128 16056 9180 16108
rect 10508 16056 10560 16108
rect 10876 16056 10928 16108
rect 11244 16056 11296 16108
rect 12532 16056 12584 16108
rect 10048 15988 10100 16040
rect 10692 15988 10744 16040
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 12808 15988 12860 16040
rect 13176 16056 13228 16108
rect 14464 16124 14516 16176
rect 15200 16056 15252 16108
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 19064 16192 19116 16244
rect 19340 16235 19392 16244
rect 19340 16201 19349 16235
rect 19349 16201 19383 16235
rect 19383 16201 19392 16235
rect 19340 16192 19392 16201
rect 22284 16192 22336 16244
rect 26240 16192 26292 16244
rect 22376 16124 22428 16176
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 17500 16056 17552 16108
rect 17868 16056 17920 16108
rect 18604 16056 18656 16108
rect 19432 16056 19484 16108
rect 17684 15988 17736 16040
rect 20444 16056 20496 16108
rect 20720 16056 20772 16108
rect 8208 15920 8260 15972
rect 8944 15920 8996 15972
rect 12624 15920 12676 15972
rect 13268 15920 13320 15972
rect 17224 15920 17276 15972
rect 20628 15988 20680 16040
rect 22652 16056 22704 16108
rect 23296 16167 23348 16176
rect 23296 16133 23305 16167
rect 23305 16133 23339 16167
rect 23339 16133 23348 16167
rect 23296 16124 23348 16133
rect 27436 16192 27488 16244
rect 25596 16056 25648 16108
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 28172 16099 28224 16108
rect 28172 16065 28181 16099
rect 28181 16065 28215 16099
rect 28215 16065 28224 16099
rect 28172 16056 28224 16065
rect 22560 15988 22612 16040
rect 24032 15988 24084 16040
rect 19432 15920 19484 15972
rect 20352 15920 20404 15972
rect 23572 15920 23624 15972
rect 23664 15963 23716 15972
rect 23664 15929 23673 15963
rect 23673 15929 23707 15963
rect 23707 15929 23716 15963
rect 23664 15920 23716 15929
rect 24124 15920 24176 15972
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 8300 15852 8352 15904
rect 9496 15852 9548 15904
rect 10324 15852 10376 15904
rect 12072 15852 12124 15904
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 13544 15852 13596 15904
rect 14648 15852 14700 15904
rect 17684 15895 17736 15904
rect 17684 15861 17693 15895
rect 17693 15861 17727 15895
rect 17727 15861 17736 15895
rect 17684 15852 17736 15861
rect 17776 15852 17828 15904
rect 20444 15852 20496 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 21824 15852 21876 15904
rect 23296 15852 23348 15904
rect 27712 15852 27764 15904
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1216 15648 1268 15700
rect 2136 15648 2188 15700
rect 2228 15648 2280 15700
rect 4068 15648 4120 15700
rect 6092 15648 6144 15700
rect 8484 15648 8536 15700
rect 14924 15648 14976 15700
rect 16028 15648 16080 15700
rect 3240 15580 3292 15632
rect 4804 15580 4856 15632
rect 7380 15580 7432 15632
rect 8300 15580 8352 15632
rect 14464 15580 14516 15632
rect 16488 15580 16540 15632
rect 17500 15648 17552 15700
rect 17868 15648 17920 15700
rect 20352 15648 20404 15700
rect 2780 15512 2832 15564
rect 3516 15512 3568 15564
rect 5724 15512 5776 15564
rect 480 15444 532 15496
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 4436 15487 4488 15496
rect 4436 15453 4445 15487
rect 4445 15453 4479 15487
rect 4479 15453 4488 15487
rect 4436 15444 4488 15453
rect 4988 15487 5040 15496
rect 4988 15453 5003 15487
rect 5003 15453 5037 15487
rect 5037 15453 5040 15487
rect 4988 15444 5040 15453
rect 5264 15444 5316 15496
rect 5540 15444 5592 15496
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 10416 15512 10468 15564
rect 10968 15512 11020 15564
rect 6000 15444 6052 15496
rect 2780 15376 2832 15428
rect 3240 15376 3292 15428
rect 4804 15376 4856 15428
rect 8300 15444 8352 15496
rect 8576 15444 8628 15496
rect 9680 15444 9732 15496
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 14188 15512 14240 15564
rect 14372 15512 14424 15564
rect 13084 15444 13136 15496
rect 13360 15444 13412 15496
rect 3056 15308 3108 15360
rect 3884 15308 3936 15360
rect 3976 15351 4028 15360
rect 3976 15317 3985 15351
rect 3985 15317 4019 15351
rect 4019 15317 4028 15351
rect 3976 15308 4028 15317
rect 5816 15308 5868 15360
rect 6460 15308 6512 15360
rect 9588 15376 9640 15428
rect 8208 15308 8260 15360
rect 8944 15308 8996 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 12808 15376 12860 15428
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 16304 15512 16356 15564
rect 16764 15512 16816 15564
rect 17684 15580 17736 15632
rect 20168 15580 20220 15632
rect 17224 15512 17276 15564
rect 18420 15512 18472 15564
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 12716 15308 12768 15360
rect 15292 15308 15344 15360
rect 18328 15376 18380 15428
rect 18420 15419 18472 15428
rect 18420 15385 18429 15419
rect 18429 15385 18463 15419
rect 18463 15385 18472 15419
rect 18420 15376 18472 15385
rect 18972 15444 19024 15496
rect 18696 15376 18748 15428
rect 18788 15376 18840 15428
rect 20076 15512 20128 15564
rect 21180 15648 21232 15700
rect 21364 15648 21416 15700
rect 21824 15623 21876 15632
rect 21824 15589 21833 15623
rect 21833 15589 21867 15623
rect 21867 15589 21876 15623
rect 21824 15580 21876 15589
rect 24952 15648 25004 15700
rect 25596 15648 25648 15700
rect 22744 15512 22796 15564
rect 25964 15623 26016 15632
rect 25964 15589 25973 15623
rect 25973 15589 26007 15623
rect 26007 15589 26016 15623
rect 25964 15580 26016 15589
rect 20168 15444 20220 15496
rect 15568 15308 15620 15360
rect 16856 15308 16908 15360
rect 17316 15308 17368 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 21548 15444 21600 15496
rect 21640 15444 21692 15496
rect 21088 15376 21140 15428
rect 24032 15444 24084 15496
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 25780 15444 25832 15496
rect 26424 15444 26476 15496
rect 27068 15487 27120 15496
rect 27068 15453 27102 15487
rect 27102 15453 27120 15487
rect 27068 15444 27120 15453
rect 21180 15308 21232 15360
rect 21548 15308 21600 15360
rect 23204 15376 23256 15428
rect 28080 15376 28132 15428
rect 23480 15308 23532 15360
rect 27528 15308 27580 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 1860 15104 1912 15156
rect 3516 15104 3568 15156
rect 5632 15104 5684 15156
rect 1676 15036 1728 15088
rect 6736 15104 6788 15156
rect 7196 15104 7248 15156
rect 7564 15147 7616 15156
rect 7564 15113 7573 15147
rect 7573 15113 7607 15147
rect 7607 15113 7616 15147
rect 7564 15104 7616 15113
rect 8208 15147 8260 15156
rect 8208 15113 8217 15147
rect 8217 15113 8251 15147
rect 8251 15113 8260 15147
rect 8208 15104 8260 15113
rect 8852 15104 8904 15156
rect 9036 15104 9088 15156
rect 12440 15104 12492 15156
rect 12992 15104 13044 15156
rect 13084 15104 13136 15156
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 4344 14968 4396 15020
rect 3332 14900 3384 14952
rect 3792 14900 3844 14952
rect 4436 14900 4488 14952
rect 5724 14900 5776 14952
rect 2688 14832 2740 14884
rect 5356 14832 5408 14884
rect 10784 15036 10836 15088
rect 6736 14968 6788 15020
rect 8300 15011 8352 15020
rect 8300 14977 8309 15011
rect 8309 14977 8343 15011
rect 8343 14977 8352 15011
rect 8300 14968 8352 14977
rect 8392 14968 8444 15020
rect 9772 14968 9824 15020
rect 10232 14968 10284 15020
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 12256 15036 12308 15088
rect 12624 14968 12676 15020
rect 13820 15036 13872 15088
rect 13360 14968 13412 15020
rect 13544 14968 13596 15020
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 14740 15104 14792 15156
rect 15016 15104 15068 15156
rect 16028 15147 16080 15156
rect 16028 15113 16037 15147
rect 16037 15113 16071 15147
rect 16071 15113 16080 15147
rect 16028 15104 16080 15113
rect 17868 15104 17920 15156
rect 20720 15104 20772 15156
rect 16856 15036 16908 15088
rect 17040 15036 17092 15088
rect 14740 14968 14792 15020
rect 8576 14900 8628 14952
rect 15752 14968 15804 15020
rect 16580 14968 16632 15020
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 18052 14968 18104 15020
rect 19800 15036 19852 15088
rect 19892 15036 19944 15088
rect 24860 15104 24912 15156
rect 28172 15104 28224 15156
rect 21640 15036 21692 15088
rect 25872 15036 25924 15088
rect 27804 15036 27856 15088
rect 18328 14968 18380 15020
rect 20536 14968 20588 15020
rect 2596 14764 2648 14816
rect 4252 14764 4304 14816
rect 9220 14832 9272 14884
rect 9680 14832 9732 14884
rect 11704 14832 11756 14884
rect 5724 14764 5776 14816
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 8852 14764 8904 14816
rect 10600 14764 10652 14816
rect 11796 14764 11848 14816
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 14556 14832 14608 14884
rect 15108 14832 15160 14884
rect 17040 14900 17092 14952
rect 18144 14900 18196 14952
rect 16120 14832 16172 14884
rect 12256 14764 12308 14816
rect 14280 14764 14332 14816
rect 15292 14764 15344 14816
rect 15936 14764 15988 14816
rect 19984 14900 20036 14952
rect 20352 14832 20404 14884
rect 21548 14968 21600 15020
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 22468 15011 22520 15020
rect 22468 14977 22503 15011
rect 22503 14977 22520 15011
rect 22468 14968 22520 14977
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 23480 14968 23532 15020
rect 20996 14900 21048 14952
rect 19800 14764 19852 14816
rect 20076 14807 20128 14816
rect 20076 14773 20085 14807
rect 20085 14773 20119 14807
rect 20119 14773 20128 14807
rect 20076 14764 20128 14773
rect 20260 14764 20312 14816
rect 20628 14764 20680 14816
rect 21272 14764 21324 14816
rect 23664 14832 23716 14884
rect 23756 14764 23808 14816
rect 23940 14943 23992 14952
rect 23940 14909 23949 14943
rect 23949 14909 23983 14943
rect 23983 14909 23992 14943
rect 23940 14900 23992 14909
rect 27528 14900 27580 14952
rect 25964 14832 26016 14884
rect 27436 14764 27488 14816
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1952 14560 2004 14612
rect 4160 14560 4212 14612
rect 5264 14560 5316 14612
rect 6368 14560 6420 14612
rect 8024 14560 8076 14612
rect 8668 14560 8720 14612
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 12716 14560 12768 14612
rect 13728 14560 13780 14612
rect 13820 14560 13872 14612
rect 15752 14560 15804 14612
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 16212 14560 16264 14612
rect 17960 14560 18012 14612
rect 20352 14560 20404 14612
rect 4068 14492 4120 14544
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 3976 14424 4028 14476
rect 2688 14288 2740 14340
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 7748 14492 7800 14544
rect 7840 14492 7892 14544
rect 5080 14424 5132 14476
rect 6920 14424 6972 14476
rect 4804 14356 4856 14408
rect 4896 14288 4948 14340
rect 5724 14356 5776 14408
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 7104 14356 7156 14408
rect 7196 14356 7248 14408
rect 9036 14424 9088 14476
rect 10232 14356 10284 14408
rect 11796 14492 11848 14544
rect 11980 14492 12032 14544
rect 12256 14492 12308 14544
rect 10876 14424 10928 14476
rect 11244 14424 11296 14476
rect 11520 14424 11572 14476
rect 12900 14424 12952 14476
rect 6460 14288 6512 14340
rect 10876 14288 10928 14340
rect 11152 14331 11204 14340
rect 11152 14297 11161 14331
rect 11161 14297 11195 14331
rect 11195 14297 11204 14331
rect 11152 14288 11204 14297
rect 11336 14331 11388 14340
rect 11336 14297 11361 14331
rect 11361 14297 11388 14331
rect 12256 14356 12308 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 11336 14288 11388 14297
rect 13268 14356 13320 14408
rect 13912 14492 13964 14544
rect 16028 14492 16080 14544
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14648 14424 14700 14476
rect 14556 14356 14608 14408
rect 15108 14356 15160 14408
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 2964 14220 3016 14272
rect 5172 14220 5224 14272
rect 7012 14220 7064 14272
rect 8760 14220 8812 14272
rect 9128 14220 9180 14272
rect 9220 14220 9272 14272
rect 9496 14220 9548 14272
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 10784 14220 10836 14272
rect 15384 14288 15436 14340
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 17040 14424 17092 14476
rect 18052 14492 18104 14544
rect 20628 14603 20680 14612
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 25964 14560 26016 14612
rect 20076 14424 20128 14476
rect 17132 14356 17184 14408
rect 11980 14220 12032 14272
rect 14188 14220 14240 14272
rect 14464 14220 14516 14272
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 18972 14356 19024 14408
rect 19616 14356 19668 14408
rect 17960 14288 18012 14340
rect 19064 14288 19116 14340
rect 19156 14220 19208 14272
rect 20168 14220 20220 14272
rect 20720 14288 20772 14340
rect 21548 14356 21600 14408
rect 22836 14492 22888 14544
rect 23388 14535 23440 14544
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 23572 14492 23624 14544
rect 22928 14356 22980 14408
rect 24952 14356 25004 14408
rect 26332 14356 26384 14408
rect 20812 14220 20864 14272
rect 22560 14288 22612 14340
rect 23112 14331 23164 14340
rect 23112 14297 23121 14331
rect 23121 14297 23155 14331
rect 23155 14297 23164 14331
rect 23112 14288 23164 14297
rect 22284 14220 22336 14272
rect 23572 14263 23624 14272
rect 23572 14229 23581 14263
rect 23581 14229 23615 14263
rect 23615 14229 23624 14263
rect 23572 14220 23624 14229
rect 23756 14220 23808 14272
rect 24492 14220 24544 14272
rect 26700 14220 26752 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2320 14016 2372 14068
rect 6460 14016 6512 14068
rect 2504 13880 2556 13932
rect 2780 13812 2832 13864
rect 4068 13948 4120 14000
rect 3884 13880 3936 13932
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 3976 13812 4028 13864
rect 4252 13812 4304 13864
rect 4896 13880 4948 13932
rect 5080 13880 5132 13932
rect 7840 14016 7892 14068
rect 8208 14016 8260 14068
rect 9220 14016 9272 14068
rect 7564 13948 7616 14000
rect 3056 13744 3108 13796
rect 3332 13787 3384 13796
rect 3332 13753 3341 13787
rect 3341 13753 3375 13787
rect 3375 13753 3384 13787
rect 3332 13744 3384 13753
rect 4896 13744 4948 13796
rect 5724 13812 5776 13864
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 9496 13948 9548 14000
rect 10140 14016 10192 14068
rect 10232 14016 10284 14068
rect 11796 14016 11848 14068
rect 11888 14016 11940 14068
rect 12716 13948 12768 14000
rect 13544 14059 13596 14068
rect 13544 14025 13553 14059
rect 13553 14025 13587 14059
rect 13587 14025 13596 14059
rect 13544 14016 13596 14025
rect 13820 14016 13872 14068
rect 8760 13880 8812 13932
rect 8024 13812 8076 13864
rect 9588 13880 9640 13932
rect 10692 13880 10744 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11152 13880 11204 13932
rect 12348 13880 12400 13932
rect 12900 13880 12952 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 15660 13991 15712 14000
rect 15660 13957 15685 13991
rect 15685 13957 15712 13991
rect 15844 14059 15896 14068
rect 15844 14025 15853 14059
rect 15853 14025 15887 14059
rect 15887 14025 15896 14059
rect 15844 14016 15896 14025
rect 16580 14016 16632 14068
rect 19064 14016 19116 14068
rect 22192 14016 22244 14068
rect 15660 13948 15712 13957
rect 17316 13948 17368 14000
rect 9772 13812 9824 13864
rect 10876 13812 10928 13864
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 6644 13744 6696 13796
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 7012 13744 7064 13753
rect 10416 13744 10468 13796
rect 11520 13744 11572 13796
rect 14188 13744 14240 13796
rect 15568 13880 15620 13932
rect 16028 13880 16080 13932
rect 16856 13880 16908 13932
rect 17960 13948 18012 14000
rect 18328 13880 18380 13932
rect 18696 13948 18748 14000
rect 20168 13991 20220 14000
rect 20168 13957 20177 13991
rect 20177 13957 20211 13991
rect 20211 13957 20220 13991
rect 20168 13948 20220 13957
rect 23572 14016 23624 14068
rect 24216 14016 24268 14068
rect 24492 14016 24544 14068
rect 28080 14059 28132 14068
rect 28080 14025 28089 14059
rect 28089 14025 28123 14059
rect 28123 14025 28132 14059
rect 28080 14016 28132 14025
rect 19156 13880 19208 13932
rect 19892 13923 19944 13932
rect 19892 13889 19901 13923
rect 19901 13889 19935 13923
rect 19935 13889 19944 13923
rect 19892 13880 19944 13889
rect 19984 13923 20036 13932
rect 19984 13889 19994 13923
rect 19994 13889 20028 13923
rect 20028 13889 20036 13923
rect 19984 13880 20036 13889
rect 15476 13812 15528 13864
rect 15752 13812 15804 13864
rect 19616 13812 19668 13864
rect 20536 13880 20588 13932
rect 21272 13880 21324 13932
rect 22468 13991 22520 14000
rect 22468 13957 22503 13991
rect 22503 13957 22520 13991
rect 25504 13991 25556 14000
rect 22468 13948 22520 13957
rect 25504 13957 25538 13991
rect 25538 13957 25556 13991
rect 25504 13948 25556 13957
rect 21548 13880 21600 13932
rect 20628 13812 20680 13864
rect 22100 13812 22152 13864
rect 16948 13744 17000 13796
rect 17500 13744 17552 13796
rect 4988 13676 5040 13728
rect 5264 13676 5316 13728
rect 5448 13676 5500 13728
rect 6460 13676 6512 13728
rect 9312 13676 9364 13728
rect 10968 13676 11020 13728
rect 12072 13676 12124 13728
rect 12624 13676 12676 13728
rect 13268 13676 13320 13728
rect 13728 13676 13780 13728
rect 15292 13676 15344 13728
rect 15660 13719 15712 13728
rect 15660 13685 15669 13719
rect 15669 13685 15703 13719
rect 15703 13685 15712 13719
rect 15660 13676 15712 13685
rect 17132 13676 17184 13728
rect 17776 13719 17828 13728
rect 17776 13685 17785 13719
rect 17785 13685 17819 13719
rect 17819 13685 17828 13719
rect 17776 13676 17828 13685
rect 18512 13676 18564 13728
rect 19616 13676 19668 13728
rect 21640 13744 21692 13796
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23112 13812 23164 13821
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 28264 13923 28316 13932
rect 28264 13889 28273 13923
rect 28273 13889 28307 13923
rect 28307 13889 28316 13923
rect 28264 13880 28316 13889
rect 24952 13812 25004 13864
rect 25136 13812 25188 13864
rect 27160 13855 27212 13864
rect 27160 13821 27169 13855
rect 27169 13821 27203 13855
rect 27203 13821 27212 13855
rect 27160 13812 27212 13821
rect 22836 13744 22888 13796
rect 22560 13676 22612 13728
rect 22744 13676 22796 13728
rect 23572 13719 23624 13728
rect 23572 13685 23581 13719
rect 23581 13685 23615 13719
rect 23615 13685 23624 13719
rect 23572 13676 23624 13685
rect 27436 13787 27488 13796
rect 27436 13753 27445 13787
rect 27445 13753 27479 13787
rect 27479 13753 27488 13787
rect 27436 13744 27488 13753
rect 25044 13676 25096 13728
rect 27620 13719 27672 13728
rect 27620 13685 27629 13719
rect 27629 13685 27663 13719
rect 27663 13685 27672 13719
rect 27620 13676 27672 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 2044 13472 2096 13524
rect 3148 13472 3200 13524
rect 5264 13472 5316 13524
rect 5816 13472 5868 13524
rect 4712 13404 4764 13456
rect 4896 13404 4948 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 5172 13336 5224 13388
rect 5448 13336 5500 13388
rect 6552 13404 6604 13456
rect 9864 13472 9916 13524
rect 11152 13472 11204 13524
rect 11336 13472 11388 13524
rect 9496 13404 9548 13456
rect 9588 13447 9640 13456
rect 9588 13413 9597 13447
rect 9597 13413 9631 13447
rect 9631 13413 9640 13447
rect 9588 13404 9640 13413
rect 12164 13404 12216 13456
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 17408 13472 17460 13524
rect 13820 13404 13872 13456
rect 16672 13404 16724 13456
rect 17776 13447 17828 13456
rect 17776 13413 17785 13447
rect 17785 13413 17819 13447
rect 17819 13413 17828 13447
rect 17776 13404 17828 13413
rect 6920 13336 6972 13388
rect 4068 13268 4120 13320
rect 3608 13200 3660 13252
rect 4620 13268 4672 13320
rect 4896 13268 4948 13320
rect 5632 13268 5684 13320
rect 4160 13132 4212 13184
rect 4620 13132 4672 13184
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 6276 13243 6328 13252
rect 6276 13209 6285 13243
rect 6285 13209 6319 13243
rect 6319 13209 6328 13243
rect 6276 13200 6328 13209
rect 6460 13243 6512 13252
rect 6460 13209 6469 13243
rect 6469 13209 6503 13243
rect 6503 13209 6512 13243
rect 6460 13200 6512 13209
rect 6368 13132 6420 13184
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 7840 13336 7892 13388
rect 10140 13336 10192 13388
rect 10968 13336 11020 13388
rect 11152 13336 11204 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 7656 13268 7708 13320
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 8484 13268 8536 13320
rect 8668 13268 8720 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 9496 13268 9548 13320
rect 10508 13268 10560 13320
rect 12348 13268 12400 13320
rect 12440 13268 12492 13320
rect 13452 13268 13504 13320
rect 8760 13132 8812 13184
rect 11336 13200 11388 13252
rect 11796 13200 11848 13252
rect 14004 13200 14056 13252
rect 15476 13200 15528 13252
rect 11152 13132 11204 13184
rect 11428 13132 11480 13184
rect 12348 13132 12400 13184
rect 13360 13132 13412 13184
rect 13452 13132 13504 13184
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 19340 13336 19392 13388
rect 17597 13311 17649 13320
rect 17597 13277 17606 13311
rect 17606 13277 17640 13311
rect 17640 13277 17649 13311
rect 17597 13268 17649 13277
rect 17960 13268 18012 13320
rect 18788 13268 18840 13320
rect 20628 13336 20680 13388
rect 21548 13472 21600 13524
rect 23112 13472 23164 13524
rect 23940 13472 23992 13524
rect 24216 13472 24268 13524
rect 20996 13404 21048 13456
rect 22744 13447 22796 13456
rect 22744 13413 22753 13447
rect 22753 13413 22787 13447
rect 22787 13413 22796 13447
rect 22744 13404 22796 13413
rect 24860 13472 24912 13524
rect 24952 13472 25004 13524
rect 26148 13472 26200 13524
rect 23940 13336 23992 13388
rect 16948 13200 17000 13252
rect 19248 13200 19300 13252
rect 19892 13200 19944 13252
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 20536 13268 20588 13320
rect 22744 13268 22796 13320
rect 20996 13200 21048 13252
rect 21088 13243 21140 13252
rect 21088 13209 21097 13243
rect 21097 13209 21131 13243
rect 21131 13209 21140 13243
rect 21088 13200 21140 13209
rect 23112 13200 23164 13252
rect 23848 13200 23900 13252
rect 24032 13268 24084 13320
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 27160 13472 27212 13524
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26700 13311 26752 13320
rect 26700 13277 26734 13311
rect 26734 13277 26752 13311
rect 26700 13268 26752 13277
rect 16028 13132 16080 13184
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 16764 13132 16816 13184
rect 18236 13132 18288 13184
rect 19524 13132 19576 13184
rect 20720 13132 20772 13184
rect 24676 13132 24728 13184
rect 28080 13200 28132 13252
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 1860 12928 1912 12980
rect 3424 12971 3476 12980
rect 3424 12937 3449 12971
rect 3449 12937 3476 12971
rect 3424 12928 3476 12937
rect 4344 12928 4396 12980
rect 5356 12928 5408 12980
rect 5724 12928 5776 12980
rect 7472 12971 7524 12980
rect 7472 12937 7481 12971
rect 7481 12937 7515 12971
rect 7515 12937 7524 12971
rect 7472 12928 7524 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 8944 12928 8996 12980
rect 10324 12928 10376 12980
rect 2320 12792 2372 12844
rect 2688 12860 2740 12912
rect 3056 12792 3108 12844
rect 4896 12860 4948 12912
rect 6276 12860 6328 12912
rect 8392 12860 8444 12912
rect 10784 12928 10836 12980
rect 10968 12928 11020 12980
rect 11152 12928 11204 12980
rect 11612 12928 11664 12980
rect 3608 12792 3660 12844
rect 4804 12792 4856 12844
rect 2964 12724 3016 12776
rect 3240 12724 3292 12776
rect 3148 12656 3200 12708
rect 4252 12724 4304 12776
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 4712 12724 4764 12733
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 6552 12792 6604 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 5356 12724 5408 12776
rect 7564 12724 7616 12776
rect 8760 12792 8812 12844
rect 13820 12928 13872 12980
rect 14004 12928 14056 12980
rect 14740 12928 14792 12980
rect 16488 12928 16540 12980
rect 18880 12971 18932 12980
rect 18880 12937 18889 12971
rect 18889 12937 18923 12971
rect 18923 12937 18932 12971
rect 18880 12928 18932 12937
rect 19156 12928 19208 12980
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 11152 12792 11204 12844
rect 11612 12792 11664 12844
rect 8668 12724 8720 12776
rect 9864 12724 9916 12776
rect 10048 12724 10100 12776
rect 11428 12724 11480 12776
rect 12900 12860 12952 12912
rect 14372 12860 14424 12912
rect 16304 12860 16356 12912
rect 12808 12835 12860 12844
rect 12808 12801 12842 12835
rect 12842 12801 12860 12835
rect 12808 12792 12860 12801
rect 13820 12792 13872 12844
rect 14280 12792 14332 12844
rect 14740 12792 14792 12844
rect 15108 12792 15160 12844
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 16212 12792 16264 12844
rect 17500 12860 17552 12912
rect 17592 12860 17644 12912
rect 17960 12903 18012 12912
rect 17960 12869 17969 12903
rect 17969 12869 18003 12903
rect 18003 12869 18012 12903
rect 17960 12860 18012 12869
rect 18144 12903 18196 12912
rect 18144 12869 18169 12903
rect 18169 12869 18196 12903
rect 19708 12928 19760 12980
rect 20076 12928 20128 12980
rect 20720 12928 20772 12980
rect 24032 12928 24084 12980
rect 18144 12860 18196 12869
rect 20812 12860 20864 12912
rect 5816 12656 5868 12708
rect 5908 12656 5960 12708
rect 6460 12656 6512 12708
rect 8208 12656 8260 12708
rect 13636 12724 13688 12776
rect 17040 12792 17092 12844
rect 17684 12792 17736 12844
rect 17592 12724 17644 12776
rect 4068 12588 4120 12640
rect 6368 12588 6420 12640
rect 6736 12588 6788 12640
rect 7840 12588 7892 12640
rect 8392 12588 8444 12640
rect 8852 12588 8904 12640
rect 9036 12588 9088 12640
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 10232 12588 10284 12640
rect 11060 12588 11112 12640
rect 12164 12588 12216 12640
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 15752 12588 15804 12640
rect 18788 12724 18840 12776
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 19156 12767 19208 12776
rect 19156 12733 19165 12767
rect 19165 12733 19199 12767
rect 19199 12733 19208 12767
rect 19156 12724 19208 12733
rect 19340 12767 19392 12776
rect 19340 12733 19349 12767
rect 19349 12733 19383 12767
rect 19383 12733 19392 12767
rect 19340 12724 19392 12733
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 20628 12792 20680 12844
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 22560 12860 22612 12912
rect 27988 12928 28040 12980
rect 28080 12971 28132 12980
rect 28080 12937 28089 12971
rect 28089 12937 28123 12971
rect 28123 12937 28132 12971
rect 28080 12928 28132 12937
rect 24584 12860 24636 12912
rect 22468 12792 22520 12844
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 23664 12792 23716 12844
rect 26424 12860 26476 12912
rect 27160 12903 27212 12912
rect 27160 12869 27169 12903
rect 27169 12869 27203 12903
rect 27203 12869 27212 12903
rect 27160 12860 27212 12869
rect 25320 12792 25372 12844
rect 27620 12792 27672 12844
rect 19984 12656 20036 12708
rect 20168 12656 20220 12708
rect 18604 12588 18656 12640
rect 19156 12588 19208 12640
rect 20904 12724 20956 12776
rect 23480 12656 23532 12708
rect 26240 12656 26292 12708
rect 20720 12588 20772 12640
rect 22376 12631 22428 12640
rect 22376 12597 22385 12631
rect 22385 12597 22419 12631
rect 22419 12597 22428 12631
rect 22376 12588 22428 12597
rect 22468 12631 22520 12640
rect 22468 12597 22477 12631
rect 22477 12597 22511 12631
rect 22511 12597 22520 12631
rect 22468 12588 22520 12597
rect 23296 12588 23348 12640
rect 26700 12588 26752 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 4252 12384 4304 12436
rect 5080 12384 5132 12436
rect 2412 12248 2464 12300
rect 3148 12248 3200 12300
rect 3884 12248 3936 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4712 12248 4764 12300
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 6092 12384 6144 12436
rect 6552 12384 6604 12436
rect 1952 12155 2004 12164
rect 1952 12121 1961 12155
rect 1961 12121 1995 12155
rect 1995 12121 2004 12155
rect 1952 12112 2004 12121
rect 2228 12112 2280 12164
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 5080 12180 5132 12232
rect 3240 12044 3292 12096
rect 4344 12044 4396 12096
rect 5908 12044 5960 12096
rect 6460 12248 6512 12300
rect 6828 12248 6880 12300
rect 6644 12180 6696 12232
rect 10140 12384 10192 12436
rect 11152 12384 11204 12436
rect 7288 12359 7340 12368
rect 7288 12325 7297 12359
rect 7297 12325 7331 12359
rect 7331 12325 7340 12359
rect 7288 12316 7340 12325
rect 7656 12316 7708 12368
rect 8116 12316 8168 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 8392 12316 8444 12368
rect 10324 12316 10376 12368
rect 11060 12316 11112 12368
rect 12348 12359 12400 12368
rect 12348 12325 12357 12359
rect 12357 12325 12391 12359
rect 12391 12325 12400 12359
rect 12348 12316 12400 12325
rect 12808 12384 12860 12436
rect 14464 12384 14516 12436
rect 14188 12316 14240 12368
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7288 12180 7340 12232
rect 7840 12180 7892 12232
rect 9220 12248 9272 12300
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 10048 12248 10100 12300
rect 10232 12180 10284 12232
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 15108 12359 15160 12368
rect 15108 12325 15117 12359
rect 15117 12325 15151 12359
rect 15151 12325 15160 12359
rect 15108 12316 15160 12325
rect 16396 12316 16448 12368
rect 18144 12384 18196 12436
rect 18328 12384 18380 12436
rect 18512 12384 18564 12436
rect 19432 12384 19484 12436
rect 19708 12384 19760 12436
rect 19892 12384 19944 12436
rect 22100 12384 22152 12436
rect 23480 12384 23532 12436
rect 23848 12384 23900 12436
rect 25044 12384 25096 12436
rect 18236 12316 18288 12368
rect 19984 12316 20036 12368
rect 20904 12316 20956 12368
rect 21548 12316 21600 12368
rect 22928 12316 22980 12368
rect 23388 12316 23440 12368
rect 23756 12316 23808 12368
rect 10692 12180 10744 12232
rect 10876 12180 10928 12232
rect 8300 12112 8352 12164
rect 9588 12112 9640 12164
rect 10416 12112 10468 12164
rect 10784 12112 10836 12164
rect 14280 12180 14332 12232
rect 14372 12180 14424 12232
rect 12072 12112 12124 12164
rect 13452 12112 13504 12164
rect 14832 12112 14884 12164
rect 15108 12180 15160 12232
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 15660 12180 15712 12232
rect 15200 12112 15252 12164
rect 16488 12155 16540 12164
rect 16488 12121 16497 12155
rect 16497 12121 16531 12155
rect 16531 12121 16540 12155
rect 16488 12112 16540 12121
rect 18328 12248 18380 12300
rect 20076 12248 20128 12300
rect 16856 12180 16908 12232
rect 20720 12180 20772 12232
rect 21456 12248 21508 12300
rect 23572 12248 23624 12300
rect 22284 12180 22336 12232
rect 16948 12112 17000 12164
rect 17960 12112 18012 12164
rect 18236 12155 18288 12164
rect 18236 12121 18245 12155
rect 18245 12121 18279 12155
rect 18279 12121 18288 12155
rect 18236 12112 18288 12121
rect 8944 12044 8996 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9864 12044 9916 12096
rect 10876 12044 10928 12096
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11796 12044 11848 12096
rect 13084 12044 13136 12096
rect 15844 12044 15896 12096
rect 16580 12044 16632 12096
rect 18144 12044 18196 12096
rect 19064 12112 19116 12164
rect 18696 12044 18748 12096
rect 19432 12155 19484 12164
rect 19432 12121 19441 12155
rect 19441 12121 19475 12155
rect 19475 12121 19484 12155
rect 19432 12112 19484 12121
rect 19984 12112 20036 12164
rect 20904 12112 20956 12164
rect 21364 12112 21416 12164
rect 23480 12180 23532 12232
rect 22468 12112 22520 12164
rect 23020 12112 23072 12164
rect 19800 12087 19852 12096
rect 19800 12053 19809 12087
rect 19809 12053 19843 12087
rect 19843 12053 19852 12087
rect 19800 12044 19852 12053
rect 20168 12044 20220 12096
rect 20536 12044 20588 12096
rect 23204 12044 23256 12096
rect 26332 12248 26384 12300
rect 26424 12248 26476 12300
rect 24676 12180 24728 12232
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 388 11840 440 11892
rect 940 11840 992 11892
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3056 11840 3108 11892
rect 3516 11840 3568 11892
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 2136 11772 2188 11824
rect 3884 11840 3936 11892
rect 4712 11840 4764 11892
rect 4160 11772 4212 11824
rect 8668 11840 8720 11892
rect 940 11704 992 11756
rect 1124 11704 1176 11756
rect 2412 11704 2464 11756
rect 664 11636 716 11688
rect 1216 11636 1268 11688
rect 2044 11636 2096 11688
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3516 11704 3568 11756
rect 2964 11636 3016 11688
rect 4712 11704 4764 11756
rect 5172 11704 5224 11756
rect 7656 11772 7708 11824
rect 8484 11772 8536 11824
rect 9680 11840 9732 11892
rect 12072 11840 12124 11892
rect 12256 11840 12308 11892
rect 5540 11704 5592 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 6460 11704 6512 11756
rect 6828 11704 6880 11756
rect 7288 11704 7340 11756
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8944 11747 8996 11756
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 11244 11772 11296 11824
rect 15476 11840 15528 11892
rect 16488 11840 16540 11892
rect 4068 11636 4120 11688
rect 1124 11568 1176 11620
rect 6644 11568 6696 11620
rect 7012 11636 7064 11688
rect 10416 11704 10468 11756
rect 1216 11500 1268 11552
rect 2872 11500 2924 11552
rect 3608 11500 3660 11552
rect 3700 11500 3752 11552
rect 6552 11500 6604 11552
rect 7472 11500 7524 11552
rect 7840 11611 7892 11620
rect 7840 11577 7849 11611
rect 7849 11577 7883 11611
rect 7883 11577 7892 11611
rect 7840 11568 7892 11577
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 10232 11636 10284 11688
rect 11612 11704 11664 11756
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 14096 11772 14148 11824
rect 14188 11772 14240 11824
rect 14372 11772 14424 11824
rect 15384 11772 15436 11824
rect 17960 11840 18012 11892
rect 18696 11840 18748 11892
rect 18972 11840 19024 11892
rect 20260 11840 20312 11892
rect 20352 11840 20404 11892
rect 21640 11840 21692 11892
rect 24860 11840 24912 11892
rect 28264 11840 28316 11892
rect 19248 11772 19300 11824
rect 20168 11772 20220 11824
rect 20720 11772 20772 11824
rect 21548 11772 21600 11824
rect 26240 11772 26292 11824
rect 27528 11772 27580 11824
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14832 11704 14884 11756
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15568 11704 15620 11756
rect 8208 11568 8260 11620
rect 8300 11500 8352 11552
rect 8944 11500 8996 11552
rect 13636 11568 13688 11620
rect 10232 11500 10284 11552
rect 13912 11500 13964 11552
rect 15384 11568 15436 11620
rect 16764 11704 16816 11756
rect 17500 11704 17552 11756
rect 19064 11704 19116 11756
rect 19800 11704 19852 11756
rect 18236 11636 18288 11688
rect 18420 11636 18472 11688
rect 18788 11568 18840 11620
rect 19984 11636 20036 11688
rect 16212 11500 16264 11552
rect 19892 11568 19944 11620
rect 21180 11568 21232 11620
rect 21548 11568 21600 11620
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 22008 11636 22060 11688
rect 26700 11704 26752 11756
rect 23664 11679 23716 11688
rect 23664 11645 23673 11679
rect 23673 11645 23707 11679
rect 23707 11645 23716 11679
rect 23664 11636 23716 11645
rect 23112 11568 23164 11620
rect 24676 11568 24728 11620
rect 22468 11500 22520 11552
rect 25136 11500 25188 11552
rect 27712 11611 27764 11620
rect 27712 11577 27721 11611
rect 27721 11577 27755 11611
rect 27755 11577 27764 11611
rect 27712 11568 27764 11577
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 3976 11339 4028 11348
rect 3976 11305 3985 11339
rect 3985 11305 4019 11339
rect 4019 11305 4028 11339
rect 3976 11296 4028 11305
rect 4896 11296 4948 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 7288 11296 7340 11348
rect 3240 11228 3292 11280
rect 3424 11228 3476 11280
rect 1860 11160 1912 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 4252 11160 4304 11212
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2320 11024 2372 11076
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2872 11024 2924 11076
rect 2964 10956 3016 11008
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 5264 11228 5316 11280
rect 5816 11160 5868 11212
rect 6460 11228 6512 11280
rect 7564 11228 7616 11280
rect 6276 11160 6328 11212
rect 6552 11160 6604 11212
rect 4896 11092 4948 11144
rect 5264 11092 5316 11144
rect 5448 11024 5500 11076
rect 5632 11024 5684 11076
rect 6092 11024 6144 11076
rect 6552 11024 6604 11076
rect 4160 10956 4212 11008
rect 4436 10956 4488 11008
rect 5908 10956 5960 11008
rect 6000 10956 6052 11008
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 9956 11296 10008 11348
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 10876 11296 10928 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 12624 11296 12676 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 13360 11296 13412 11348
rect 13912 11296 13964 11348
rect 14924 11296 14976 11348
rect 15476 11296 15528 11348
rect 15936 11296 15988 11348
rect 16672 11296 16724 11348
rect 12532 11228 12584 11280
rect 8668 11160 8720 11212
rect 10232 11092 10284 11144
rect 9404 11067 9456 11076
rect 9404 11033 9413 11067
rect 9413 11033 9447 11067
rect 9447 11033 9456 11067
rect 9404 11024 9456 11033
rect 11980 11160 12032 11212
rect 15660 11228 15712 11280
rect 15844 11228 15896 11280
rect 11796 11092 11848 11144
rect 11888 11092 11940 11144
rect 13544 11160 13596 11212
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 14832 11160 14884 11212
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 18236 11228 18288 11280
rect 20168 11296 20220 11348
rect 19340 11228 19392 11280
rect 24032 11339 24084 11348
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 26240 11339 26292 11348
rect 26240 11305 26249 11339
rect 26249 11305 26283 11339
rect 26283 11305 26292 11339
rect 26240 11296 26292 11305
rect 21640 11228 21692 11280
rect 22008 11271 22060 11280
rect 22008 11237 22017 11271
rect 22017 11237 22051 11271
rect 22051 11237 22060 11271
rect 22008 11228 22060 11237
rect 22560 11228 22612 11280
rect 17500 11160 17552 11212
rect 12992 11092 13044 11144
rect 8576 10956 8628 11008
rect 11060 11024 11112 11076
rect 13636 11092 13688 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 13728 11024 13780 11076
rect 15200 11067 15252 11076
rect 15200 11033 15235 11067
rect 15235 11033 15252 11067
rect 15200 11024 15252 11033
rect 15936 11024 15988 11076
rect 16028 11067 16080 11076
rect 16028 11033 16037 11067
rect 16037 11033 16071 11067
rect 16071 11033 16080 11067
rect 16028 11024 16080 11033
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 17776 11092 17828 11144
rect 19800 11092 19852 11144
rect 20076 11092 20128 11144
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 19616 11024 19668 11033
rect 20352 11024 20404 11076
rect 20720 11092 20772 11144
rect 21180 11092 21232 11144
rect 23204 11092 23256 11144
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 26700 11092 26752 11144
rect 26976 11092 27028 11144
rect 20904 11024 20956 11076
rect 21088 11067 21140 11076
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 21456 11067 21508 11076
rect 21456 11033 21465 11067
rect 21465 11033 21499 11067
rect 21499 11033 21508 11067
rect 21456 11024 21508 11033
rect 24676 11024 24728 11076
rect 25136 11067 25188 11076
rect 25136 11033 25170 11067
rect 25170 11033 25188 11067
rect 25136 11024 25188 11033
rect 9680 10956 9732 11008
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 12440 10956 12492 11008
rect 12992 10956 13044 11008
rect 15844 10956 15896 11008
rect 16120 10956 16172 11008
rect 17040 10956 17092 11008
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 18328 10956 18380 11008
rect 19248 10956 19300 11008
rect 19892 10956 19944 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 1952 10795 2004 10804
rect 1952 10761 1977 10795
rect 1977 10761 2004 10795
rect 1952 10752 2004 10761
rect 3424 10752 3476 10804
rect 5264 10795 5316 10804
rect 5264 10761 5289 10795
rect 5289 10761 5316 10795
rect 5264 10752 5316 10761
rect 5540 10752 5592 10804
rect 2228 10684 2280 10736
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 3240 10684 3292 10736
rect 6000 10684 6052 10736
rect 7472 10684 7524 10736
rect 8760 10684 8812 10736
rect 5632 10616 5684 10668
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 6920 10616 6972 10668
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 8668 10616 8720 10668
rect 9680 10616 9732 10668
rect 12808 10752 12860 10804
rect 12900 10752 12952 10804
rect 15200 10752 15252 10804
rect 15292 10752 15344 10804
rect 17040 10795 17092 10804
rect 17040 10761 17065 10795
rect 17065 10761 17092 10795
rect 17040 10752 17092 10761
rect 17224 10795 17276 10804
rect 17224 10761 17233 10795
rect 17233 10761 17267 10795
rect 17267 10761 17276 10795
rect 17224 10752 17276 10761
rect 18236 10752 18288 10804
rect 10876 10684 10928 10736
rect 13544 10684 13596 10736
rect 10968 10659 11020 10668
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 12256 10616 12308 10668
rect 13636 10616 13688 10668
rect 13912 10616 13964 10668
rect 14372 10616 14424 10668
rect 2412 10548 2464 10600
rect 3424 10548 3476 10600
rect 1676 10480 1728 10532
rect 2136 10412 2188 10464
rect 4344 10412 4396 10464
rect 5448 10548 5500 10600
rect 11152 10548 11204 10600
rect 6092 10412 6144 10464
rect 7840 10412 7892 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10876 10480 10928 10532
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15384 10616 15436 10668
rect 16120 10727 16172 10736
rect 16120 10693 16145 10727
rect 16145 10693 16172 10727
rect 16120 10684 16172 10693
rect 15752 10548 15804 10600
rect 16488 10616 16540 10668
rect 16948 10684 17000 10736
rect 18144 10727 18196 10736
rect 18144 10693 18153 10727
rect 18153 10693 18187 10727
rect 18187 10693 18196 10727
rect 18144 10684 18196 10693
rect 18788 10684 18840 10736
rect 19432 10684 19484 10736
rect 19984 10727 20036 10736
rect 19984 10693 20009 10727
rect 20009 10693 20036 10727
rect 20444 10752 20496 10804
rect 22560 10752 22612 10804
rect 23664 10752 23716 10804
rect 25044 10795 25096 10804
rect 25044 10761 25053 10795
rect 25053 10761 25087 10795
rect 25087 10761 25096 10795
rect 25044 10752 25096 10761
rect 19984 10684 20036 10693
rect 19340 10616 19392 10668
rect 20536 10616 20588 10668
rect 19524 10548 19576 10600
rect 19800 10548 19852 10600
rect 20260 10548 20312 10600
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 22652 10616 22704 10668
rect 22928 10616 22980 10668
rect 21088 10548 21140 10600
rect 22100 10548 22152 10600
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 17776 10480 17828 10532
rect 23664 10591 23716 10600
rect 23664 10557 23673 10591
rect 23673 10557 23707 10591
rect 23707 10557 23716 10591
rect 23664 10548 23716 10557
rect 22560 10480 22612 10532
rect 11796 10412 11848 10464
rect 12348 10412 12400 10464
rect 15200 10412 15252 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 16948 10412 17000 10464
rect 17316 10412 17368 10464
rect 18972 10412 19024 10464
rect 19248 10412 19300 10464
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 26792 10480 26844 10532
rect 23848 10412 23900 10464
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 3976 10208 4028 10260
rect 7380 10208 7432 10260
rect 7748 10208 7800 10260
rect 8392 10208 8444 10260
rect 10048 10208 10100 10260
rect 10508 10208 10560 10260
rect 11060 10208 11112 10260
rect 11980 10208 12032 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 2136 10140 2188 10192
rect 2780 10140 2832 10192
rect 9220 10140 9272 10192
rect 9864 10140 9916 10192
rect 15292 10208 15344 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16580 10208 16632 10260
rect 17684 10208 17736 10260
rect 19248 10208 19300 10260
rect 20444 10208 20496 10260
rect 20812 10208 20864 10260
rect 17224 10140 17276 10192
rect 18788 10140 18840 10192
rect 20352 10140 20404 10192
rect 20996 10183 21048 10192
rect 20996 10149 21005 10183
rect 21005 10149 21039 10183
rect 21039 10149 21048 10183
rect 20996 10140 21048 10149
rect 21088 10140 21140 10192
rect 21548 10140 21600 10192
rect 21732 10140 21784 10192
rect 2964 10072 3016 10124
rect 480 10004 532 10056
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 3516 10004 3568 10056
rect 2412 9936 2464 9988
rect 4344 10004 4396 10056
rect 5632 10072 5684 10124
rect 6000 10072 6052 10124
rect 8208 10072 8260 10124
rect 8392 10072 8444 10124
rect 3700 9936 3752 9988
rect 5540 10004 5592 10056
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6736 10004 6788 10056
rect 6920 10004 6972 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 1584 9868 1636 9920
rect 2044 9868 2096 9920
rect 5264 9868 5316 9920
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 7196 9936 7248 9988
rect 8484 10004 8536 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9864 10004 9916 10056
rect 12440 10072 12492 10124
rect 12716 10072 12768 10124
rect 11612 10004 11664 10056
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 6828 9868 6880 9920
rect 8300 9936 8352 9988
rect 8944 9936 8996 9988
rect 10324 9936 10376 9988
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 10048 9868 10100 9920
rect 10876 9868 10928 9920
rect 11152 9936 11204 9988
rect 12164 9936 12216 9988
rect 12716 9979 12768 9988
rect 12716 9945 12725 9979
rect 12725 9945 12759 9979
rect 12759 9945 12768 9979
rect 12716 9936 12768 9945
rect 13636 10072 13688 10124
rect 16948 10072 17000 10124
rect 19248 10072 19300 10124
rect 21364 10072 21416 10124
rect 21824 10072 21876 10124
rect 22836 10072 22888 10124
rect 23204 10140 23256 10192
rect 24032 10140 24084 10192
rect 23296 10072 23348 10124
rect 13452 10004 13504 10056
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 17040 10004 17092 10056
rect 19432 10047 19484 10056
rect 16948 9936 17000 9988
rect 17224 9979 17276 9988
rect 17224 9945 17233 9979
rect 17233 9945 17267 9979
rect 17267 9945 17276 9979
rect 17224 9936 17276 9945
rect 12440 9868 12492 9920
rect 13636 9868 13688 9920
rect 15936 9868 15988 9920
rect 16856 9868 16908 9920
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 19984 10004 20036 10056
rect 22100 10004 22152 10056
rect 22192 10004 22244 10056
rect 22468 10004 22520 10056
rect 20628 9979 20680 9988
rect 20628 9945 20637 9979
rect 20637 9945 20671 9979
rect 20671 9945 20680 9979
rect 20628 9936 20680 9945
rect 19708 9868 19760 9920
rect 21548 9868 21600 9920
rect 21824 9936 21876 9988
rect 25136 10047 25188 10056
rect 25136 10013 25145 10047
rect 25145 10013 25179 10047
rect 25179 10013 25188 10047
rect 25136 10004 25188 10013
rect 26700 10004 26752 10056
rect 23940 9911 23992 9920
rect 23940 9877 23949 9911
rect 23949 9877 23983 9911
rect 23983 9877 23992 9911
rect 23940 9868 23992 9877
rect 24860 9936 24912 9988
rect 26240 9936 26292 9988
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 2964 9664 3016 9716
rect 3976 9664 4028 9716
rect 1400 9596 1452 9648
rect 2780 9596 2832 9648
rect 3240 9596 3292 9648
rect 3700 9596 3752 9648
rect 6920 9664 6972 9716
rect 8576 9664 8628 9716
rect 4988 9596 5040 9648
rect 6552 9596 6604 9648
rect 7288 9596 7340 9648
rect 9588 9664 9640 9716
rect 1676 9528 1728 9580
rect 2228 9528 2280 9580
rect 4068 9528 4120 9580
rect 3516 9460 3568 9512
rect 4344 9528 4396 9580
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 5724 9528 5776 9580
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 9404 9596 9456 9648
rect 9956 9596 10008 9648
rect 10140 9596 10192 9648
rect 10416 9596 10468 9648
rect 11612 9596 11664 9648
rect 4988 9460 5040 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 10968 9528 11020 9580
rect 11704 9528 11756 9580
rect 12164 9639 12216 9648
rect 12164 9605 12199 9639
rect 12199 9605 12216 9639
rect 12164 9596 12216 9605
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 12808 9596 12860 9648
rect 13176 9596 13228 9648
rect 14832 9664 14884 9716
rect 15476 9664 15528 9716
rect 20996 9664 21048 9716
rect 24032 9664 24084 9716
rect 24492 9664 24544 9716
rect 25136 9664 25188 9716
rect 26700 9664 26752 9716
rect 13360 9528 13412 9580
rect 14188 9596 14240 9648
rect 14280 9596 14332 9648
rect 14004 9528 14056 9580
rect 15108 9639 15160 9648
rect 15108 9605 15117 9639
rect 15117 9605 15151 9639
rect 15151 9605 15160 9639
rect 15108 9596 15160 9605
rect 15752 9528 15804 9580
rect 16488 9528 16540 9580
rect 17224 9528 17276 9580
rect 17408 9596 17460 9648
rect 17960 9528 18012 9580
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 10232 9392 10284 9444
rect 14464 9460 14516 9512
rect 14556 9460 14608 9512
rect 940 9324 992 9376
rect 3516 9324 3568 9376
rect 4068 9324 4120 9376
rect 4160 9324 4212 9376
rect 4344 9324 4396 9376
rect 4896 9324 4948 9376
rect 5080 9324 5132 9376
rect 8852 9324 8904 9376
rect 9588 9324 9640 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 13452 9392 13504 9444
rect 15108 9460 15160 9512
rect 15292 9460 15344 9512
rect 15936 9460 15988 9512
rect 18880 9596 18932 9648
rect 19800 9596 19852 9648
rect 20628 9596 20680 9648
rect 21456 9596 21508 9648
rect 22652 9596 22704 9648
rect 22744 9596 22796 9648
rect 26240 9596 26292 9648
rect 19340 9528 19392 9580
rect 21088 9528 21140 9580
rect 22284 9528 22336 9580
rect 22836 9571 22888 9580
rect 22836 9537 22845 9571
rect 22845 9537 22879 9571
rect 22879 9537 22888 9571
rect 22836 9528 22888 9537
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 23664 9528 23716 9580
rect 24492 9571 24544 9580
rect 24492 9537 24501 9571
rect 24501 9537 24535 9571
rect 24535 9537 24544 9571
rect 24492 9528 24544 9537
rect 20076 9460 20128 9512
rect 12072 9324 12124 9376
rect 12624 9324 12676 9376
rect 12900 9324 12952 9376
rect 13084 9324 13136 9376
rect 13912 9324 13964 9376
rect 15844 9392 15896 9444
rect 19708 9392 19760 9444
rect 22008 9435 22060 9444
rect 22008 9401 22017 9435
rect 22017 9401 22051 9435
rect 22051 9401 22060 9435
rect 22008 9392 22060 9401
rect 24400 9392 24452 9444
rect 26516 9571 26568 9580
rect 26516 9537 26525 9571
rect 26525 9537 26559 9571
rect 26559 9537 26568 9571
rect 26516 9528 26568 9537
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17960 9367 18012 9376
rect 17960 9333 17969 9367
rect 17969 9333 18003 9367
rect 18003 9333 18012 9367
rect 17960 9324 18012 9333
rect 20628 9324 20680 9376
rect 21272 9324 21324 9376
rect 21364 9367 21416 9376
rect 21364 9333 21373 9367
rect 21373 9333 21407 9367
rect 21407 9333 21416 9367
rect 21364 9324 21416 9333
rect 22744 9324 22796 9376
rect 23756 9324 23808 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 1768 9120 1820 9172
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3424 9120 3476 9172
rect 4712 9120 4764 9172
rect 4804 9120 4856 9172
rect 6828 9120 6880 9172
rect 7288 9120 7340 9172
rect 2688 9052 2740 9104
rect 5080 9052 5132 9104
rect 5724 9052 5776 9104
rect 1032 8916 1084 8968
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 4896 8984 4948 9036
rect 4528 8916 4580 8968
rect 7012 8984 7064 9036
rect 7748 9120 7800 9172
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 8300 9095 8352 9104
rect 8300 9061 8309 9095
rect 8309 9061 8343 9095
rect 8343 9061 8352 9095
rect 8300 9052 8352 9061
rect 8852 9052 8904 9104
rect 10140 9120 10192 9172
rect 11612 9120 11664 9172
rect 11888 9120 11940 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 12992 9163 13044 9172
rect 12992 9129 13001 9163
rect 13001 9129 13035 9163
rect 13035 9129 13044 9163
rect 12992 9120 13044 9129
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 13820 9120 13872 9172
rect 14464 9120 14516 9172
rect 14648 9120 14700 9172
rect 14740 9120 14792 9172
rect 14924 9120 14976 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 2688 8848 2740 8900
rect 2872 8848 2924 8900
rect 3608 8848 3660 8900
rect 5540 8916 5592 8968
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 10508 9052 10560 9104
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 17224 9120 17276 9172
rect 13820 8984 13872 9036
rect 15016 8984 15068 9036
rect 7656 8916 7708 8968
rect 6460 8891 6512 8900
rect 6460 8857 6469 8891
rect 6469 8857 6503 8891
rect 6503 8857 6512 8891
rect 6460 8848 6512 8857
rect 9036 8916 9088 8968
rect 10600 8916 10652 8968
rect 9404 8848 9456 8900
rect 9588 8891 9640 8900
rect 9588 8857 9597 8891
rect 9597 8857 9631 8891
rect 9631 8857 9640 8891
rect 9588 8848 9640 8857
rect 3240 8823 3292 8832
rect 3240 8789 3265 8823
rect 3265 8789 3292 8823
rect 3240 8780 3292 8789
rect 4160 8780 4212 8832
rect 4620 8780 4672 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7012 8780 7064 8832
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 8300 8780 8352 8832
rect 10784 8848 10836 8900
rect 11336 8891 11388 8900
rect 11336 8857 11345 8891
rect 11345 8857 11379 8891
rect 11379 8857 11388 8891
rect 11336 8848 11388 8857
rect 12624 8916 12676 8968
rect 13636 8916 13688 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 15476 8916 15528 8968
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 22836 9120 22888 9172
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 24768 9120 24820 9172
rect 27988 9120 28040 9172
rect 19432 8984 19484 9036
rect 10416 8780 10468 8832
rect 10600 8780 10652 8832
rect 12256 8848 12308 8900
rect 14280 8891 14332 8900
rect 14280 8857 14289 8891
rect 14289 8857 14323 8891
rect 14323 8857 14332 8891
rect 14280 8848 14332 8857
rect 18880 8916 18932 8968
rect 13176 8780 13228 8832
rect 13728 8780 13780 8832
rect 15108 8780 15160 8832
rect 19156 8848 19208 8900
rect 22376 8984 22428 9036
rect 19524 8848 19576 8900
rect 20260 8891 20312 8900
rect 20260 8857 20269 8891
rect 20269 8857 20303 8891
rect 20303 8857 20312 8891
rect 20260 8848 20312 8857
rect 20444 8891 20496 8900
rect 20444 8857 20453 8891
rect 20453 8857 20487 8891
rect 20487 8857 20496 8891
rect 20444 8848 20496 8857
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 21548 8916 21600 8968
rect 22376 8848 22428 8900
rect 16028 8780 16080 8832
rect 16304 8780 16356 8832
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 19064 8780 19116 8832
rect 20904 8780 20956 8832
rect 22468 8780 22520 8832
rect 26700 9027 26752 9036
rect 26700 8993 26709 9027
rect 26709 8993 26743 9027
rect 26743 8993 26752 9027
rect 26700 8984 26752 8993
rect 24676 8916 24728 8968
rect 26792 8916 26844 8968
rect 22744 8848 22796 8900
rect 23112 8848 23164 8900
rect 23572 8848 23624 8900
rect 24952 8780 25004 8832
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 664 8576 716 8628
rect 4344 8576 4396 8628
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 5908 8576 5960 8628
rect 1308 8508 1360 8560
rect 2320 8508 2372 8560
rect 1676 8440 1728 8492
rect 3792 8508 3844 8560
rect 5448 8508 5500 8560
rect 5540 8551 5592 8560
rect 5540 8517 5549 8551
rect 5549 8517 5583 8551
rect 5583 8517 5592 8551
rect 5540 8508 5592 8517
rect 5632 8508 5684 8560
rect 6000 8508 6052 8560
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4620 8440 4672 8492
rect 4712 8440 4764 8492
rect 4896 8440 4948 8492
rect 8484 8508 8536 8560
rect 9036 8508 9088 8560
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 11060 8576 11112 8628
rect 9404 8508 9456 8560
rect 11796 8508 11848 8560
rect 4344 8372 4396 8424
rect 5632 8372 5684 8424
rect 6184 8304 6236 8356
rect 7564 8304 7616 8356
rect 8300 8304 8352 8356
rect 8484 8304 8536 8356
rect 8852 8304 8904 8356
rect 10416 8440 10468 8492
rect 10968 8440 11020 8492
rect 14740 8576 14792 8628
rect 15568 8619 15620 8628
rect 15568 8585 15593 8619
rect 15593 8585 15620 8619
rect 15568 8576 15620 8585
rect 14188 8508 14240 8560
rect 15384 8551 15436 8560
rect 15384 8517 15393 8551
rect 15393 8517 15427 8551
rect 15427 8517 15436 8551
rect 15384 8508 15436 8517
rect 15844 8576 15896 8628
rect 16304 8576 16356 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 18144 8576 18196 8628
rect 16028 8508 16080 8560
rect 16856 8551 16908 8560
rect 16856 8517 16865 8551
rect 16865 8517 16899 8551
rect 16899 8517 16908 8551
rect 16856 8508 16908 8517
rect 17776 8508 17828 8560
rect 21916 8576 21968 8628
rect 13452 8440 13504 8492
rect 9588 8372 9640 8424
rect 10784 8372 10836 8424
rect 13636 8440 13688 8492
rect 14464 8483 14516 8492
rect 14464 8449 14471 8483
rect 14471 8449 14516 8483
rect 14464 8440 14516 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14188 8372 14240 8424
rect 15292 8440 15344 8492
rect 22100 8576 22152 8628
rect 18788 8440 18840 8492
rect 19340 8483 19392 8492
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 25228 8551 25280 8560
rect 25228 8517 25262 8551
rect 25262 8517 25280 8551
rect 25228 8508 25280 8517
rect 20628 8440 20680 8492
rect 15936 8372 15988 8424
rect 16672 8372 16724 8424
rect 17868 8372 17920 8424
rect 22284 8372 22336 8424
rect 23112 8415 23164 8424
rect 23112 8381 23121 8415
rect 23121 8381 23155 8415
rect 23155 8381 23164 8415
rect 23112 8372 23164 8381
rect 24676 8372 24728 8424
rect 13176 8304 13228 8356
rect 14464 8304 14516 8356
rect 4068 8236 4120 8288
rect 6368 8236 6420 8288
rect 7840 8236 7892 8288
rect 11152 8236 11204 8288
rect 12624 8236 12676 8288
rect 12900 8236 12952 8288
rect 13544 8236 13596 8288
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 16764 8236 16816 8288
rect 17408 8236 17460 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 19340 8304 19392 8356
rect 19800 8304 19852 8356
rect 20168 8347 20220 8356
rect 20168 8313 20177 8347
rect 20177 8313 20211 8347
rect 20211 8313 20220 8347
rect 20168 8304 20220 8313
rect 19432 8236 19484 8288
rect 19524 8236 19576 8288
rect 21088 8236 21140 8288
rect 21180 8236 21232 8288
rect 21548 8236 21600 8288
rect 26332 8347 26384 8356
rect 26332 8313 26341 8347
rect 26341 8313 26375 8347
rect 26375 8313 26384 8347
rect 26332 8304 26384 8313
rect 23480 8236 23532 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 4344 8032 4396 8084
rect 4896 8032 4948 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 2320 7828 2372 7880
rect 5632 7896 5684 7948
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5264 7828 5316 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6184 7964 6236 8016
rect 7104 8032 7156 8084
rect 8760 8032 8812 8084
rect 9128 8032 9180 8084
rect 9588 8032 9640 8084
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 10692 8032 10744 8084
rect 13636 8032 13688 8084
rect 15108 8032 15160 8084
rect 18052 8032 18104 8084
rect 18512 8032 18564 8084
rect 18788 8032 18840 8084
rect 19156 8032 19208 8084
rect 19524 8032 19576 8084
rect 20536 8032 20588 8084
rect 20720 8032 20772 8084
rect 7840 8007 7892 8016
rect 7840 7973 7849 8007
rect 7849 7973 7883 8007
rect 7883 7973 7892 8007
rect 7840 7964 7892 7973
rect 11980 7964 12032 8016
rect 6000 7828 6052 7880
rect 16028 7964 16080 8016
rect 16212 7964 16264 8016
rect 17960 7964 18012 8016
rect 21548 8032 21600 8084
rect 23112 8032 23164 8084
rect 24860 8032 24912 8084
rect 27160 8075 27212 8084
rect 27160 8041 27169 8075
rect 27169 8041 27203 8075
rect 27203 8041 27212 8075
rect 27160 8032 27212 8041
rect 28356 7964 28408 8016
rect 9404 7828 9456 7880
rect 6552 7803 6604 7812
rect 6552 7769 6561 7803
rect 6561 7769 6595 7803
rect 6595 7769 6604 7803
rect 6552 7760 6604 7769
rect 8760 7760 8812 7812
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 11152 7828 11204 7880
rect 15844 7896 15896 7948
rect 15936 7896 15988 7948
rect 5264 7692 5316 7744
rect 7380 7692 7432 7744
rect 7748 7692 7800 7744
rect 9588 7692 9640 7744
rect 11244 7692 11296 7744
rect 13084 7828 13136 7880
rect 12164 7760 12216 7812
rect 12808 7760 12860 7812
rect 14188 7828 14240 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16120 7828 16172 7880
rect 16672 7896 16724 7948
rect 16488 7828 16540 7880
rect 17132 7760 17184 7812
rect 18512 7803 18564 7812
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 13636 7692 13688 7744
rect 15844 7692 15896 7744
rect 18512 7769 18521 7803
rect 18521 7769 18555 7803
rect 18555 7769 18564 7803
rect 18512 7760 18564 7769
rect 19616 7828 19668 7880
rect 19892 7828 19944 7880
rect 19984 7828 20036 7880
rect 21548 7896 21600 7948
rect 22468 7896 22520 7948
rect 25136 7896 25188 7948
rect 22560 7828 22612 7880
rect 23848 7828 23900 7880
rect 23940 7828 23992 7880
rect 26424 7828 26476 7880
rect 18880 7692 18932 7744
rect 19432 7803 19484 7812
rect 19432 7769 19441 7803
rect 19441 7769 19475 7803
rect 19475 7769 19484 7803
rect 19432 7760 19484 7769
rect 19616 7735 19668 7744
rect 19616 7701 19641 7735
rect 19641 7701 19668 7735
rect 20628 7760 20680 7812
rect 24492 7760 24544 7812
rect 19616 7692 19668 7701
rect 21548 7692 21600 7744
rect 23204 7692 23256 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 5540 7488 5592 7540
rect 6276 7488 6328 7540
rect 7012 7488 7064 7540
rect 1676 7420 1728 7472
rect 756 7284 808 7336
rect 5264 7420 5316 7472
rect 6920 7420 6972 7472
rect 3976 7395 4028 7404
rect 3976 7361 4010 7395
rect 4010 7361 4028 7395
rect 3976 7352 4028 7361
rect 5632 7352 5684 7404
rect 4712 7216 4764 7268
rect 3700 7148 3752 7200
rect 6644 7352 6696 7404
rect 6460 7284 6512 7336
rect 6736 7216 6788 7268
rect 9036 7488 9088 7540
rect 12808 7488 12860 7540
rect 16028 7488 16080 7540
rect 16948 7488 17000 7540
rect 18144 7488 18196 7540
rect 19616 7488 19668 7540
rect 20628 7488 20680 7540
rect 20904 7488 20956 7540
rect 7288 7420 7340 7472
rect 7472 7352 7524 7404
rect 7656 7352 7708 7404
rect 8392 7352 8444 7404
rect 9680 7420 9732 7472
rect 12256 7352 12308 7404
rect 12900 7463 12952 7472
rect 12900 7429 12909 7463
rect 12909 7429 12943 7463
rect 12943 7429 12952 7463
rect 12900 7420 12952 7429
rect 14648 7420 14700 7472
rect 14832 7420 14884 7472
rect 15016 7352 15068 7404
rect 16396 7420 16448 7472
rect 17960 7420 18012 7472
rect 8116 7284 8168 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18788 7463 18840 7472
rect 18788 7429 18797 7463
rect 18797 7429 18831 7463
rect 18831 7429 18840 7463
rect 18788 7420 18840 7429
rect 19892 7420 19944 7472
rect 21732 7488 21784 7540
rect 22284 7488 22336 7540
rect 22744 7531 22796 7540
rect 22744 7497 22753 7531
rect 22753 7497 22787 7531
rect 22787 7497 22796 7531
rect 22744 7488 22796 7497
rect 18604 7352 18656 7404
rect 19156 7352 19208 7404
rect 19432 7352 19484 7404
rect 19984 7352 20036 7404
rect 20720 7395 20772 7404
rect 20720 7361 20729 7395
rect 20729 7361 20763 7395
rect 20763 7361 20772 7395
rect 20720 7352 20772 7361
rect 23480 7420 23532 7472
rect 22192 7352 22244 7404
rect 22652 7352 22704 7404
rect 23204 7352 23256 7404
rect 24676 7352 24728 7404
rect 8484 7259 8536 7268
rect 8484 7225 8493 7259
rect 8493 7225 8527 7259
rect 8527 7225 8536 7259
rect 8484 7216 8536 7225
rect 7656 7191 7708 7200
rect 7656 7157 7665 7191
rect 7665 7157 7699 7191
rect 7699 7157 7708 7191
rect 7656 7148 7708 7157
rect 8576 7148 8628 7200
rect 10508 7259 10560 7268
rect 10508 7225 10517 7259
rect 10517 7225 10551 7259
rect 10551 7225 10560 7259
rect 10508 7216 10560 7225
rect 15292 7216 15344 7268
rect 18236 7284 18288 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 9496 7148 9548 7200
rect 10416 7148 10468 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 14372 7148 14424 7200
rect 16120 7148 16172 7200
rect 18236 7148 18288 7200
rect 18604 7148 18656 7200
rect 22284 7284 22336 7336
rect 22560 7284 22612 7336
rect 23756 7284 23808 7336
rect 19984 7259 20036 7268
rect 19984 7225 19993 7259
rect 19993 7225 20027 7259
rect 20027 7225 20036 7259
rect 19984 7216 20036 7225
rect 20536 7216 20588 7268
rect 21548 7216 21600 7268
rect 20260 7148 20312 7200
rect 23572 7216 23624 7268
rect 26516 7216 26568 7268
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 4896 6944 4948 6996
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 8760 6944 8812 6996
rect 9220 6944 9272 6996
rect 9956 6944 10008 6996
rect 10508 6944 10560 6996
rect 12164 6987 12216 6996
rect 12164 6953 12173 6987
rect 12173 6953 12207 6987
rect 12207 6953 12216 6987
rect 12164 6944 12216 6953
rect 12716 6944 12768 6996
rect 13452 6944 13504 6996
rect 3240 6808 3292 6860
rect 1676 6740 1728 6792
rect 5724 6808 5776 6860
rect 10968 6876 11020 6928
rect 5264 6740 5316 6792
rect 848 6672 900 6724
rect 4804 6672 4856 6724
rect 7472 6808 7524 6860
rect 9772 6808 9824 6860
rect 7196 6740 7248 6792
rect 7748 6740 7800 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 9220 6740 9272 6792
rect 10692 6783 10744 6792
rect 10692 6749 10699 6783
rect 10699 6749 10744 6783
rect 10692 6740 10744 6749
rect 11244 6740 11296 6792
rect 8392 6672 8444 6724
rect 9312 6672 9364 6724
rect 10324 6672 10376 6724
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 12900 6876 12952 6928
rect 14004 6876 14056 6928
rect 14464 6944 14516 6996
rect 14832 6987 14884 6996
rect 14832 6953 14841 6987
rect 14841 6953 14875 6987
rect 14875 6953 14884 6987
rect 14832 6944 14884 6953
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 15016 6876 15068 6928
rect 15108 6876 15160 6928
rect 17040 6944 17092 6996
rect 17132 6944 17184 6996
rect 16488 6919 16540 6928
rect 16488 6885 16497 6919
rect 16497 6885 16531 6919
rect 16531 6885 16540 6919
rect 16488 6876 16540 6885
rect 17224 6876 17276 6928
rect 20536 6944 20588 6996
rect 20720 6944 20772 6996
rect 23112 6987 23164 6996
rect 23112 6953 23121 6987
rect 23121 6953 23155 6987
rect 23155 6953 23164 6987
rect 23112 6944 23164 6953
rect 18696 6808 18748 6860
rect 19156 6808 19208 6860
rect 19248 6808 19300 6860
rect 20628 6919 20680 6928
rect 20628 6885 20637 6919
rect 20637 6885 20671 6919
rect 20671 6885 20680 6919
rect 20628 6876 20680 6885
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 19984 6808 20036 6860
rect 21732 6851 21784 6860
rect 21732 6817 21741 6851
rect 21741 6817 21775 6851
rect 21775 6817 21784 6851
rect 21732 6808 21784 6817
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13268 6740 13320 6792
rect 13636 6740 13688 6792
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 4712 6604 4764 6656
rect 5632 6604 5684 6656
rect 6000 6604 6052 6656
rect 6368 6604 6420 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 9772 6604 9824 6656
rect 11060 6604 11112 6656
rect 13728 6672 13780 6724
rect 15108 6740 15160 6792
rect 15844 6740 15896 6792
rect 16856 6740 16908 6792
rect 15476 6715 15528 6724
rect 15476 6681 15501 6715
rect 15501 6681 15528 6715
rect 15476 6672 15528 6681
rect 16120 6715 16172 6724
rect 16120 6681 16129 6715
rect 16129 6681 16163 6715
rect 16163 6681 16172 6715
rect 16120 6672 16172 6681
rect 14372 6604 14424 6656
rect 14648 6647 14700 6656
rect 14648 6613 14673 6647
rect 14673 6613 14700 6647
rect 14648 6604 14700 6613
rect 15660 6604 15712 6656
rect 17868 6672 17920 6724
rect 16948 6604 17000 6656
rect 19340 6672 19392 6724
rect 19524 6604 19576 6656
rect 20168 6740 20220 6792
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 24676 6740 24728 6792
rect 21640 6672 21692 6724
rect 24952 6672 25004 6724
rect 25136 6672 25188 6724
rect 20720 6604 20772 6656
rect 24768 6604 24820 6656
rect 26424 6783 26476 6792
rect 26424 6749 26433 6783
rect 26433 6749 26467 6783
rect 26467 6749 26476 6783
rect 26424 6740 26476 6749
rect 26516 6740 26568 6792
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 4620 6400 4672 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 5264 6400 5316 6452
rect 5356 6400 5408 6452
rect 6368 6400 6420 6452
rect 8392 6400 8444 6452
rect 9220 6443 9272 6452
rect 9220 6409 9229 6443
rect 9229 6409 9263 6443
rect 9263 6409 9272 6443
rect 9220 6400 9272 6409
rect 9312 6400 9364 6452
rect 3700 6375 3752 6384
rect 3700 6341 3709 6375
rect 3709 6341 3743 6375
rect 3743 6341 3752 6375
rect 3700 6332 3752 6341
rect 4344 6332 4396 6384
rect 4712 6375 4764 6384
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 4988 6332 5040 6384
rect 1676 6264 1728 6316
rect 4252 6264 4304 6316
rect 2964 6196 3016 6248
rect 4896 6264 4948 6316
rect 5080 6264 5132 6316
rect 8944 6332 8996 6384
rect 9772 6332 9824 6384
rect 10048 6375 10100 6384
rect 10048 6341 10082 6375
rect 10082 6341 10100 6375
rect 10048 6332 10100 6341
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 10324 6264 10376 6316
rect 11060 6264 11112 6316
rect 11796 6307 11848 6316
rect 11796 6273 11806 6307
rect 11806 6273 11840 6307
rect 11840 6273 11848 6307
rect 12164 6400 12216 6452
rect 13360 6400 13412 6452
rect 15200 6400 15252 6452
rect 17592 6400 17644 6452
rect 17868 6400 17920 6452
rect 12440 6332 12492 6384
rect 15292 6332 15344 6384
rect 11796 6264 11848 6273
rect 6460 6196 6512 6248
rect 9128 6196 9180 6248
rect 10784 6196 10836 6248
rect 12348 6264 12400 6316
rect 13452 6264 13504 6316
rect 15200 6264 15252 6316
rect 16672 6332 16724 6384
rect 17684 6332 17736 6384
rect 18236 6375 18288 6384
rect 18236 6341 18245 6375
rect 18245 6341 18279 6375
rect 18279 6341 18288 6375
rect 18236 6332 18288 6341
rect 18972 6400 19024 6452
rect 25136 6400 25188 6452
rect 25228 6400 25280 6452
rect 19616 6332 19668 6384
rect 19984 6332 20036 6384
rect 21364 6332 21416 6384
rect 22100 6332 22152 6384
rect 22836 6332 22888 6384
rect 23388 6375 23440 6384
rect 23388 6341 23397 6375
rect 23397 6341 23431 6375
rect 23431 6341 23440 6375
rect 23388 6332 23440 6341
rect 15476 6264 15528 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16212 6264 16264 6316
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 4344 6128 4396 6180
rect 4988 6060 5040 6112
rect 5540 6060 5592 6112
rect 7196 6060 7248 6112
rect 7380 6060 7432 6112
rect 8944 6060 8996 6112
rect 10876 6128 10928 6180
rect 13636 6196 13688 6248
rect 14832 6196 14884 6248
rect 15292 6196 15344 6248
rect 16856 6196 16908 6248
rect 17132 6196 17184 6248
rect 17960 6264 18012 6316
rect 18696 6264 18748 6316
rect 19064 6307 19116 6316
rect 19064 6273 19073 6307
rect 19073 6273 19107 6307
rect 19107 6273 19116 6307
rect 19064 6264 19116 6273
rect 19248 6264 19300 6316
rect 19708 6196 19760 6248
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 22192 6264 22244 6316
rect 23204 6264 23256 6316
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 26608 6443 26660 6452
rect 26608 6409 26617 6443
rect 26617 6409 26651 6443
rect 26651 6409 26660 6443
rect 26608 6400 26660 6409
rect 21088 6196 21140 6248
rect 21272 6196 21324 6248
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 24676 6196 24728 6248
rect 25044 6196 25096 6248
rect 12716 6128 12768 6180
rect 12164 6060 12216 6112
rect 14096 6060 14148 6112
rect 14648 6128 14700 6180
rect 16212 6128 16264 6180
rect 17316 6128 17368 6180
rect 17592 6128 17644 6180
rect 18052 6128 18104 6180
rect 20628 6128 20680 6180
rect 20996 6171 21048 6180
rect 20996 6137 21005 6171
rect 21005 6137 21039 6171
rect 21039 6137 21048 6171
rect 20996 6128 21048 6137
rect 24216 6128 24268 6180
rect 14556 6060 14608 6112
rect 17868 6060 17920 6112
rect 18788 6060 18840 6112
rect 23388 6060 23440 6112
rect 23572 6060 23624 6112
rect 27068 6060 27120 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 2964 5856 3016 5908
rect 3332 5856 3384 5908
rect 1216 5788 1268 5840
rect 6736 5856 6788 5908
rect 4068 5788 4120 5840
rect 5448 5788 5500 5840
rect 9772 5856 9824 5908
rect 10048 5856 10100 5908
rect 12900 5856 12952 5908
rect 12992 5856 13044 5908
rect 572 5720 624 5772
rect 480 5652 532 5704
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 8208 5788 8260 5840
rect 8392 5788 8444 5840
rect 9128 5788 9180 5840
rect 10232 5788 10284 5840
rect 10876 5788 10928 5840
rect 17224 5856 17276 5908
rect 15752 5788 15804 5840
rect 21272 5856 21324 5908
rect 17592 5788 17644 5840
rect 20628 5788 20680 5840
rect 21088 5788 21140 5840
rect 23480 5856 23532 5908
rect 23940 5856 23992 5908
rect 24492 5856 24544 5908
rect 22744 5788 22796 5840
rect 3884 5652 3936 5704
rect 4344 5652 4396 5704
rect 7196 5720 7248 5772
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6092 5652 6144 5704
rect 7564 5652 7616 5704
rect 8760 5652 8812 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 13176 5720 13228 5772
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 14556 5720 14608 5772
rect 14832 5720 14884 5772
rect 10876 5652 10928 5704
rect 11060 5652 11112 5704
rect 2412 5627 2464 5636
rect 2412 5593 2421 5627
rect 2421 5593 2455 5627
rect 2455 5593 2464 5627
rect 2412 5584 2464 5593
rect 3792 5584 3844 5636
rect 5264 5584 5316 5636
rect 8576 5584 8628 5636
rect 9772 5584 9824 5636
rect 10600 5584 10652 5636
rect 12992 5584 13044 5636
rect 13176 5627 13228 5636
rect 13176 5593 13185 5627
rect 13185 5593 13219 5627
rect 13219 5593 13228 5627
rect 13176 5584 13228 5593
rect 13268 5627 13320 5636
rect 13268 5593 13277 5627
rect 13277 5593 13311 5627
rect 13311 5593 13320 5627
rect 13268 5584 13320 5593
rect 14096 5584 14148 5636
rect 3700 5516 3752 5568
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 7012 5516 7064 5568
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 9680 5516 9732 5568
rect 14004 5516 14056 5568
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 16212 5720 16264 5772
rect 17960 5652 18012 5704
rect 18972 5652 19024 5704
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 22928 5720 22980 5772
rect 20628 5652 20680 5704
rect 22744 5652 22796 5704
rect 23388 5652 23440 5704
rect 14280 5627 14332 5636
rect 14280 5593 14289 5627
rect 14289 5593 14323 5627
rect 14323 5593 14332 5627
rect 14280 5584 14332 5593
rect 16120 5627 16172 5636
rect 16120 5593 16129 5627
rect 16129 5593 16163 5627
rect 16163 5593 16172 5627
rect 16120 5584 16172 5593
rect 16580 5584 16632 5636
rect 16948 5584 17000 5636
rect 18420 5627 18472 5636
rect 18420 5593 18429 5627
rect 18429 5593 18463 5627
rect 18463 5593 18472 5627
rect 18420 5584 18472 5593
rect 19340 5584 19392 5636
rect 19800 5584 19852 5636
rect 22192 5584 22244 5636
rect 15476 5516 15528 5568
rect 16028 5516 16080 5568
rect 17040 5516 17092 5568
rect 20168 5516 20220 5568
rect 20536 5516 20588 5568
rect 24216 5584 24268 5636
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 26424 5720 26476 5772
rect 24676 5516 24728 5568
rect 24860 5627 24912 5636
rect 24860 5593 24894 5627
rect 24894 5593 24912 5627
rect 24860 5584 24912 5593
rect 26148 5584 26200 5636
rect 26240 5516 26292 5568
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 3792 5312 3844 5364
rect 3976 5312 4028 5364
rect 4804 5312 4856 5364
rect 5356 5312 5408 5364
rect 5448 5244 5500 5296
rect 1676 5176 1728 5228
rect 4160 5176 4212 5228
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 5908 5244 5960 5296
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 8852 5244 8904 5296
rect 9588 5244 9640 5296
rect 10784 5244 10836 5296
rect 12624 5312 12676 5364
rect 14096 5312 14148 5364
rect 13636 5244 13688 5296
rect 14832 5312 14884 5364
rect 16672 5244 16724 5296
rect 17316 5244 17368 5296
rect 17960 5287 18012 5296
rect 17960 5253 17995 5287
rect 17995 5253 18012 5287
rect 19800 5312 19852 5364
rect 17960 5244 18012 5253
rect 19340 5244 19392 5296
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 26792 5312 26844 5364
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 6092 5176 6144 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6736 5176 6788 5228
rect 9128 5176 9180 5228
rect 4988 5040 5040 5092
rect 5356 5040 5408 5092
rect 5816 5083 5868 5092
rect 5816 5049 5825 5083
rect 5825 5049 5859 5083
rect 5859 5049 5868 5083
rect 5816 5040 5868 5049
rect 6644 5040 6696 5092
rect 9128 5040 9180 5092
rect 9312 5040 9364 5092
rect 9864 5176 9916 5228
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 9772 5108 9824 5160
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 13360 5176 13412 5228
rect 15660 5176 15712 5228
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 6460 4972 6512 5024
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 14188 5108 14240 5160
rect 15476 5108 15528 5160
rect 17132 5040 17184 5092
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 20720 5176 20772 5228
rect 21640 5176 21692 5228
rect 20444 5108 20496 5160
rect 22744 5176 22796 5228
rect 24676 5219 24728 5228
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 26240 5176 26292 5228
rect 27344 5219 27396 5228
rect 27344 5185 27353 5219
rect 27353 5185 27387 5219
rect 27387 5185 27396 5219
rect 27344 5176 27396 5185
rect 25136 5108 25188 5160
rect 20076 5040 20128 5092
rect 20536 5040 20588 5092
rect 15660 4972 15712 5024
rect 16856 4972 16908 5024
rect 18420 4972 18472 5024
rect 20720 4972 20772 5024
rect 20996 4972 21048 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 388 4768 440 4820
rect 4344 4768 4396 4820
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 8576 4768 8628 4820
rect 10600 4768 10652 4820
rect 11152 4768 11204 4820
rect 17592 4768 17644 4820
rect 1676 4632 1728 4684
rect 5540 4700 5592 4752
rect 8668 4700 8720 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 15568 4700 15620 4752
rect 16396 4700 16448 4752
rect 17224 4700 17276 4752
rect 18052 4700 18104 4752
rect 3700 4632 3752 4684
rect 3884 4496 3936 4548
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 6828 4564 6880 4616
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 11152 4632 11204 4684
rect 11888 4564 11940 4616
rect 15384 4632 15436 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16948 4632 17000 4684
rect 20536 4768 20588 4820
rect 27712 4811 27764 4820
rect 27712 4777 27721 4811
rect 27721 4777 27755 4811
rect 27755 4777 27764 4811
rect 27712 4768 27764 4777
rect 12716 4564 12768 4616
rect 14372 4564 14424 4616
rect 14556 4564 14608 4616
rect 4344 4428 4396 4480
rect 7104 4496 7156 4548
rect 7748 4496 7800 4548
rect 9496 4496 9548 4548
rect 11796 4496 11848 4548
rect 12348 4496 12400 4548
rect 13728 4496 13780 4548
rect 8392 4428 8444 4480
rect 12164 4428 12216 4480
rect 12900 4428 12952 4480
rect 13820 4428 13872 4480
rect 15476 4496 15528 4548
rect 18880 4564 18932 4616
rect 19432 4564 19484 4616
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 22376 4743 22428 4752
rect 22376 4709 22385 4743
rect 22385 4709 22419 4743
rect 22419 4709 22428 4743
rect 22376 4700 22428 4709
rect 21640 4632 21692 4684
rect 23204 4607 23256 4616
rect 23204 4573 23213 4607
rect 23213 4573 23247 4607
rect 23247 4573 23256 4607
rect 23204 4564 23256 4573
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23480 4564 23532 4573
rect 25136 4632 25188 4684
rect 27252 4632 27304 4684
rect 27620 4607 27672 4616
rect 27620 4573 27629 4607
rect 27629 4573 27663 4607
rect 27663 4573 27672 4607
rect 27620 4564 27672 4573
rect 19340 4496 19392 4548
rect 14648 4471 14700 4480
rect 14648 4437 14657 4471
rect 14657 4437 14691 4471
rect 14691 4437 14700 4471
rect 14648 4428 14700 4437
rect 14740 4428 14792 4480
rect 18236 4428 18288 4480
rect 21272 4428 21324 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 3516 4156 3568 4208
rect 10140 4224 10192 4276
rect 15384 4224 15436 4276
rect 16120 4224 16172 4276
rect 1676 4088 1728 4140
rect 1124 4020 1176 4072
rect 6276 4156 6328 4208
rect 6828 4156 6880 4208
rect 4160 4088 4212 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4344 4020 4396 4072
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6460 4088 6512 4140
rect 7472 4156 7524 4208
rect 7748 4156 7800 4208
rect 12532 4156 12584 4208
rect 8760 4088 8812 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 9588 4088 9640 4140
rect 13820 4156 13872 4208
rect 14740 4156 14792 4208
rect 16856 4199 16908 4208
rect 16856 4165 16865 4199
rect 16865 4165 16899 4199
rect 16899 4165 16908 4199
rect 16856 4156 16908 4165
rect 21640 4224 21692 4276
rect 17868 4156 17920 4208
rect 2780 3952 2832 4004
rect 4252 3952 4304 4004
rect 5172 3952 5224 4004
rect 480 3884 532 3936
rect 2412 3884 2464 3936
rect 3976 3884 4028 3936
rect 5356 3884 5408 3936
rect 6736 3884 6788 3936
rect 9220 4020 9272 4072
rect 12348 4020 12400 4072
rect 16948 4088 17000 4140
rect 13268 4020 13320 4072
rect 15384 4020 15436 4072
rect 20720 4156 20772 4208
rect 24676 4224 24728 4276
rect 7012 3884 7064 3936
rect 7472 3884 7524 3936
rect 9956 3952 10008 4004
rect 10508 3995 10560 4004
rect 10508 3961 10517 3995
rect 10517 3961 10551 3995
rect 10551 3961 10560 3995
rect 10508 3952 10560 3961
rect 13912 3952 13964 4004
rect 14280 3952 14332 4004
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 15568 3884 15620 3936
rect 17776 3884 17828 3936
rect 19524 3884 19576 3936
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 21548 4088 21600 4140
rect 22192 4088 22244 4140
rect 22652 4088 22704 4140
rect 23204 4131 23256 4140
rect 23204 4097 23238 4131
rect 23238 4097 23256 4131
rect 23204 4088 23256 4097
rect 23388 4156 23440 4208
rect 25596 4156 25648 4208
rect 23480 4088 23532 4140
rect 24768 4131 24820 4140
rect 24768 4097 24777 4131
rect 24777 4097 24811 4131
rect 24811 4097 24820 4131
rect 24768 4088 24820 4097
rect 20444 3995 20496 4004
rect 20444 3961 20453 3995
rect 20453 3961 20487 3995
rect 20487 3961 20496 3995
rect 20444 3952 20496 3961
rect 22836 4020 22888 4072
rect 22284 3995 22336 4004
rect 22284 3961 22293 3995
rect 22293 3961 22327 3995
rect 22327 3961 22336 3995
rect 22284 3952 22336 3961
rect 22744 3952 22796 4004
rect 23940 4020 23992 4072
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 24216 3952 24268 4004
rect 20536 3884 20588 3936
rect 22560 3884 22612 3936
rect 26700 3884 26752 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 2504 3680 2556 3732
rect 4804 3680 4856 3732
rect 1676 3544 1728 3596
rect 5724 3612 5776 3664
rect 6552 3655 6604 3664
rect 6552 3621 6561 3655
rect 6561 3621 6595 3655
rect 6595 3621 6604 3655
rect 6552 3612 6604 3621
rect 6736 3612 6788 3664
rect 4068 3544 4120 3596
rect 5816 3544 5868 3596
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 6644 3544 6696 3596
rect 2964 3408 3016 3460
rect 4988 3408 5040 3460
rect 5080 3408 5132 3460
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6920 3476 6972 3528
rect 7288 3612 7340 3664
rect 12072 3612 12124 3664
rect 16488 3680 16540 3732
rect 16948 3723 17000 3732
rect 16948 3689 16957 3723
rect 16957 3689 16991 3723
rect 16991 3689 17000 3723
rect 16948 3680 17000 3689
rect 19340 3680 19392 3732
rect 19524 3680 19576 3732
rect 20168 3680 20220 3732
rect 12808 3612 12860 3664
rect 13084 3612 13136 3664
rect 17684 3655 17736 3664
rect 17684 3621 17693 3655
rect 17693 3621 17727 3655
rect 17727 3621 17736 3655
rect 17684 3612 17736 3621
rect 17868 3612 17920 3664
rect 19800 3655 19852 3664
rect 19800 3621 19809 3655
rect 19809 3621 19843 3655
rect 19843 3621 19852 3655
rect 19800 3612 19852 3621
rect 20628 3655 20680 3664
rect 20628 3621 20637 3655
rect 20637 3621 20671 3655
rect 20671 3621 20680 3655
rect 20628 3612 20680 3621
rect 20812 3612 20864 3664
rect 25044 3680 25096 3732
rect 8668 3544 8720 3596
rect 6644 3408 6696 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 6276 3340 6328 3392
rect 9036 3476 9088 3528
rect 9496 3476 9548 3528
rect 10140 3476 10192 3528
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 22560 3544 22612 3596
rect 24400 3544 24452 3596
rect 24768 3544 24820 3596
rect 28356 3723 28408 3732
rect 28356 3689 28365 3723
rect 28365 3689 28399 3723
rect 28399 3689 28408 3723
rect 28356 3680 28408 3689
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 13176 3476 13228 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 13728 3476 13780 3528
rect 15476 3476 15528 3528
rect 15660 3476 15712 3528
rect 18236 3476 18288 3528
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 27068 3476 27120 3528
rect 9312 3408 9364 3460
rect 10324 3408 10376 3460
rect 10416 3340 10468 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 15292 3340 15344 3392
rect 15936 3408 15988 3460
rect 20076 3408 20128 3460
rect 21548 3408 21600 3460
rect 21916 3408 21968 3460
rect 23020 3408 23072 3460
rect 24860 3408 24912 3460
rect 25044 3408 25096 3460
rect 16764 3340 16816 3392
rect 17040 3340 17092 3392
rect 19616 3340 19668 3392
rect 21364 3340 21416 3392
rect 21456 3340 21508 3392
rect 22284 3340 22336 3392
rect 24032 3340 24084 3392
rect 26516 3383 26568 3392
rect 26516 3349 26525 3383
rect 26525 3349 26559 3383
rect 26559 3349 26568 3383
rect 26516 3340 26568 3349
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 3608 3136 3660 3188
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 2136 3068 2188 3120
rect 1860 3000 1912 3052
rect 4160 3068 4212 3120
rect 4068 3000 4120 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 6552 3068 6604 3120
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 2964 2864 3016 2916
rect 2780 2796 2832 2848
rect 7472 3068 7524 3120
rect 7012 3000 7064 3052
rect 9588 3068 9640 3120
rect 9680 3068 9732 3120
rect 12716 3136 12768 3188
rect 13636 3136 13688 3188
rect 14372 3136 14424 3188
rect 17408 3136 17460 3188
rect 20260 3136 20312 3188
rect 20444 3136 20496 3188
rect 21732 3136 21784 3188
rect 26516 3136 26568 3188
rect 10600 3000 10652 3052
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 15476 3068 15528 3120
rect 15660 3068 15712 3120
rect 16856 3068 16908 3120
rect 17316 3111 17368 3120
rect 17316 3077 17325 3111
rect 17325 3077 17359 3111
rect 17359 3077 17368 3111
rect 17316 3068 17368 3077
rect 20904 3068 20956 3120
rect 21548 3068 21600 3120
rect 24124 3068 24176 3120
rect 13268 3000 13320 3052
rect 11244 2932 11296 2984
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 15476 2932 15528 2984
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 21916 3000 21968 3052
rect 17592 2932 17644 2984
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 4988 2796 5040 2848
rect 6736 2796 6788 2848
rect 9772 2864 9824 2916
rect 12532 2864 12584 2916
rect 9496 2796 9548 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 13544 2796 13596 2848
rect 17960 2864 18012 2916
rect 20260 2864 20312 2916
rect 21732 2864 21784 2916
rect 23388 2907 23440 2916
rect 23388 2873 23397 2907
rect 23397 2873 23431 2907
rect 23431 2873 23440 2907
rect 23388 2864 23440 2873
rect 15844 2796 15896 2848
rect 22284 2796 22336 2848
rect 22652 2796 22704 2848
rect 24400 2975 24452 2984
rect 24400 2941 24409 2975
rect 24409 2941 24443 2975
rect 24443 2941 24452 2975
rect 24400 2932 24452 2941
rect 25780 2907 25832 2916
rect 25780 2873 25789 2907
rect 25789 2873 25823 2907
rect 25823 2873 25832 2907
rect 25780 2864 25832 2873
rect 26240 2907 26292 2916
rect 26240 2873 26249 2907
rect 26249 2873 26283 2907
rect 26283 2873 26292 2907
rect 26240 2864 26292 2873
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 6552 2592 6604 2644
rect 4712 2567 4764 2576
rect 4712 2533 4721 2567
rect 4721 2533 4755 2567
rect 4755 2533 4764 2567
rect 4712 2524 4764 2533
rect 7380 2592 7432 2644
rect 9956 2592 10008 2644
rect 10508 2592 10560 2644
rect 11244 2592 11296 2644
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 15384 2592 15436 2644
rect 16396 2592 16448 2644
rect 17408 2592 17460 2644
rect 17684 2592 17736 2644
rect 21180 2592 21232 2644
rect 12624 2524 12676 2576
rect 13268 2524 13320 2576
rect 15476 2524 15528 2576
rect 17500 2524 17552 2576
rect 18696 2524 18748 2576
rect 19432 2567 19484 2576
rect 19432 2533 19441 2567
rect 19441 2533 19475 2567
rect 19475 2533 19484 2567
rect 19432 2524 19484 2533
rect 21640 2524 21692 2576
rect 25688 2592 25740 2644
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 1676 2388 1728 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 7012 2388 7064 2440
rect 10968 2456 11020 2508
rect 7196 2320 7248 2372
rect 8208 2388 8260 2440
rect 9680 2388 9732 2440
rect 10140 2388 10192 2440
rect 11244 2388 11296 2440
rect 15200 2456 15252 2508
rect 17868 2456 17920 2508
rect 20444 2456 20496 2508
rect 22100 2456 22152 2508
rect 22560 2456 22612 2508
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 14648 2388 14700 2440
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 15476 2388 15528 2440
rect 15568 2388 15620 2440
rect 17408 2388 17460 2440
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18144 2388 18196 2440
rect 18604 2388 18656 2440
rect 18880 2388 18932 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19708 2388 19760 2440
rect 20168 2388 20220 2440
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 21640 2388 21692 2440
rect 23388 2388 23440 2440
rect 24400 2388 24452 2440
rect 26792 2388 26844 2440
rect 9220 2320 9272 2372
rect 15200 2320 15252 2372
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 8392 2252 8444 2304
rect 11704 2252 11756 2304
rect 17500 2252 17552 2304
rect 21272 2320 21324 2372
rect 24952 2320 25004 2372
rect 20444 2252 20496 2304
rect 22376 2252 22428 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 3516 2091 3568 2100
rect 3516 2057 3525 2091
rect 3525 2057 3559 2091
rect 3559 2057 3568 2091
rect 3516 2048 3568 2057
rect 4160 2048 4212 2100
rect 7104 2048 7156 2100
rect 9128 2048 9180 2100
rect 11152 2091 11204 2100
rect 11152 2057 11161 2091
rect 11161 2057 11195 2091
rect 11195 2057 11204 2091
rect 11152 2048 11204 2057
rect 2596 1980 2648 2032
rect 6644 1980 6696 2032
rect 7656 1980 7708 2032
rect 9496 1980 9548 2032
rect 12348 2023 12400 2032
rect 12348 1989 12357 2023
rect 12357 1989 12391 2023
rect 12391 1989 12400 2023
rect 12348 1980 12400 1989
rect 5264 1912 5316 1964
rect 6000 1955 6052 1964
rect 6000 1921 6009 1955
rect 6009 1921 6043 1955
rect 6043 1921 6052 1955
rect 6000 1912 6052 1921
rect 6552 1912 6604 1964
rect 7104 1912 7156 1964
rect 8944 1912 8996 1964
rect 9680 1912 9732 1964
rect 10968 1912 11020 1964
rect 12532 1980 12584 2032
rect 14464 1980 14516 2032
rect 15936 1980 15988 2032
rect 16488 1980 16540 2032
rect 17500 1980 17552 2032
rect 4712 1708 4764 1760
rect 13268 1955 13320 1964
rect 13268 1921 13277 1955
rect 13277 1921 13311 1955
rect 13311 1921 13320 1955
rect 13268 1912 13320 1921
rect 17408 1912 17460 1964
rect 17684 1912 17736 1964
rect 18604 1912 18656 1964
rect 7380 1819 7432 1828
rect 7380 1785 7389 1819
rect 7389 1785 7423 1819
rect 7423 1785 7432 1819
rect 7380 1776 7432 1785
rect 12256 1776 12308 1828
rect 12716 1819 12768 1828
rect 12716 1785 12725 1819
rect 12725 1785 12759 1819
rect 12759 1785 12768 1819
rect 12716 1776 12768 1785
rect 14280 1776 14332 1828
rect 15568 1819 15620 1828
rect 15568 1785 15577 1819
rect 15577 1785 15611 1819
rect 15611 1785 15620 1819
rect 15568 1776 15620 1785
rect 17868 1776 17920 1828
rect 15108 1708 15160 1760
rect 17224 1708 17276 1760
rect 17960 1708 18012 1760
rect 22560 1980 22612 2032
rect 23848 1980 23900 2032
rect 20904 1912 20956 1964
rect 21364 1955 21416 1964
rect 21364 1921 21373 1955
rect 21373 1921 21407 1955
rect 21407 1921 21416 1955
rect 21364 1912 21416 1921
rect 21548 1912 21600 1964
rect 26332 2091 26384 2100
rect 26332 2057 26341 2091
rect 26341 2057 26375 2091
rect 26375 2057 26384 2091
rect 26332 2048 26384 2057
rect 26516 1955 26568 1964
rect 26516 1921 26525 1955
rect 26525 1921 26559 1955
rect 26559 1921 26568 1955
rect 26516 1912 26568 1921
rect 20628 1844 20680 1896
rect 23848 1887 23900 1896
rect 23848 1853 23857 1887
rect 23857 1853 23891 1887
rect 23891 1853 23900 1887
rect 23848 1844 23900 1853
rect 21640 1776 21692 1828
rect 23388 1819 23440 1828
rect 23388 1785 23397 1819
rect 23397 1785 23431 1819
rect 23431 1785 23440 1819
rect 23388 1776 23440 1785
rect 25688 1819 25740 1828
rect 25688 1785 25697 1819
rect 25697 1785 25731 1819
rect 25731 1785 25740 1819
rect 25688 1776 25740 1785
rect 22652 1708 22704 1760
rect 23480 1708 23532 1760
rect 4423 1606 4475 1658
rect 4487 1606 4539 1658
rect 4551 1606 4603 1658
rect 4615 1606 4667 1658
rect 4679 1606 4731 1658
rect 11369 1606 11421 1658
rect 11433 1606 11485 1658
rect 11497 1606 11549 1658
rect 11561 1606 11613 1658
rect 11625 1606 11677 1658
rect 18315 1606 18367 1658
rect 18379 1606 18431 1658
rect 18443 1606 18495 1658
rect 18507 1606 18559 1658
rect 18571 1606 18623 1658
rect 25261 1606 25313 1658
rect 25325 1606 25377 1658
rect 25389 1606 25441 1658
rect 25453 1606 25505 1658
rect 25517 1606 25569 1658
rect 6368 1504 6420 1556
rect 9772 1479 9824 1488
rect 9772 1445 9781 1479
rect 9781 1445 9815 1479
rect 9815 1445 9824 1479
rect 9772 1436 9824 1445
rect 14556 1436 14608 1488
rect 17316 1436 17368 1488
rect 1584 1411 1636 1420
rect 1584 1377 1593 1411
rect 1593 1377 1627 1411
rect 1627 1377 1636 1411
rect 1584 1368 1636 1377
rect 4160 1411 4212 1420
rect 4160 1377 4169 1411
rect 4169 1377 4203 1411
rect 4203 1377 4212 1411
rect 4160 1368 4212 1377
rect 2780 1300 2832 1352
rect 6736 1300 6788 1352
rect 10324 1300 10376 1352
rect 8208 1232 8260 1284
rect 10692 1300 10744 1352
rect 11060 1300 11112 1352
rect 11244 1368 11296 1420
rect 11796 1300 11848 1352
rect 5816 1164 5868 1216
rect 5908 1207 5960 1216
rect 5908 1173 5917 1207
rect 5917 1173 5951 1207
rect 5951 1173 5960 1207
rect 5908 1164 5960 1173
rect 7748 1164 7800 1216
rect 9956 1207 10008 1216
rect 9956 1173 9965 1207
rect 9965 1173 9999 1207
rect 9999 1173 10008 1207
rect 9956 1164 10008 1173
rect 10876 1232 10928 1284
rect 14464 1411 14516 1420
rect 14464 1377 14473 1411
rect 14473 1377 14507 1411
rect 14507 1377 14516 1411
rect 14464 1368 14516 1377
rect 15200 1300 15252 1352
rect 15660 1368 15712 1420
rect 18144 1504 18196 1556
rect 18696 1504 18748 1556
rect 23480 1504 23532 1556
rect 15844 1300 15896 1352
rect 17040 1343 17092 1352
rect 17040 1309 17049 1343
rect 17049 1309 17083 1343
rect 17083 1309 17092 1343
rect 17040 1300 17092 1309
rect 17408 1300 17460 1352
rect 17592 1300 17644 1352
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 23848 1368 23900 1420
rect 15108 1164 15160 1216
rect 21456 1343 21508 1352
rect 21456 1309 21465 1343
rect 21465 1309 21499 1343
rect 21499 1309 21508 1343
rect 21456 1300 21508 1309
rect 22560 1300 22612 1352
rect 18880 1207 18932 1216
rect 18880 1173 18889 1207
rect 18889 1173 18923 1207
rect 18923 1173 18932 1207
rect 18880 1164 18932 1173
rect 20812 1207 20864 1216
rect 20812 1173 20821 1207
rect 20821 1173 20855 1207
rect 20855 1173 20864 1207
rect 20812 1164 20864 1173
rect 23204 1232 23256 1284
rect 23388 1207 23440 1216
rect 23388 1173 23397 1207
rect 23397 1173 23431 1207
rect 23431 1173 23440 1207
rect 23388 1164 23440 1173
rect 24032 1343 24084 1352
rect 24032 1309 24041 1343
rect 24041 1309 24075 1343
rect 24075 1309 24084 1343
rect 24032 1300 24084 1309
rect 24860 1343 24912 1352
rect 24860 1309 24894 1343
rect 24894 1309 24912 1343
rect 24860 1300 24912 1309
rect 26608 1343 26660 1352
rect 26608 1309 26617 1343
rect 26617 1309 26651 1343
rect 26651 1309 26660 1343
rect 26608 1300 26660 1309
rect 27344 1343 27396 1352
rect 27344 1309 27353 1343
rect 27353 1309 27387 1343
rect 27387 1309 27396 1343
rect 27344 1300 27396 1309
rect 25044 1164 25096 1216
rect 25596 1164 25648 1216
rect 26424 1207 26476 1216
rect 26424 1173 26433 1207
rect 26433 1173 26467 1207
rect 26467 1173 26476 1207
rect 26424 1164 26476 1173
rect 27160 1207 27212 1216
rect 27160 1173 27169 1207
rect 27169 1173 27203 1207
rect 27203 1173 27212 1207
rect 27160 1164 27212 1173
rect 7896 1062 7948 1114
rect 7960 1062 8012 1114
rect 8024 1062 8076 1114
rect 8088 1062 8140 1114
rect 8152 1062 8204 1114
rect 14842 1062 14894 1114
rect 14906 1062 14958 1114
rect 14970 1062 15022 1114
rect 15034 1062 15086 1114
rect 15098 1062 15150 1114
rect 21788 1062 21840 1114
rect 21852 1062 21904 1114
rect 21916 1062 21968 1114
rect 21980 1062 22032 1114
rect 22044 1062 22096 1114
rect 28734 1062 28786 1114
rect 28798 1062 28850 1114
rect 28862 1062 28914 1114
rect 28926 1062 28978 1114
rect 28990 1062 29042 1114
rect 10968 960 11020 1012
rect 26424 960 26476 1012
rect 9956 892 10008 944
rect 26608 892 26660 944
rect 4068 824 4120 876
rect 27160 824 27212 876
rect 5908 756 5960 808
rect 26700 756 26752 808
rect 16764 688 16816 740
rect 20812 688 20864 740
rect 3976 620 4028 672
rect 15568 552 15620 604
rect 18880 552 18932 604
rect 19064 552 19116 604
rect 23388 688 23440 740
rect 27344 620 27396 672
<< metal2 >>
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 12808 33584 12860 33590
rect 12808 33526 12860 33532
rect 9220 33516 9272 33522
rect 9220 33458 9272 33464
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 2332 32570 2360 32846
rect 2320 32564 2372 32570
rect 2320 32506 2372 32512
rect 3332 32496 3384 32502
rect 3332 32438 3384 32444
rect 2872 32428 2924 32434
rect 2872 32370 2924 32376
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 2688 32360 2740 32366
rect 2688 32302 2740 32308
rect 1584 31136 1636 31142
rect 1584 31078 1636 31084
rect 1596 30734 1624 31078
rect 2424 30734 2452 32302
rect 2700 31890 2728 32302
rect 2884 32230 2912 32370
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 2872 32224 2924 32230
rect 2872 32166 2924 32172
rect 2884 31890 2912 32166
rect 2596 31884 2648 31890
rect 2596 31826 2648 31832
rect 2688 31884 2740 31890
rect 2688 31826 2740 31832
rect 2872 31884 2924 31890
rect 2872 31826 2924 31832
rect 2502 31376 2558 31385
rect 2502 31311 2504 31320
rect 2556 31311 2558 31320
rect 2504 31282 2556 31288
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 2412 30728 2464 30734
rect 2412 30670 2464 30676
rect 2136 30320 2188 30326
rect 2134 30288 2136 30297
rect 2188 30288 2190 30297
rect 1952 30252 2004 30258
rect 1952 30194 2004 30200
rect 2044 30252 2096 30258
rect 2134 30223 2190 30232
rect 2320 30252 2372 30258
rect 2044 30194 2096 30200
rect 2320 30194 2372 30200
rect 1860 30048 1912 30054
rect 1860 29990 1912 29996
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 478 28248 534 28257
rect 478 28183 534 28192
rect 492 27674 520 28183
rect 480 27668 532 27674
rect 480 27610 532 27616
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 1412 24818 1440 25774
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 480 23588 532 23594
rect 480 23530 532 23536
rect 492 22137 520 23530
rect 1308 23044 1360 23050
rect 1308 22986 1360 22992
rect 478 22128 534 22137
rect 478 22063 534 22072
rect 572 21956 624 21962
rect 572 21898 624 21904
rect 480 21480 532 21486
rect 480 21422 532 21428
rect 492 20097 520 21422
rect 478 20088 534 20097
rect 478 20023 534 20032
rect 584 18057 612 21898
rect 938 20904 994 20913
rect 938 20839 994 20848
rect 848 19712 900 19718
rect 848 19654 900 19660
rect 570 18048 626 18057
rect 570 17983 626 17992
rect 478 16008 534 16017
rect 478 15943 534 15952
rect 492 15502 520 15943
rect 480 15496 532 15502
rect 480 15438 532 15444
rect 478 13968 534 13977
rect 478 13903 534 13912
rect 492 12434 520 13903
rect 754 12744 810 12753
rect 754 12679 810 12688
rect 492 12406 612 12434
rect 388 11892 440 11898
rect 388 11834 440 11840
rect 400 4826 428 11834
rect 480 10056 532 10062
rect 480 9998 532 10004
rect 492 9897 520 9998
rect 478 9888 534 9897
rect 478 9823 534 9832
rect 478 5808 534 5817
rect 584 5778 612 12406
rect 664 11688 716 11694
rect 664 11630 716 11636
rect 676 8634 704 11630
rect 664 8628 716 8634
rect 664 8570 716 8576
rect 768 7342 796 12679
rect 756 7336 808 7342
rect 756 7278 808 7284
rect 860 6730 888 19654
rect 952 11898 980 20839
rect 1320 20602 1348 22986
rect 1308 20596 1360 20602
rect 1308 20538 1360 20544
rect 1124 20392 1176 20398
rect 1124 20334 1176 20340
rect 1032 17876 1084 17882
rect 1032 17818 1084 17824
rect 940 11892 992 11898
rect 940 11834 992 11840
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 9382 980 11698
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 1044 8974 1072 17818
rect 1136 11762 1164 20334
rect 1308 18080 1360 18086
rect 1308 18022 1360 18028
rect 1216 15700 1268 15706
rect 1216 15642 1268 15648
rect 1124 11756 1176 11762
rect 1124 11698 1176 11704
rect 1228 11694 1256 15642
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1124 11620 1176 11626
rect 1124 11562 1176 11568
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 848 6724 900 6730
rect 848 6666 900 6672
rect 478 5743 534 5752
rect 572 5772 624 5778
rect 492 5710 520 5743
rect 572 5714 624 5720
rect 480 5704 532 5710
rect 480 5646 532 5652
rect 388 4820 440 4826
rect 388 4762 440 4768
rect 1136 4078 1164 11562
rect 1216 11552 1268 11558
rect 1216 11494 1268 11500
rect 1228 5846 1256 11494
rect 1320 8566 1348 18022
rect 1412 16289 1440 24754
rect 1504 22098 1532 29446
rect 1872 28558 1900 29990
rect 1964 29578 1992 30194
rect 1952 29572 2004 29578
rect 1952 29514 2004 29520
rect 2056 29510 2084 30194
rect 2044 29504 2096 29510
rect 2044 29446 2096 29452
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1964 28082 1992 28358
rect 2332 28218 2360 30194
rect 2412 29640 2464 29646
rect 2410 29608 2412 29617
rect 2464 29608 2466 29617
rect 2410 29543 2466 29552
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 1780 27402 1808 28018
rect 1964 27470 1992 28018
rect 2044 28008 2096 28014
rect 2044 27950 2096 27956
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1780 26994 1808 27338
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1780 26382 1808 26930
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 1688 25770 1716 26250
rect 1780 26234 1808 26318
rect 1780 26206 1900 26234
rect 1872 25838 1900 26206
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1676 25764 1728 25770
rect 1676 25706 1728 25712
rect 1964 25294 1992 27406
rect 2056 25294 2084 27950
rect 2412 27396 2464 27402
rect 2412 27338 2464 27344
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1872 24954 1900 25162
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 1964 24834 1992 25230
rect 1860 24812 1912 24818
rect 1964 24806 2084 24834
rect 1860 24754 1912 24760
rect 1768 23792 1820 23798
rect 1766 23760 1768 23769
rect 1820 23760 1822 23769
rect 1766 23695 1822 23704
rect 1872 23322 1900 24754
rect 2056 24750 2084 24806
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 2056 24206 2084 24686
rect 2148 24206 2176 26862
rect 2424 26042 2452 27338
rect 2516 27062 2544 31078
rect 2608 29306 2636 31826
rect 3068 31754 3096 32302
rect 3148 32224 3200 32230
rect 3148 32166 3200 32172
rect 3056 31748 3108 31754
rect 3056 31690 3108 31696
rect 3068 31278 3096 31690
rect 3160 31482 3188 32166
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3252 31210 3280 32302
rect 3344 32026 3372 32438
rect 4816 32366 4844 33254
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 4804 32360 4856 32366
rect 3422 32328 3478 32337
rect 4804 32302 4856 32308
rect 3422 32263 3478 32272
rect 4252 32292 4304 32298
rect 3436 32026 3464 32263
rect 4304 32252 4384 32280
rect 4252 32234 4304 32240
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 3424 32020 3476 32026
rect 3424 31962 3476 31968
rect 4356 31958 4384 32252
rect 4423 32124 4731 32133
rect 4423 32122 4429 32124
rect 4485 32122 4509 32124
rect 4565 32122 4589 32124
rect 4645 32122 4669 32124
rect 4725 32122 4731 32124
rect 4485 32070 4487 32122
rect 4667 32070 4669 32122
rect 4423 32068 4429 32070
rect 4485 32068 4509 32070
rect 4565 32068 4589 32070
rect 4645 32068 4669 32070
rect 4725 32068 4731 32070
rect 4423 32059 4731 32068
rect 4252 31952 4304 31958
rect 4252 31894 4304 31900
rect 4344 31952 4396 31958
rect 4344 31894 4396 31900
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 4160 31816 4212 31822
rect 4160 31758 4212 31764
rect 3240 31204 3292 31210
rect 3240 31146 3292 31152
rect 2778 30696 2834 30705
rect 2778 30631 2834 30640
rect 2792 29850 2820 30631
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2596 29300 2648 29306
rect 2596 29242 2648 29248
rect 2884 27130 2912 30194
rect 3252 29782 3280 31146
rect 3884 30864 3936 30870
rect 3330 30832 3386 30841
rect 3884 30806 3936 30812
rect 3330 30767 3332 30776
rect 3384 30767 3386 30776
rect 3332 30738 3384 30744
rect 3240 29776 3292 29782
rect 3240 29718 3292 29724
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3160 28422 3188 29650
rect 3792 29232 3844 29238
rect 3792 29174 3844 29180
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3148 28416 3200 28422
rect 3148 28358 3200 28364
rect 3160 28218 3188 28358
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2504 27056 2556 27062
rect 2504 26998 2556 27004
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2226 25120 2282 25129
rect 2226 25055 2282 25064
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1504 21865 1532 22034
rect 1780 22030 1808 22714
rect 1872 22250 1900 23054
rect 2056 22574 2084 24142
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2148 22642 2176 23666
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2134 22264 2190 22273
rect 1872 22222 2084 22250
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1872 22030 1900 22063
rect 1768 22024 1820 22030
rect 1768 21966 1820 21972
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1490 21856 1546 21865
rect 1490 21791 1546 21800
rect 1504 20262 1532 21791
rect 1780 21622 1808 21966
rect 1768 21616 1820 21622
rect 1768 21558 1820 21564
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 20942 1716 21286
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16590 1624 16934
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1398 16280 1454 16289
rect 1398 16215 1454 16224
rect 1596 14074 1624 16526
rect 1688 15094 1716 20402
rect 1780 19310 1808 21422
rect 1952 21412 2004 21418
rect 1952 21354 2004 21360
rect 1964 19854 1992 21354
rect 2056 21078 2084 22222
rect 2134 22199 2190 22208
rect 2148 22030 2176 22199
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2240 21894 2268 25055
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2332 21842 2360 25774
rect 2596 25764 2648 25770
rect 2596 25706 2648 25712
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24750 2544 25230
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2608 23798 2636 25706
rect 2976 24886 3004 25774
rect 2964 24880 3016 24886
rect 2964 24822 3016 24828
rect 2976 23866 3004 24822
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2412 23248 2464 23254
rect 2412 23190 2464 23196
rect 2424 22438 2452 23190
rect 2976 23186 3004 23802
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2962 23080 3018 23089
rect 2962 23015 2964 23024
rect 3016 23015 3018 23024
rect 2964 22986 3016 22992
rect 3068 22982 3096 24006
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2240 21554 2268 21830
rect 2332 21814 2452 21842
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 2056 20942 2084 21014
rect 2044 20936 2096 20942
rect 2424 20913 2452 21814
rect 2516 21593 2544 22918
rect 2686 22808 2742 22817
rect 2686 22743 2688 22752
rect 2740 22743 2742 22752
rect 2688 22714 2740 22720
rect 2594 22536 2650 22545
rect 2594 22471 2650 22480
rect 2502 21584 2558 21593
rect 2502 21519 2504 21528
rect 2556 21519 2558 21528
rect 2504 21490 2556 21496
rect 2608 21146 2636 22471
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2884 22234 2912 22374
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 2870 22128 2926 22137
rect 3068 22094 3096 22918
rect 3252 22760 3280 28494
rect 3700 27940 3752 27946
rect 3700 27882 3752 27888
rect 3608 27668 3660 27674
rect 3608 27610 3660 27616
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3344 24698 3372 27270
rect 3516 26920 3568 26926
rect 3516 26862 3568 26868
rect 3424 25968 3476 25974
rect 3422 25936 3424 25945
rect 3476 25936 3478 25945
rect 3422 25871 3478 25880
rect 3344 24670 3464 24698
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 2870 22063 2926 22072
rect 2976 22066 3096 22094
rect 3160 22732 3280 22760
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2778 21992 2834 22001
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2044 20878 2096 20884
rect 2410 20904 2466 20913
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1768 18760 1820 18766
rect 1872 18748 1900 19722
rect 1952 19372 2004 19378
rect 2056 19360 2084 20878
rect 2228 20868 2280 20874
rect 2410 20839 2466 20848
rect 2228 20810 2280 20816
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2148 20369 2176 20402
rect 2134 20360 2190 20369
rect 2134 20295 2190 20304
rect 2240 20233 2268 20810
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2226 20224 2282 20233
rect 2226 20159 2282 20168
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2004 19332 2084 19360
rect 1952 19314 2004 19320
rect 2044 19236 2096 19242
rect 2044 19178 2096 19184
rect 1820 18720 1900 18748
rect 1768 18702 1820 18708
rect 1780 16794 1808 18702
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1872 17610 1900 18566
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 1780 14249 1808 16050
rect 1872 15162 1900 17546
rect 2056 17320 2084 19178
rect 2240 18834 2268 19654
rect 2332 19378 2360 20742
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2424 19553 2452 20538
rect 2502 20496 2558 20505
rect 2502 20431 2558 20440
rect 2410 19544 2466 19553
rect 2516 19514 2544 20431
rect 2596 19984 2648 19990
rect 2700 19972 2728 21966
rect 2778 21927 2834 21936
rect 2648 19944 2728 19972
rect 2596 19926 2648 19932
rect 2792 19904 2820 21927
rect 2884 20806 2912 22063
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2884 19961 2912 20470
rect 2700 19876 2820 19904
rect 2870 19952 2926 19961
rect 2870 19887 2926 19896
rect 2410 19479 2466 19488
rect 2504 19508 2556 19514
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2134 18456 2190 18465
rect 2134 18391 2136 18400
rect 2188 18391 2190 18400
rect 2136 18362 2188 18368
rect 2424 18290 2452 19479
rect 2504 19450 2556 19456
rect 2700 19378 2728 19876
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2792 19514 2820 19722
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2608 18766 2636 19246
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2608 17678 2636 18702
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2228 17332 2280 17338
rect 2056 17292 2176 17320
rect 2148 17202 2176 17292
rect 2228 17274 2280 17280
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16726 1992 17070
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1964 15026 1992 16662
rect 2056 15026 2084 17138
rect 2240 16590 2268 17274
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2148 15706 2176 15982
rect 2240 15706 2268 16526
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2332 15026 2360 17138
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2134 14512 2190 14521
rect 2134 14447 2190 14456
rect 2148 14414 2176 14447
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1766 14240 1822 14249
rect 1766 14175 1822 14184
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 10538 1716 13262
rect 1872 12986 1900 14350
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1950 13968 2006 13977
rect 1950 13903 2006 13912
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1964 12288 1992 13903
rect 2056 13530 2084 14214
rect 2332 14074 2360 14962
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2332 12345 2360 12786
rect 1872 12260 1992 12288
rect 2318 12336 2374 12345
rect 2424 12306 2452 17546
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 16522 2544 17138
rect 2608 16522 2636 17614
rect 2700 17338 2728 18226
rect 2792 17882 2820 18634
rect 2884 18630 2912 19790
rect 2976 19174 3004 22066
rect 3054 21992 3110 22001
rect 3054 21927 3110 21936
rect 3068 21894 3096 21927
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3054 21584 3110 21593
rect 3054 21519 3056 21528
rect 3108 21519 3110 21528
rect 3056 21490 3108 21496
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3068 18850 3096 20946
rect 3160 20505 3188 22732
rect 3238 22672 3294 22681
rect 3238 22607 3240 22616
rect 3292 22607 3294 22616
rect 3240 22578 3292 22584
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 22273 3280 22374
rect 3238 22264 3294 22273
rect 3238 22199 3294 22208
rect 3240 21956 3292 21962
rect 3240 21898 3292 21904
rect 3252 21078 3280 21898
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3252 20942 3280 21014
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3146 20496 3202 20505
rect 3146 20431 3202 20440
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 19514 3188 20198
rect 3252 19514 3280 20402
rect 3344 19854 3372 24550
rect 3436 23848 3464 24670
rect 3528 24410 3556 26862
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3436 23820 3556 23848
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3436 21146 3464 23666
rect 3528 22438 3556 23820
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3620 21690 3648 27610
rect 3712 25906 3740 27882
rect 3804 26586 3832 29174
rect 3896 28626 3924 30806
rect 3988 30394 4016 31758
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4066 30152 4122 30161
rect 4066 30087 4122 30096
rect 4080 29850 4108 30087
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 4172 29646 4200 31758
rect 4264 30598 4292 31894
rect 4344 31680 4396 31686
rect 4344 31622 4396 31628
rect 4528 31680 4580 31686
rect 4528 31622 4580 31628
rect 4356 31142 4384 31622
rect 4540 31482 4568 31622
rect 4528 31476 4580 31482
rect 4528 31418 4580 31424
rect 4816 31346 4844 32302
rect 5184 32298 5212 32506
rect 6644 32360 6696 32366
rect 6644 32302 6696 32308
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5184 31686 5212 32234
rect 5264 31952 5316 31958
rect 5262 31920 5264 31929
rect 5316 31920 5318 31929
rect 5262 31855 5318 31864
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5184 31482 5212 31622
rect 5172 31476 5224 31482
rect 5172 31418 5224 31424
rect 5184 31346 5212 31418
rect 4804 31340 4856 31346
rect 4804 31282 4856 31288
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 4344 31136 4396 31142
rect 4344 31078 4396 31084
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 4344 30660 4396 30666
rect 4344 30602 4396 30608
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 4160 29640 4212 29646
rect 4160 29582 4212 29588
rect 3976 29232 4028 29238
rect 3976 29174 4028 29180
rect 3884 28620 3936 28626
rect 3884 28562 3936 28568
rect 3884 28144 3936 28150
rect 3884 28086 3936 28092
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3790 26208 3846 26217
rect 3790 26143 3846 26152
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3700 23180 3752 23186
rect 3700 23122 3752 23128
rect 3712 22778 3740 23122
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3700 22636 3752 22642
rect 3700 22578 3752 22584
rect 3712 22234 3740 22578
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3804 22098 3832 26143
rect 3896 24800 3924 28086
rect 3988 27606 4016 29174
rect 4160 29028 4212 29034
rect 4160 28970 4212 28976
rect 4172 28665 4200 28970
rect 4158 28656 4214 28665
rect 4158 28591 4214 28600
rect 4356 28529 4384 30602
rect 5184 30598 5212 31282
rect 5736 31278 5764 31758
rect 6104 31346 6132 31758
rect 6092 31340 6144 31346
rect 6092 31282 6144 31288
rect 5724 31272 5776 31278
rect 5724 31214 5776 31220
rect 5736 30734 5764 31214
rect 6104 30870 6132 31282
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6092 30864 6144 30870
rect 6092 30806 6144 30812
rect 5724 30728 5776 30734
rect 5724 30670 5776 30676
rect 5172 30592 5224 30598
rect 5172 30534 5224 30540
rect 4896 30252 4948 30258
rect 4896 30194 4948 30200
rect 4804 30184 4856 30190
rect 4804 30126 4856 30132
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4710 29200 4766 29209
rect 4816 29170 4844 30126
rect 4710 29135 4766 29144
rect 4804 29164 4856 29170
rect 4724 29102 4752 29135
rect 4804 29106 4856 29112
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 4816 28558 4844 29106
rect 4804 28552 4856 28558
rect 4342 28520 4398 28529
rect 4804 28494 4856 28500
rect 4342 28455 4398 28464
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 4080 27606 4108 28018
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4264 27470 4292 28358
rect 4252 27464 4304 27470
rect 4252 27406 4304 27412
rect 4356 27316 4384 28358
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 4908 27402 4936 30194
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 5000 29102 5028 29582
rect 5184 29510 5212 30534
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 5264 29776 5316 29782
rect 5264 29718 5316 29724
rect 5172 29504 5224 29510
rect 5172 29446 5224 29452
rect 5184 29306 5212 29446
rect 5172 29300 5224 29306
rect 5172 29242 5224 29248
rect 4988 29096 5040 29102
rect 4988 29038 5040 29044
rect 4988 28484 5040 28490
rect 4988 28426 5040 28432
rect 5080 28484 5132 28490
rect 5080 28426 5132 28432
rect 5000 27470 5028 28426
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 4264 27288 4384 27316
rect 4066 26888 4122 26897
rect 4066 26823 4068 26832
rect 4120 26823 4122 26832
rect 4160 26852 4212 26858
rect 4068 26794 4120 26800
rect 4160 26794 4212 26800
rect 4172 26450 4200 26794
rect 4160 26444 4212 26450
rect 4160 26386 4212 26392
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4080 24818 4108 26250
rect 4068 24812 4120 24818
rect 3896 24772 4016 24800
rect 3988 24596 4016 24772
rect 4068 24754 4120 24760
rect 4068 24608 4120 24614
rect 3988 24568 4068 24596
rect 4068 24550 4120 24556
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3974 24168 4030 24177
rect 3896 23866 3924 24142
rect 3974 24103 4030 24112
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3988 23798 4016 24103
rect 3976 23792 4028 23798
rect 3976 23734 4028 23740
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 3896 22522 3924 23666
rect 4068 23588 4120 23594
rect 4068 23530 4120 23536
rect 4080 23322 4108 23530
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4080 22574 4108 22918
rect 3976 22568 4028 22574
rect 3896 22516 3976 22522
rect 3896 22510 4028 22516
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 3896 22494 4016 22510
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3528 20602 3556 20878
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3422 19952 3478 19961
rect 3422 19887 3478 19896
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3160 19394 3188 19450
rect 3160 19366 3280 19394
rect 3068 18822 3188 18850
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2962 18592 3018 18601
rect 2962 18527 3018 18536
rect 2976 18408 3004 18527
rect 2884 18380 3004 18408
rect 2884 18290 2912 18380
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2792 16726 2820 17070
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 16232 2636 16458
rect 2516 16204 2636 16232
rect 2516 16114 2544 16204
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2608 14822 2636 16050
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 2780 15564 2832 15570
rect 2700 15502 2728 15535
rect 2780 15506 2832 15512
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2792 15434 2820 15506
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2318 12271 2374 12280
rect 2412 12300 2464 12306
rect 1766 12064 1822 12073
rect 1766 11999 1822 12008
rect 1780 11830 1808 11999
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1872 11218 1900 12260
rect 2412 12242 2464 12248
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1858 11112 1914 11121
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1400 9648 1452 9654
rect 1398 9616 1400 9625
rect 1452 9616 1454 9625
rect 1398 9551 1454 9560
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1216 5840 1268 5846
rect 1216 5782 1268 5788
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 480 3936 532 3942
rect 480 3878 532 3884
rect 492 3777 520 3878
rect 478 3768 534 3777
rect 478 3703 534 3712
rect 1596 3058 1624 9862
rect 1688 9586 1716 10474
rect 1780 9625 1808 11086
rect 1858 11047 1860 11056
rect 1912 11047 1914 11056
rect 1860 11018 1912 11024
rect 1964 10810 1992 12106
rect 2148 11830 2176 12174
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9761 1900 9998
rect 2056 9926 2084 11630
rect 2148 10470 2176 11766
rect 2240 10742 2268 12106
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1858 9752 1914 9761
rect 1858 9687 1914 9696
rect 1766 9616 1822 9625
rect 1676 9580 1728 9586
rect 1766 9551 1822 9560
rect 1676 9522 1728 9528
rect 1688 8498 1716 9522
rect 1766 9208 1822 9217
rect 1766 9143 1768 9152
rect 1820 9143 1822 9152
rect 1768 9114 1820 9120
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7954 1716 8434
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 7478 1716 7890
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1688 6798 1716 7414
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6322 1716 6734
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1688 5234 1716 6258
rect 1858 5808 1914 5817
rect 1858 5743 1860 5752
rect 1912 5743 1914 5752
rect 1860 5714 1912 5720
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 4690 1716 5170
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4146 1716 4626
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3602 1716 4082
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1688 2774 1716 3538
rect 1872 3058 1900 5714
rect 2148 3126 2176 10134
rect 2240 9586 2268 10678
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2332 8566 2360 11018
rect 2424 10606 2452 11698
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2318 8256 2374 8265
rect 2318 8191 2374 8200
rect 2332 7886 2360 8191
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2424 5794 2452 9930
rect 2516 9178 2544 13874
rect 2608 10742 2636 14758
rect 2700 14346 2728 14826
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2688 12912 2740 12918
rect 2792 12866 2820 13806
rect 2740 12860 2820 12866
rect 2688 12854 2820 12860
rect 2700 12838 2820 12854
rect 2792 11914 2820 12838
rect 2884 12481 2912 14962
rect 2976 14278 3004 18226
rect 3068 15910 3096 18702
rect 3160 18086 3188 18822
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3252 17898 3280 19366
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3344 18057 3372 18702
rect 3330 18048 3386 18057
rect 3330 17983 3386 17992
rect 3252 17870 3372 17898
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3252 17270 3280 17614
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 3068 13802 3096 15302
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3068 12850 3096 13738
rect 3160 13530 3188 16526
rect 3252 15638 3280 17206
rect 3344 16998 3372 17870
rect 3436 17746 3464 19887
rect 3528 19417 3556 20402
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3620 19258 3648 19790
rect 3528 19230 3648 19258
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2870 12472 2926 12481
rect 2870 12407 2926 12416
rect 2792 11886 2912 11914
rect 2976 11898 3004 12718
rect 3068 12594 3096 12786
rect 3160 12714 3188 13466
rect 3252 12782 3280 15370
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 13802 3372 14894
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3436 12986 3464 17546
rect 3528 15570 3556 19230
rect 3712 19174 3740 20810
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19446 3832 20198
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3620 18222 3648 19110
rect 3792 18760 3844 18766
rect 3790 18728 3792 18737
rect 3844 18728 3846 18737
rect 3790 18663 3846 18672
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3620 16572 3648 18158
rect 3712 16697 3740 18294
rect 3790 17640 3846 17649
rect 3790 17575 3846 17584
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 3804 16590 3832 17575
rect 3792 16584 3844 16590
rect 3620 16544 3740 16572
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3528 15314 3556 15506
rect 3528 15286 3648 15314
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3424 12980 3476 12986
rect 3344 12940 3424 12968
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3068 12566 3188 12594
rect 3160 12306 3188 12566
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2594 10432 2650 10441
rect 2594 10367 2650 10376
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2608 8974 2636 10367
rect 2700 9110 2728 11086
rect 2792 10198 2820 11698
rect 2884 11558 2912 11886
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8650 2728 8842
rect 2792 8650 2820 9590
rect 2884 8906 2912 11018
rect 2976 11014 3004 11630
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10130 3004 10950
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 9722 3004 10066
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2700 8622 2820 8650
rect 2424 5766 2544 5794
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2424 3942 2452 5578
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2516 3738 2544 5766
rect 2792 4010 2820 8622
rect 3068 8090 3096 11834
rect 3160 10441 3188 12242
rect 3252 12102 3280 12718
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11286 3280 12038
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3146 10432 3202 10441
rect 3146 10367 3202 10376
rect 3252 9654 3280 10678
rect 3240 9648 3292 9654
rect 3146 9616 3202 9625
rect 3240 9590 3292 9596
rect 3146 9551 3202 9560
rect 3160 8956 3188 9551
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 9081 3280 9114
rect 3238 9072 3294 9081
rect 3238 9007 3294 9016
rect 3160 8928 3280 8956
rect 3252 8838 3280 8928
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2962 6760 3018 6769
rect 2962 6695 3018 6704
rect 2976 6662 3004 6695
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2976 5914 3004 6190
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 2976 2922 3004 3402
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1596 2746 1716 2774
rect 1596 2446 1624 2746
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1688 2446 1716 2479
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1596 1426 1624 2382
rect 2596 2032 2648 2038
rect 2594 2000 2596 2009
rect 2648 2000 2650 2009
rect 2594 1935 2650 1944
rect 1584 1420 1636 1426
rect 1584 1362 1636 1368
rect 2792 1358 2820 2790
rect 3068 2774 3096 7919
rect 3252 6866 3280 8774
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3344 5914 3372 12940
rect 3424 12922 3476 12928
rect 3528 11898 3556 15098
rect 3620 13258 3648 15286
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3620 12850 3648 13194
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3436 11150 3464 11222
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10810 3464 11086
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 9178 3464 10542
rect 3528 10062 3556 11698
rect 3712 11558 3740 16544
rect 3792 16526 3844 16532
rect 3896 16250 3924 22494
rect 4172 21554 4200 23462
rect 4264 23236 4292 27288
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4816 26081 4844 26930
rect 4802 26072 4858 26081
rect 4802 26007 4858 26016
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4816 24721 4844 25842
rect 4908 25265 4936 27338
rect 5000 26994 5028 27406
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 5000 26518 5028 26930
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 5092 26382 5120 28426
rect 5184 28218 5212 29242
rect 5276 29170 5304 29718
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5172 28212 5224 28218
rect 5172 28154 5224 28160
rect 5184 28082 5212 28154
rect 5172 28076 5224 28082
rect 5172 28018 5224 28024
rect 5184 27606 5212 28018
rect 5264 28008 5316 28014
rect 5262 27976 5264 27985
rect 5316 27976 5318 27985
rect 5262 27911 5318 27920
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 5276 27470 5304 27911
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5368 26382 5396 29582
rect 5552 29034 5580 30330
rect 5736 29714 5764 30670
rect 6000 30184 6052 30190
rect 6000 30126 6052 30132
rect 5816 30116 5868 30122
rect 5816 30058 5868 30064
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5828 29594 5856 30058
rect 5736 29578 5856 29594
rect 5724 29572 5856 29578
rect 5776 29566 5856 29572
rect 5724 29514 5776 29520
rect 5540 29028 5592 29034
rect 5540 28970 5592 28976
rect 5448 28960 5500 28966
rect 5448 28902 5500 28908
rect 5080 26376 5132 26382
rect 5264 26376 5316 26382
rect 5080 26318 5132 26324
rect 5262 26344 5264 26353
rect 5356 26376 5408 26382
rect 5316 26344 5318 26353
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 4894 25256 4950 25265
rect 4894 25191 4950 25200
rect 4802 24712 4858 24721
rect 4802 24647 4858 24656
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4816 24392 4844 24647
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4632 24364 4844 24392
rect 4344 24132 4396 24138
rect 4344 24074 4396 24080
rect 4356 23633 4384 24074
rect 4632 23866 4660 24364
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4436 23860 4488 23866
rect 4436 23802 4488 23808
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4342 23624 4398 23633
rect 4342 23559 4398 23568
rect 4448 23508 4476 23802
rect 4724 23662 4752 24142
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4356 23480 4476 23508
rect 4356 23304 4384 23480
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4356 23276 4568 23304
rect 4264 23208 4476 23236
rect 4448 23118 4476 23208
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4264 21554 4292 22918
rect 4344 22500 4396 22506
rect 4540 22488 4568 23276
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4632 22545 4660 23054
rect 4396 22460 4568 22488
rect 4618 22536 4674 22545
rect 4618 22471 4674 22480
rect 4344 22442 4396 22448
rect 4356 21962 4384 22442
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4344 21956 4396 21962
rect 4344 21898 4396 21904
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3988 20058 4016 21422
rect 4724 21332 4752 22170
rect 4816 22030 4844 24006
rect 4908 23526 4936 24550
rect 5000 24206 5028 26250
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4894 23352 4950 23361
rect 4894 23287 4950 23296
rect 4908 22817 4936 23287
rect 5000 23118 5028 24142
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4894 22808 4950 22817
rect 5000 22778 5028 23054
rect 4894 22743 4950 22752
rect 4988 22772 5040 22778
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4908 21962 4936 22743
rect 4988 22714 5040 22720
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4896 21616 4948 21622
rect 4896 21558 4948 21564
rect 4724 21304 4844 21332
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3974 19952 4030 19961
rect 3974 19887 4030 19896
rect 3988 19854 4016 19887
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 3988 17814 4016 19382
rect 4080 18086 4108 20742
rect 4172 20398 4200 21014
rect 4436 20936 4488 20942
rect 4434 20904 4436 20913
rect 4488 20904 4490 20913
rect 4434 20839 4490 20848
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4158 20224 4214 20233
rect 4158 20159 4214 20168
rect 4172 19854 4200 20159
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4172 18970 4200 19314
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4264 18902 4292 20470
rect 4356 18902 4384 20742
rect 4712 20528 4764 20534
rect 4434 20496 4490 20505
rect 4816 20516 4844 21304
rect 4764 20488 4844 20516
rect 4712 20470 4764 20476
rect 4434 20431 4436 20440
rect 4488 20431 4490 20440
rect 4436 20402 4488 20408
rect 4724 20262 4752 20470
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4712 19848 4764 19854
rect 4434 19816 4490 19825
rect 4712 19790 4764 19796
rect 4434 19751 4490 19760
rect 4448 19514 4476 19751
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4724 19281 4752 19790
rect 4816 19786 4844 20266
rect 4908 20058 4936 21558
rect 5000 20602 5028 22510
rect 5092 22234 5120 26318
rect 5356 26318 5408 26324
rect 5262 26279 5318 26288
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5368 24993 5396 25094
rect 5354 24984 5410 24993
rect 5264 24948 5316 24954
rect 5184 24908 5264 24936
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5092 20942 5120 21966
rect 5184 21554 5212 24908
rect 5354 24919 5410 24928
rect 5264 24890 5316 24896
rect 5460 24886 5488 28902
rect 5736 28082 5764 29514
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 6012 28014 6040 30126
rect 6104 29782 6132 30806
rect 6092 29776 6144 29782
rect 6092 29718 6144 29724
rect 6000 28008 6052 28014
rect 6000 27950 6052 27956
rect 5908 27940 5960 27946
rect 5908 27882 5960 27888
rect 5920 27849 5948 27882
rect 5906 27840 5962 27849
rect 5906 27775 5962 27784
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5552 25430 5580 27406
rect 5644 25906 5672 27406
rect 5736 27334 5764 27542
rect 6012 27470 6040 27950
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 6092 27056 6144 27062
rect 6092 26998 6144 27004
rect 5908 26852 5960 26858
rect 5908 26794 5960 26800
rect 5816 26512 5868 26518
rect 5816 26454 5868 26460
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5540 25424 5592 25430
rect 5540 25366 5592 25372
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5276 21690 5304 24142
rect 5368 22409 5396 24754
rect 5460 24410 5488 24822
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5540 24200 5592 24206
rect 5538 24168 5540 24177
rect 5592 24168 5594 24177
rect 5538 24103 5594 24112
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5552 22778 5580 23054
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5354 22400 5410 22409
rect 5354 22335 5410 22344
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5368 22098 5396 22170
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 21049 5212 21490
rect 5368 21457 5396 21830
rect 5460 21554 5488 22442
rect 5540 21888 5592 21894
rect 5538 21856 5540 21865
rect 5592 21856 5594 21865
rect 5538 21791 5594 21800
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5354 21448 5410 21457
rect 5354 21383 5410 21392
rect 5460 21332 5488 21490
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5276 21304 5488 21332
rect 5276 21078 5304 21304
rect 5446 21176 5502 21185
rect 5446 21111 5448 21120
rect 5500 21111 5502 21120
rect 5448 21082 5500 21088
rect 5552 21078 5580 21422
rect 5264 21072 5316 21078
rect 5170 21040 5226 21049
rect 5540 21072 5592 21078
rect 5264 21014 5316 21020
rect 5354 21040 5410 21049
rect 5170 20975 5226 20984
rect 5540 21014 5592 21020
rect 5354 20975 5410 20984
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5092 20602 5120 20878
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 5078 20496 5134 20505
rect 4988 20460 5040 20466
rect 5078 20431 5134 20440
rect 4988 20402 5040 20408
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4710 19272 4766 19281
rect 4710 19207 4766 19216
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4436 18896 4488 18902
rect 4816 18850 4844 19450
rect 4436 18838 4488 18844
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4172 17882 4200 18770
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 4068 17604 4120 17610
rect 3988 17564 4068 17592
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3804 15473 3832 16186
rect 3988 15586 4016 17564
rect 4068 17546 4120 17552
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4172 16697 4200 17138
rect 4158 16688 4214 16697
rect 4158 16623 4214 16632
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4172 16266 4200 16458
rect 4264 16454 4292 18702
rect 4344 18284 4396 18290
rect 4448 18272 4476 18838
rect 4724 18822 4844 18850
rect 4724 18766 4752 18822
rect 4908 18766 4936 19790
rect 5000 19553 5028 20402
rect 4986 19544 5042 19553
rect 4986 19479 5042 19488
rect 5000 19378 5028 19479
rect 5092 19446 5120 20431
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5184 19514 5212 19858
rect 5276 19553 5304 20878
rect 5262 19544 5318 19553
rect 5172 19508 5224 19514
rect 5262 19479 5318 19488
rect 5172 19450 5224 19456
rect 5080 19440 5132 19446
rect 5080 19382 5132 19388
rect 4988 19372 5040 19378
rect 5264 19372 5316 19378
rect 4988 19314 5040 19320
rect 5184 19332 5264 19360
rect 5000 18902 5028 19314
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4988 18896 5040 18902
rect 4988 18838 5040 18844
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4528 18420 4580 18426
rect 4580 18380 4844 18408
rect 4528 18362 4580 18368
rect 4396 18244 4476 18272
rect 4528 18284 4580 18290
rect 4344 18226 4396 18232
rect 4528 18226 4580 18232
rect 4816 18272 4844 18380
rect 4908 18290 4936 18702
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4896 18284 4948 18290
rect 4816 18244 4896 18272
rect 4540 18193 4568 18226
rect 4620 18216 4672 18222
rect 4526 18184 4582 18193
rect 4620 18158 4672 18164
rect 4526 18119 4582 18128
rect 4632 18068 4660 18158
rect 4356 18040 4660 18068
rect 4356 17882 4384 18040
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4342 17776 4398 17785
rect 4342 17711 4344 17720
rect 4396 17711 4398 17720
rect 4344 17682 4396 17688
rect 4816 17320 4844 18244
rect 4896 18226 4948 18232
rect 5000 17921 5028 18362
rect 4986 17912 5042 17921
rect 4986 17847 5042 17856
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4724 17292 4844 17320
rect 4724 17202 4752 17292
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4436 17128 4488 17134
rect 4356 17088 4436 17116
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4356 16266 4384 17088
rect 4436 17070 4488 17076
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4712 16516 4764 16522
rect 4816 16504 4844 17138
rect 4764 16476 4844 16504
rect 4712 16458 4764 16464
rect 4172 16238 4292 16266
rect 4356 16238 4568 16266
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15706 4108 16050
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3896 15558 4016 15586
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3896 15366 3924 15558
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9518 3556 9998
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3528 5545 3556 9318
rect 3620 8906 3648 11494
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3712 9654 3740 9930
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3514 5536 3570 5545
rect 3514 5471 3570 5480
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 2976 2746 3096 2774
rect 2976 2650 3004 2746
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3528 2106 3556 4150
rect 3620 3194 3648 8842
rect 3712 8498 3740 9590
rect 3804 8566 3832 14894
rect 3988 14482 4016 15302
rect 4080 14550 4108 15642
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 14618 4200 15438
rect 4264 14822 4292 16238
rect 4540 15892 4568 16238
rect 4724 16114 4752 16458
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4540 15864 4844 15892
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4816 15638 4844 15864
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 4080 14006 4108 14486
rect 4160 14408 4212 14414
rect 4264 14396 4292 14758
rect 4212 14368 4292 14396
rect 4160 14350 4212 14356
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3896 12306 3924 13874
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3896 11898 3924 12242
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3988 11354 4016 13806
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12646 4108 13262
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4172 11830 4200 13126
rect 4264 12782 4292 13806
rect 4356 12986 4384 14962
rect 4448 14958 4476 15438
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4816 14600 4844 15370
rect 4908 15348 4936 17614
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 15502 5028 17478
rect 5092 17202 5120 19110
rect 5184 18737 5212 19332
rect 5264 19314 5316 19320
rect 5170 18728 5226 18737
rect 5170 18663 5226 18672
rect 5184 17678 5212 18663
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5276 17202 5304 18566
rect 5368 18426 5396 20975
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5460 20505 5488 20878
rect 5446 20496 5502 20505
rect 5446 20431 5502 20440
rect 5448 20392 5500 20398
rect 5446 20360 5448 20369
rect 5500 20360 5502 20369
rect 5446 20295 5502 20304
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5460 19378 5488 19926
rect 5552 19553 5580 20198
rect 5644 19922 5672 24346
rect 5736 23798 5764 26182
rect 5828 25242 5856 26454
rect 5920 26042 5948 26794
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 5908 25764 5960 25770
rect 5908 25706 5960 25712
rect 5920 25362 5948 25706
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5828 25214 5948 25242
rect 5814 24848 5870 24857
rect 5814 24783 5816 24792
rect 5868 24783 5870 24792
rect 5816 24754 5868 24760
rect 5920 24274 5948 25214
rect 6012 24886 6040 26522
rect 6104 24954 6132 26998
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 5908 24268 5960 24274
rect 5828 24228 5908 24256
rect 5724 23792 5776 23798
rect 5724 23734 5776 23740
rect 5736 23361 5764 23734
rect 5828 23497 5856 24228
rect 5908 24210 5960 24216
rect 6012 24138 6040 24550
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 6104 24018 6132 24074
rect 5920 23990 6132 24018
rect 5814 23488 5870 23497
rect 5814 23423 5870 23432
rect 5722 23352 5778 23361
rect 5828 23322 5856 23423
rect 5722 23287 5778 23296
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5722 23216 5778 23225
rect 5722 23151 5778 23160
rect 5736 23118 5764 23151
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5736 22137 5764 23054
rect 5816 23044 5868 23050
rect 5816 22986 5868 22992
rect 5722 22128 5778 22137
rect 5722 22063 5778 22072
rect 5828 22030 5856 22986
rect 5920 22098 5948 23990
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6196 23066 6224 26862
rect 6288 23866 6316 27406
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 6380 26382 6408 27270
rect 6472 26450 6500 31214
rect 6564 30734 6592 31758
rect 6656 31278 6684 32302
rect 6644 31272 6696 31278
rect 6644 31214 6696 31220
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 6736 30660 6788 30666
rect 6736 30602 6788 30608
rect 6748 29170 6776 30602
rect 6840 30258 6868 30670
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 6736 29164 6788 29170
rect 6656 29124 6736 29152
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 6368 25356 6420 25362
rect 6368 25298 6420 25304
rect 6380 24886 6408 25298
rect 6472 25294 6500 25842
rect 6564 25401 6592 29038
rect 6656 27334 6684 29124
rect 6736 29106 6788 29112
rect 6736 29028 6788 29034
rect 6736 28970 6788 28976
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6656 26489 6684 26930
rect 6642 26480 6698 26489
rect 6642 26415 6698 26424
rect 6644 26308 6696 26314
rect 6644 26250 6696 26256
rect 6550 25392 6606 25401
rect 6550 25327 6606 25336
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6550 25256 6606 25265
rect 6472 24954 6500 25230
rect 6550 25191 6606 25200
rect 6564 25158 6592 25191
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6368 24880 6420 24886
rect 6368 24822 6420 24828
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6368 24676 6420 24682
rect 6368 24618 6420 24624
rect 6380 23866 6408 24618
rect 6564 24138 6592 24822
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6460 24064 6512 24070
rect 6458 24032 6460 24041
rect 6512 24032 6514 24041
rect 6458 23967 6514 23976
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6012 22574 6040 23054
rect 6196 23038 6316 23066
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5816 22024 5868 22030
rect 5736 21984 5816 22012
rect 5736 20466 5764 21984
rect 5816 21966 5868 21972
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5632 19712 5684 19718
rect 5630 19680 5632 19689
rect 5684 19680 5686 19689
rect 5630 19615 5686 19624
rect 5538 19544 5594 19553
rect 5538 19479 5594 19488
rect 5552 19378 5580 19479
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18601 5580 19110
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5538 18592 5594 18601
rect 5538 18527 5594 18536
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5644 17882 5672 18634
rect 5736 18630 5764 20402
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17202 5396 17478
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5276 17082 5304 17138
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5172 17060 5224 17066
rect 5276 17054 5396 17082
rect 5172 17002 5224 17008
rect 4988 15496 5040 15502
rect 5092 15484 5120 17002
rect 5184 16454 5212 17002
rect 5368 16794 5396 17054
rect 5552 16794 5580 17818
rect 5644 17678 5672 17818
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5736 17524 5764 17750
rect 5644 17496 5764 17524
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5276 16114 5304 16662
rect 5644 16436 5672 17496
rect 5828 17338 5856 21490
rect 5920 20534 5948 22034
rect 6104 21350 6132 22918
rect 6196 22710 6224 22918
rect 6184 22704 6236 22710
rect 6184 22646 6236 22652
rect 6288 22001 6316 23038
rect 6380 22556 6408 23598
rect 6472 22710 6500 23666
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6460 22704 6512 22710
rect 6460 22646 6512 22652
rect 6380 22528 6500 22556
rect 6366 22400 6422 22409
rect 6366 22335 6422 22344
rect 6274 21992 6330 22001
rect 6274 21927 6330 21936
rect 6288 21690 6316 21927
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 5908 20528 5960 20534
rect 6380 20482 6408 22335
rect 6472 21962 6500 22528
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6564 21894 6592 23190
rect 6656 23186 6684 26250
rect 6748 25294 6776 28970
rect 6828 28552 6880 28558
rect 6826 28520 6828 28529
rect 6880 28520 6882 28529
rect 6826 28455 6882 28464
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6840 26926 6868 28018
rect 6932 27538 6960 33254
rect 7012 32428 7064 32434
rect 7012 32370 7064 32376
rect 7024 31754 7052 32370
rect 7472 32360 7524 32366
rect 7472 32302 7524 32308
rect 7196 32292 7248 32298
rect 7196 32234 7248 32240
rect 7024 31726 7144 31754
rect 7012 30320 7064 30326
rect 7012 30262 7064 30268
rect 7116 30274 7144 31726
rect 7208 31414 7236 32234
rect 7196 31408 7248 31414
rect 7196 31350 7248 31356
rect 7484 31278 7512 32302
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 7484 30598 7512 31214
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7024 28966 7052 30262
rect 7116 30246 7236 30274
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 7024 28082 7052 28902
rect 7012 28076 7064 28082
rect 7012 28018 7064 28024
rect 7024 27946 7052 28018
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 6920 27532 6972 27538
rect 6920 27474 6972 27480
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 6918 27024 6974 27033
rect 7024 26994 7052 27338
rect 6918 26959 6974 26968
rect 7012 26988 7064 26994
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 25430 6868 26862
rect 6932 26840 6960 26959
rect 7012 26930 7064 26936
rect 7012 26852 7064 26858
rect 6932 26812 7012 26840
rect 7012 26794 7064 26800
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6932 25770 6960 26318
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6736 25288 6788 25294
rect 6840 25265 6868 25366
rect 6736 25230 6788 25236
rect 6826 25256 6882 25265
rect 6826 25191 6882 25200
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6748 22522 6776 23802
rect 6840 23118 6868 25094
rect 6932 24818 6960 25094
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6932 23905 6960 24754
rect 7024 24177 7052 26794
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 6918 23896 6974 23905
rect 6918 23831 6974 23840
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 23633 7052 23666
rect 7010 23624 7066 23633
rect 6920 23588 6972 23594
rect 7010 23559 7066 23568
rect 6920 23530 6972 23536
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6748 22494 6868 22522
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21078 6592 21830
rect 6656 21622 6684 21898
rect 6748 21622 6776 22374
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6642 21040 6698 21049
rect 6642 20975 6644 20984
rect 6696 20975 6698 20984
rect 6644 20946 6696 20952
rect 6748 20534 6776 21558
rect 5908 20470 5960 20476
rect 6012 20454 6408 20482
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 18154 5948 19790
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 6012 17338 6040 20454
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6104 19854 6132 20266
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6104 19174 6132 19382
rect 6196 19378 6224 19722
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6104 18698 6132 19110
rect 6196 18766 6224 19314
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 18692 6144 18698
rect 6092 18634 6144 18640
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6090 17912 6146 17921
rect 6090 17847 6146 17856
rect 6104 17542 6132 17847
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5816 17332 5868 17338
rect 6000 17332 6052 17338
rect 5816 17274 5868 17280
rect 5920 17292 6000 17320
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5828 17105 5856 17138
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16590 5856 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5724 16448 5776 16454
rect 5644 16408 5724 16436
rect 5724 16390 5776 16396
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5264 15496 5316 15502
rect 5092 15456 5264 15484
rect 4988 15438 5040 15444
rect 5264 15438 5316 15444
rect 4908 15320 5212 15348
rect 4540 14572 4844 14600
rect 4540 14414 4568 14572
rect 5184 14498 5212 15320
rect 5276 14618 5304 15438
rect 5368 14890 5396 16118
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5552 15502 5580 15846
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5644 15162 5672 15846
rect 5736 15570 5764 16390
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5736 14958 5764 15506
rect 5828 15366 5856 16526
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5080 14476 5132 14482
rect 5184 14470 5304 14498
rect 5080 14418 5132 14424
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4540 14249 4568 14350
rect 4526 14240 4582 14249
rect 4526 14175 4582 14184
rect 4712 13932 4764 13938
rect 4816 13920 4844 14350
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4908 13938 4936 14282
rect 5092 13938 5120 14418
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 4764 13892 4844 13920
rect 4712 13874 4764 13880
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 13190 4660 13262
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4342 12880 4398 12889
rect 4342 12815 4398 12824
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4264 12442 4292 12718
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4356 12102 4384 12815
rect 4724 12782 4752 13398
rect 4816 12850 4844 13892
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4908 13462 4936 13738
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12918 4936 13262
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4712 12776 4764 12782
rect 4764 12724 4844 12730
rect 4712 12718 4844 12724
rect 4724 12702 4844 12718
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4816 12434 4844 12702
rect 4724 12406 4844 12434
rect 4724 12306 4752 12406
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3974 10296 4030 10305
rect 3974 10231 3976 10240
rect 4028 10231 4030 10240
rect 3976 10202 4028 10208
rect 3988 9874 4016 10202
rect 3896 9846 4016 9874
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 6390 3740 7142
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3712 5574 3740 6326
rect 3896 6118 3924 9846
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3988 9042 4016 9658
rect 4080 9586 4108 11630
rect 4172 11121 4200 11766
rect 4356 11234 4384 12038
rect 4724 11898 4752 12242
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4724 11762 4752 11834
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4252 11212 4304 11218
rect 4356 11206 4476 11234
rect 4252 11154 4304 11160
rect 4158 11112 4214 11121
rect 4158 11047 4214 11056
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4172 9382 4200 10950
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4080 8294 4108 9318
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8498 4200 8774
rect 4264 8514 4292 11154
rect 4344 11144 4396 11150
rect 4342 11112 4344 11121
rect 4396 11112 4398 11121
rect 4342 11047 4398 11056
rect 4448 11014 4476 11206
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4356 10062 4384 10406
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4356 9382 4384 9522
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 8634 4384 9318
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4816 9178 4844 12174
rect 4908 11354 4936 12854
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4908 9466 4936 11086
rect 5000 9654 5028 13670
rect 5092 12850 5120 13874
rect 5184 13394 5212 14214
rect 5276 13734 5304 14470
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5092 12442 5120 12786
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5078 12336 5134 12345
rect 5078 12271 5134 12280
rect 5092 12238 5120 12271
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4988 9512 5040 9518
rect 4908 9460 4988 9466
rect 4908 9454 5040 9460
rect 4908 9438 5028 9454
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8634 4568 8910
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4160 8492 4212 8498
rect 4264 8486 4384 8514
rect 4632 8498 4660 8774
rect 4724 8498 4752 9114
rect 4908 9042 4936 9318
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4160 8434 4212 8440
rect 4356 8430 4384 8486
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4356 8090 4384 8366
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4908 8090 4936 8434
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4908 7970 4936 8026
rect 4816 7942 4936 7970
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5794 3924 6054
rect 3804 5766 3924 5794
rect 3804 5642 3832 5766
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 4690 3740 5510
rect 3804 5370 3832 5578
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3896 4554 3924 5646
rect 3988 5370 4016 7346
rect 4710 7304 4766 7313
rect 4710 7239 4712 7248
rect 4764 7239 4766 7248
rect 4712 7210 4764 7216
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4816 6730 4844 7942
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4908 7002 4936 7822
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4618 6488 4674 6497
rect 4618 6423 4620 6432
rect 4672 6423 4674 6432
rect 4620 6394 4672 6400
rect 4724 6390 4752 6598
rect 4816 6458 4844 6666
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5000 6390 5028 9438
rect 5092 9382 5120 12174
rect 5184 11762 5212 13223
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5276 11286 5304 13466
rect 5368 12986 5396 14826
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5736 14414 5764 14758
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 13870 5764 14350
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13728 5500 13734
rect 5828 13682 5856 15302
rect 5920 13841 5948 17292
rect 6000 17274 6052 17280
rect 6104 17218 6132 17478
rect 6012 17190 6132 17218
rect 6012 16114 6040 17190
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 15502 6040 15914
rect 6104 15706 6132 16526
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5906 13832 5962 13841
rect 5906 13767 5962 13776
rect 5448 13670 5500 13676
rect 5460 13394 5488 13670
rect 5736 13654 5856 13682
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 11280 5316 11286
rect 5184 11240 5264 11268
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4158 6216 4214 6225
rect 4158 6151 4214 6160
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 2780 1352 2832 1358
rect 2780 1294 2832 1300
rect 3988 678 4016 3878
rect 4080 3602 4108 5782
rect 4172 5234 4200 6151
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 4146 4200 5170
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4264 4010 4292 6258
rect 4356 6186 4384 6326
rect 5092 6322 5120 9046
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5710 4384 6122
rect 4802 6080 4858 6089
rect 4423 6012 4731 6021
rect 4802 6015 4858 6024
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4816 5370 4844 6015
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4356 4826 4384 5170
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4908 4622 4936 6258
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5000 5817 5028 6054
rect 4986 5808 5042 5817
rect 4986 5743 5042 5752
rect 5000 5098 5028 5743
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4986 4856 5042 4865
rect 4986 4791 4988 4800
rect 5040 4791 5042 4800
rect 4988 4762 5040 4768
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4078 4384 4422
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4816 3738 4844 4082
rect 5092 4049 5120 5510
rect 5078 4040 5134 4049
rect 5184 4010 5212 11240
rect 5264 11222 5316 11228
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 10810 5304 11086
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9586 5304 9862
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 7886 5304 9522
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7478 5304 7686
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5276 6798 5304 7414
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5368 6458 5396 12718
rect 5460 11082 5488 13126
rect 5644 12424 5672 13262
rect 5736 12986 5764 13654
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5552 12396 5672 12424
rect 5552 12084 5580 12396
rect 5552 12056 5672 12084
rect 5644 11762 5672 12056
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5552 11234 5580 11698
rect 5736 11354 5764 12786
rect 5828 12714 5856 13466
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5920 12594 5948 12650
rect 5828 12566 5948 12594
rect 5724 11348 5776 11354
rect 5828 11336 5856 12566
rect 5906 12472 5962 12481
rect 5906 12407 5908 12416
rect 5960 12407 5962 12416
rect 6092 12436 6144 12442
rect 5908 12378 5960 12384
rect 6092 12378 6144 12384
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11529 5948 12038
rect 5906 11520 5962 11529
rect 5906 11455 5962 11464
rect 5828 11308 5948 11336
rect 5724 11290 5776 11296
rect 5552 11206 5764 11234
rect 5448 11076 5500 11082
rect 5632 11076 5684 11082
rect 5448 11018 5500 11024
rect 5552 11036 5632 11064
rect 5552 10962 5580 11036
rect 5632 11018 5684 11024
rect 5460 10934 5580 10962
rect 5460 10606 5488 10934
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5552 10062 5580 10746
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10130 5672 10610
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 8974 5580 9998
rect 5632 9988 5684 9994
rect 5736 9976 5764 11206
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5684 9948 5764 9976
rect 5632 9930 5684 9936
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5644 8566 5672 9930
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9110 5764 9522
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5448 8560 5500 8566
rect 5540 8560 5592 8566
rect 5448 8502 5500 8508
rect 5538 8528 5540 8537
rect 5632 8560 5684 8566
rect 5592 8528 5594 8537
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5276 5642 5304 6394
rect 5460 6338 5488 8502
rect 5632 8502 5684 8508
rect 5538 8463 5594 8472
rect 5632 8424 5684 8430
rect 5538 8392 5594 8401
rect 5632 8366 5684 8372
rect 5538 8327 5594 8336
rect 5552 7546 5580 8327
rect 5644 7954 5672 8366
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5736 7886 5764 9046
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 6662 5672 7346
rect 5736 6866 5764 7822
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5368 6310 5488 6338
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5368 5370 5396 6310
rect 5446 6216 5502 6225
rect 5446 6151 5502 6160
rect 5460 5846 5488 6151
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5078 3975 5134 3984
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5368 3942 5396 5034
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3126 4200 3334
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4080 882 4108 2994
rect 4172 2106 4200 3062
rect 5000 2854 5028 3402
rect 5092 2990 5120 3402
rect 5460 3398 5488 5238
rect 5552 4758 5580 6054
rect 5828 5710 5856 11154
rect 5920 11098 5948 11308
rect 5920 11070 6040 11098
rect 6104 11082 6132 12378
rect 6012 11014 6040 11070
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5920 10146 5948 10950
rect 6012 10742 6040 10950
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5920 10130 6040 10146
rect 5920 10124 6052 10130
rect 5920 10118 6000 10124
rect 6000 10066 6052 10072
rect 5908 10056 5960 10062
rect 5906 10024 5908 10033
rect 5960 10024 5962 10033
rect 5906 9959 5962 9968
rect 6012 9897 6040 10066
rect 5998 9888 6054 9897
rect 5998 9823 6054 9832
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5644 3913 5672 4082
rect 5630 3904 5686 3913
rect 5630 3839 5686 3848
rect 5736 3670 5764 5510
rect 5920 5302 5948 8570
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6012 7886 6040 8502
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5814 5128 5870 5137
rect 5814 5063 5816 5072
rect 5868 5063 5870 5072
rect 5816 5034 5868 5040
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 3528 5776 3534
rect 5722 3496 5724 3505
rect 5776 3496 5778 3505
rect 5722 3431 5778 3440
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5354 3088 5410 3097
rect 5354 3023 5356 3032
rect 5408 3023 5410 3032
rect 5356 2994 5408 3000
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 4172 1426 4200 2042
rect 4724 1766 4752 2518
rect 5264 2440 5316 2446
rect 4802 2408 4858 2417
rect 5264 2382 5316 2388
rect 4802 2343 4858 2352
rect 4816 2310 4844 2343
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 5276 1970 5304 2382
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 4712 1760 4764 1766
rect 4712 1702 4764 1708
rect 4423 1660 4731 1669
rect 4423 1658 4429 1660
rect 4485 1658 4509 1660
rect 4565 1658 4589 1660
rect 4645 1658 4669 1660
rect 4725 1658 4731 1660
rect 4485 1606 4487 1658
rect 4667 1606 4669 1658
rect 4423 1604 4429 1606
rect 4485 1604 4509 1606
rect 4565 1604 4589 1606
rect 4645 1604 4669 1606
rect 4725 1604 4731 1606
rect 4423 1595 4731 1604
rect 4160 1420 4212 1426
rect 4160 1362 4212 1368
rect 5828 1222 5856 3538
rect 6012 1970 6040 6598
rect 6104 5710 6132 10406
rect 6196 8362 6224 18566
rect 6288 16182 6316 20198
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6458 18184 6514 18193
rect 6368 18148 6420 18154
rect 6458 18119 6514 18128
rect 6368 18090 6420 18096
rect 6380 16590 6408 18090
rect 6472 17882 6500 18119
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6564 17610 6592 19246
rect 6748 18834 6776 19858
rect 6840 18902 6868 22494
rect 6932 22234 6960 23530
rect 6920 22228 6972 22234
rect 7024 22216 7052 23559
rect 7116 22438 7144 30126
rect 7208 29170 7236 30246
rect 7380 30116 7432 30122
rect 7380 30058 7432 30064
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7208 28994 7236 29106
rect 7208 28966 7328 28994
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7208 28218 7236 28698
rect 7196 28212 7248 28218
rect 7196 28154 7248 28160
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 7208 23746 7236 27814
rect 7300 26518 7328 28966
rect 7392 28218 7420 30058
rect 7484 29646 7512 30534
rect 7576 30394 7604 31758
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 7668 30326 7696 33322
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 8300 32836 8352 32842
rect 8300 32778 8352 32784
rect 7896 32668 8204 32677
rect 7896 32666 7902 32668
rect 7958 32666 7982 32668
rect 8038 32666 8062 32668
rect 8118 32666 8142 32668
rect 8198 32666 8204 32668
rect 7958 32614 7960 32666
rect 8140 32614 8142 32666
rect 7896 32612 7902 32614
rect 7958 32612 7982 32614
rect 8038 32612 8062 32614
rect 8118 32612 8142 32614
rect 8198 32612 8204 32614
rect 7896 32603 8204 32612
rect 7748 32292 7800 32298
rect 7748 32234 7800 32240
rect 7760 31958 7788 32234
rect 8312 31958 8340 32778
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 7748 31952 7800 31958
rect 7748 31894 7800 31900
rect 8300 31952 8352 31958
rect 8300 31894 8352 31900
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 8312 31521 8340 31758
rect 8404 31754 8432 32438
rect 8496 31958 8524 33050
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 8484 31952 8536 31958
rect 8482 31920 8484 31929
rect 8536 31920 8538 31929
rect 8482 31855 8538 31864
rect 8404 31726 8708 31754
rect 8298 31512 8354 31521
rect 7840 31476 7892 31482
rect 8298 31447 8354 31456
rect 7840 31418 7892 31424
rect 7852 31210 7880 31418
rect 7840 31204 7892 31210
rect 7840 31146 7892 31152
rect 8312 30734 8340 31447
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 7656 30320 7708 30326
rect 7576 30268 7656 30274
rect 7576 30262 7708 30268
rect 7576 30246 7696 30262
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7576 29170 7604 30246
rect 7656 30184 7708 30190
rect 7654 30152 7656 30161
rect 7708 30152 7710 30161
rect 7654 30087 7710 30096
rect 8576 29776 8628 29782
rect 8576 29718 8628 29724
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 8312 29170 8340 29650
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29306 8524 29446
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8298 29064 8354 29073
rect 8588 29034 8616 29718
rect 8298 28999 8354 29008
rect 8576 29028 8628 29034
rect 7748 28688 7800 28694
rect 7748 28630 7800 28636
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7380 28212 7432 28218
rect 7380 28154 7432 28160
rect 7380 28076 7432 28082
rect 7380 28018 7432 28024
rect 7288 26512 7340 26518
rect 7288 26454 7340 26460
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7300 25401 7328 25638
rect 7286 25392 7342 25401
rect 7286 25327 7342 25336
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7300 25129 7328 25162
rect 7286 25120 7342 25129
rect 7286 25055 7342 25064
rect 7392 24954 7420 28018
rect 7484 28014 7512 28494
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7484 27334 7512 27542
rect 7472 27328 7524 27334
rect 7472 27270 7524 27276
rect 7484 26042 7512 27270
rect 7760 26994 7788 28630
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7668 25702 7696 26862
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7562 25528 7618 25537
rect 7472 25492 7524 25498
rect 7562 25463 7618 25472
rect 7472 25434 7524 25440
rect 7380 24948 7432 24954
rect 7380 24890 7432 24896
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7380 24744 7432 24750
rect 7380 24686 7432 24692
rect 7300 23866 7328 24686
rect 7392 24206 7420 24686
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7208 23718 7328 23746
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7208 22506 7236 22986
rect 7196 22500 7248 22506
rect 7196 22442 7248 22448
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7024 22188 7144 22216
rect 6920 22170 6972 22176
rect 6932 22098 6960 22170
rect 7010 22128 7066 22137
rect 6920 22092 6972 22098
rect 7010 22063 7066 22072
rect 6920 22034 6972 22040
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6932 21350 6960 21490
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 17660 6684 18702
rect 6826 18048 6882 18057
rect 6826 17983 6882 17992
rect 6736 17672 6788 17678
rect 6656 17632 6736 17660
rect 6736 17614 6788 17620
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17338 6592 17546
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6380 14618 6408 16526
rect 6472 16454 6500 17138
rect 6748 16998 6776 17614
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6748 16658 6776 16934
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6460 16176 6512 16182
rect 6458 16144 6460 16153
rect 6512 16144 6514 16153
rect 6458 16079 6514 16088
rect 6472 15366 6500 16079
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6380 14414 6408 14554
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6288 12918 6316 13194
rect 6380 13190 6408 14350
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6472 14074 6500 14282
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6472 13977 6500 14010
rect 6458 13968 6514 13977
rect 6458 13903 6514 13912
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 13258 6500 13670
rect 6564 13462 6592 16594
rect 6656 15337 6684 16594
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6748 15026 6776 15098
rect 6736 15020 6788 15026
rect 6656 14980 6736 15008
rect 6656 13802 6684 14980
rect 6736 14962 6788 14968
rect 6734 13968 6790 13977
rect 6734 13903 6790 13912
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6288 11218 6316 12854
rect 6472 12714 6500 13194
rect 6564 13002 6592 13398
rect 6564 12974 6684 13002
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6380 11098 6408 12582
rect 6458 12472 6514 12481
rect 6564 12442 6592 12786
rect 6458 12407 6514 12416
rect 6552 12436 6604 12442
rect 6472 12306 6500 12407
rect 6656 12434 6684 12974
rect 6748 12646 6776 13903
rect 6840 12850 6868 17983
rect 6932 17898 6960 21286
rect 7024 21146 7052 22063
rect 7116 22030 7144 22188
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7102 21584 7158 21593
rect 7102 21519 7104 21528
rect 7156 21519 7158 21528
rect 7104 21490 7156 21496
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7010 20632 7066 20641
rect 7010 20567 7066 20576
rect 7024 19334 7052 20567
rect 7102 20224 7158 20233
rect 7102 20159 7158 20168
rect 7116 19854 7144 20159
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7024 19306 7144 19334
rect 7116 18222 7144 19306
rect 7194 19272 7250 19281
rect 7194 19207 7250 19216
rect 7208 18698 7236 19207
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7208 18426 7236 18634
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6932 17870 7144 17898
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 7024 16794 7052 17750
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16250 7052 16390
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7010 16144 7066 16153
rect 7116 16114 7144 17870
rect 7208 17610 7236 18362
rect 7300 18290 7328 23718
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7392 23322 7420 23666
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 22166 7420 22510
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 7378 21856 7434 21865
rect 7378 21791 7434 21800
rect 7392 20466 7420 21791
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 19446 7420 20198
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 17066 7236 17546
rect 7300 17202 7328 18226
rect 7392 17338 7420 19382
rect 7484 19378 7512 25434
rect 7576 21146 7604 25463
rect 7654 25256 7710 25265
rect 7654 25191 7710 25200
rect 7668 24410 7696 25191
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7668 22234 7696 24210
rect 7760 22778 7788 26318
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 8312 26024 8340 28999
rect 8576 28970 8628 28976
rect 8484 28144 8536 28150
rect 8484 28086 8536 28092
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8404 26586 8432 27270
rect 8496 26994 8524 28086
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8496 26432 8524 26930
rect 8680 26518 8708 31726
rect 9048 31482 9076 32302
rect 9036 31476 9088 31482
rect 9036 31418 9088 31424
rect 9048 31346 9076 31418
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 9048 30802 9076 31282
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 9036 30796 9088 30802
rect 9036 30738 9088 30744
rect 9140 29646 9168 31214
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 8772 28014 8800 29106
rect 9036 29028 9088 29034
rect 9036 28970 9088 28976
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 9048 27878 9076 28970
rect 9140 28422 9168 29242
rect 9232 29170 9260 33458
rect 10048 33244 10100 33250
rect 10048 33186 10100 33192
rect 9496 32904 9548 32910
rect 9496 32846 9548 32852
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9416 31249 9444 31282
rect 9402 31240 9458 31249
rect 9402 31175 9458 31184
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9140 28218 9168 28358
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8668 26512 8720 26518
rect 8668 26454 8720 26460
rect 8220 25996 8340 26024
rect 8404 26404 8524 26432
rect 8220 25906 8248 25996
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 7840 25764 7892 25770
rect 7840 25706 7892 25712
rect 8116 25764 8168 25770
rect 8116 25706 8168 25712
rect 7852 25226 7880 25706
rect 7932 25696 7984 25702
rect 8128 25673 8156 25706
rect 7932 25638 7984 25644
rect 8114 25664 8170 25673
rect 7944 25294 7972 25638
rect 8114 25599 8170 25608
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 8220 25158 8248 25434
rect 8404 25158 8432 26404
rect 8956 26353 8984 26862
rect 8942 26344 8998 26353
rect 8942 26279 8998 26288
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8588 26042 8616 26182
rect 8758 26072 8814 26081
rect 8576 26036 8628 26042
rect 8758 26007 8814 26016
rect 8576 25978 8628 25984
rect 8772 25906 8800 26007
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8588 25362 8616 25774
rect 8772 25498 8800 25842
rect 9048 25838 9076 27814
rect 9140 27470 9168 28154
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 27130 9168 27406
rect 9232 27334 9260 28018
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9126 26480 9182 26489
rect 9126 26415 9128 26424
rect 9180 26415 9182 26424
rect 9128 26386 9180 26392
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8760 25220 8812 25226
rect 8760 25162 8812 25168
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7852 24410 7880 24890
rect 7930 24712 7986 24721
rect 7930 24647 7932 24656
rect 7984 24647 7986 24656
rect 7932 24618 7984 24624
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7852 23118 7880 23598
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7944 23186 7972 23462
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7484 19242 7512 19314
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7484 18766 7512 18906
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7576 17785 7604 20402
rect 7668 20040 7696 21626
rect 7760 21554 7788 22510
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 8312 21350 8340 24074
rect 8404 24070 8432 25094
rect 8496 24886 8524 25094
rect 8772 24954 8800 25162
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 8864 24682 8892 24822
rect 8852 24676 8904 24682
rect 8852 24618 8904 24624
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8404 23322 8432 23598
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8404 22234 8432 23258
rect 8496 23225 8524 24006
rect 8588 23662 8616 24346
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8588 23497 8616 23598
rect 8574 23488 8630 23497
rect 8574 23423 8630 23432
rect 8482 23216 8538 23225
rect 8482 23151 8538 23160
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8496 22094 8524 23151
rect 8404 22066 8524 22094
rect 8404 22030 8432 22066
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 20058 7880 20198
rect 8312 20058 8340 20810
rect 8404 20058 8432 20878
rect 8496 20777 8524 21966
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8482 20768 8538 20777
rect 8482 20703 8538 20712
rect 7840 20052 7892 20058
rect 7668 20012 7788 20040
rect 7654 19952 7710 19961
rect 7654 19887 7710 19896
rect 7668 19378 7696 19887
rect 7760 19496 7788 20012
rect 7840 19994 7892 20000
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 7760 19468 7880 19496
rect 7746 19408 7802 19417
rect 7656 19372 7708 19378
rect 7746 19343 7802 19352
rect 7656 19314 7708 19320
rect 7562 17776 7618 17785
rect 7472 17740 7524 17746
rect 7562 17711 7618 17720
rect 7472 17682 7524 17688
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7010 16079 7066 16088
rect 7104 16108 7156 16114
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 14482 6960 15846
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6932 13394 6960 14418
rect 7024 14278 7052 16079
rect 7104 16050 7156 16056
rect 7208 15162 7236 16730
rect 7484 16504 7512 17682
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7576 16794 7604 17206
rect 7668 17184 7696 19314
rect 7760 18970 7788 19343
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7852 18902 7880 19468
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 8220 18766 8248 19110
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18193 7788 18566
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8128 18290 8156 18362
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 7746 18184 7802 18193
rect 7746 18119 7802 18128
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7760 17678 7788 18022
rect 7852 17814 7880 18022
rect 8312 17882 8340 19207
rect 8588 18426 8616 20878
rect 8680 20874 8708 24550
rect 8772 24313 8800 24550
rect 8758 24304 8814 24313
rect 8758 24239 8814 24248
rect 8852 24268 8904 24274
rect 8852 24210 8904 24216
rect 8864 23730 8892 24210
rect 9048 24206 9076 24550
rect 9140 24206 9168 25910
rect 9232 25294 9260 26726
rect 9324 26246 9352 27066
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9324 24954 9352 25910
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9128 24200 9180 24206
rect 9180 24160 9260 24188
rect 9128 24142 9180 24148
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8864 22098 8892 23666
rect 9126 23080 9182 23089
rect 9126 23015 9182 23024
rect 9140 22982 9168 23015
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8772 20618 8800 21490
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8680 20590 8800 20618
rect 8680 19786 8708 20590
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8864 20262 8892 20334
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 19825 8892 20198
rect 8850 19816 8906 19825
rect 8668 19780 8720 19786
rect 8850 19751 8906 19760
rect 8668 19722 8720 19728
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7852 17678 7880 17750
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 8116 17196 8168 17202
rect 7668 17156 7972 17184
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7668 16590 7696 17002
rect 7944 16590 7972 17156
rect 8312 17184 8340 17546
rect 8404 17202 8432 17818
rect 8496 17678 8524 18226
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8168 17156 8340 17184
rect 8392 17196 8444 17202
rect 8116 17138 8168 17144
rect 8392 17138 8444 17144
rect 8128 17105 8156 17138
rect 8114 17096 8170 17105
rect 8114 17031 8170 17040
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16726 8340 16934
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 7656 16584 7708 16590
rect 7932 16584 7984 16590
rect 7656 16526 7708 16532
rect 7746 16552 7802 16561
rect 7564 16516 7616 16522
rect 7484 16476 7564 16504
rect 7932 16526 7984 16532
rect 7746 16487 7748 16496
rect 7564 16458 7616 16464
rect 7800 16487 7802 16496
rect 7748 16458 7800 16464
rect 7562 16280 7618 16289
rect 7562 16215 7618 16224
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7196 14408 7248 14414
rect 7300 14396 7328 16050
rect 7576 16046 7604 16215
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7562 15600 7618 15609
rect 7248 14368 7328 14396
rect 7196 14350 7248 14356
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7024 13705 7052 13738
rect 7010 13696 7066 13705
rect 7010 13631 7066 13640
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6918 13288 6974 13297
rect 6918 13223 6974 13232
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6932 12730 6960 13223
rect 6840 12702 6960 12730
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6656 12406 6776 12434
rect 6552 12378 6604 12384
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6458 12064 6514 12073
rect 6458 11999 6514 12008
rect 6472 11762 6500 11999
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11286 6500 11698
rect 6656 11626 6684 12174
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6288 11070 6408 11098
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6184 8016 6236 8022
rect 6182 7984 6184 7993
rect 6236 7984 6238 7993
rect 6182 7919 6238 7928
rect 6288 7546 6316 11070
rect 6472 8906 6500 11222
rect 6564 11218 6592 11494
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 9761 6592 11018
rect 6550 9752 6606 9761
rect 6550 9687 6606 9696
rect 6564 9654 6592 9687
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6656 8974 6684 11562
rect 6748 10674 6776 12406
rect 6840 12306 6868 12702
rect 6918 12472 6974 12481
rect 6918 12407 6974 12416
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 12209 6868 12242
rect 6826 12200 6882 12209
rect 6826 12135 6882 12144
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6736 10056 6788 10062
rect 6840 10044 6868 11698
rect 6932 10674 6960 12407
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6932 10062 6960 10610
rect 6788 10016 6868 10044
rect 6920 10056 6972 10062
rect 6736 9998 6788 10004
rect 6920 9998 6972 10004
rect 6748 8974 6776 9998
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9178 6868 9862
rect 6932 9722 6960 9998
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7024 9042 7052 11630
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6182 6352 6238 6361
rect 6182 6287 6238 6296
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 5234 6132 5646
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6196 3602 6224 6287
rect 6288 4214 6316 7482
rect 6380 7188 6408 8230
rect 6472 7342 6500 8842
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6380 7160 6500 7188
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6380 6458 6408 6598
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6288 3398 6316 4150
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 6380 1562 6408 6394
rect 6472 6254 6500 7160
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4146 6500 4966
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6564 3670 6592 7754
rect 6656 7410 6684 8910
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6748 7274 6776 8910
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6932 8498 6960 8774
rect 7024 8498 7052 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 7546 7052 8434
rect 7116 8090 7144 14350
rect 7208 13977 7236 14350
rect 7194 13968 7250 13977
rect 7194 13903 7250 13912
rect 7392 13326 7420 15574
rect 7562 15535 7618 15544
rect 7470 15192 7526 15201
rect 7576 15162 7604 15535
rect 7470 15127 7526 15136
rect 7564 15156 7616 15162
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12753 7328 13126
rect 7484 12986 7512 15127
rect 7564 15098 7616 15104
rect 7760 14634 7788 16458
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8312 16114 8340 16662
rect 8404 16182 8432 17138
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8404 16028 8432 16118
rect 8404 16000 8616 16028
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8220 15366 8248 15914
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15638 8340 15846
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8300 15496 8352 15502
rect 8352 15444 8432 15450
rect 8300 15438 8432 15444
rect 8312 15422 8432 15438
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7760 14606 7880 14634
rect 8036 14618 8064 14758
rect 7852 14550 7880 14606
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7576 13841 7604 13942
rect 7562 13832 7618 13841
rect 7562 13767 7618 13776
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7286 12744 7342 12753
rect 7286 12679 7342 12688
rect 7286 12472 7342 12481
rect 7286 12407 7342 12416
rect 7300 12374 7328 12407
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7208 12073 7236 12174
rect 7194 12064 7250 12073
rect 7194 11999 7250 12008
rect 7300 11762 7328 12174
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7194 10704 7250 10713
rect 7194 10639 7196 10648
rect 7248 10639 7250 10648
rect 7196 10610 7248 10616
rect 7208 9994 7236 10610
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7300 9654 7328 11290
rect 7392 10266 7420 12786
rect 7564 12776 7616 12782
rect 7562 12744 7564 12753
rect 7616 12744 7618 12753
rect 7562 12679 7618 12688
rect 7668 12617 7696 13262
rect 7654 12608 7710 12617
rect 7654 12543 7710 12552
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7668 11830 7696 12310
rect 7760 11880 7788 14486
rect 8220 14385 8248 15098
rect 8404 15026 8432 15422
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8206 14376 8262 14385
rect 8206 14311 8262 14320
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 7852 13394 7880 14010
rect 7930 13968 7986 13977
rect 8220 13938 8248 14010
rect 7930 13903 7932 13912
rect 7984 13903 7986 13912
rect 8208 13932 8260 13938
rect 7932 13874 7984 13880
rect 8208 13874 8260 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13433 8064 13806
rect 8022 13424 8078 13433
rect 7840 13388 7892 13394
rect 8022 13359 8078 13368
rect 7840 13330 7892 13336
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12238 7880 12582
rect 8220 12434 8248 12650
rect 8128 12406 8248 12434
rect 8128 12374 8156 12406
rect 8116 12368 8168 12374
rect 8208 12368 8260 12374
rect 8116 12310 8168 12316
rect 8206 12336 8208 12345
rect 8260 12336 8262 12345
rect 8206 12271 8262 12280
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8312 12170 8340 14962
rect 8404 12918 8432 14962
rect 8496 13326 8524 15642
rect 8588 15502 8616 16000
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12986 8524 13262
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12374 8432 12582
rect 8392 12368 8444 12374
rect 8588 12322 8616 14894
rect 8680 14618 8708 19722
rect 8956 19378 8984 21286
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8852 18896 8904 18902
rect 8758 18864 8814 18873
rect 8852 18838 8904 18844
rect 8758 18799 8814 18808
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8680 13569 8708 14554
rect 8772 14278 8800 18799
rect 8864 18290 8892 18838
rect 8956 18698 8984 19314
rect 9048 18873 9076 22578
rect 9232 19854 9260 24160
rect 9324 23662 9352 24754
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9310 23352 9366 23361
rect 9310 23287 9366 23296
rect 9324 23186 9352 23287
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9324 22681 9352 23122
rect 9310 22672 9366 22681
rect 9310 22607 9366 22616
rect 9416 22137 9444 26862
rect 9508 26042 9536 32846
rect 9956 32564 10008 32570
rect 9956 32506 10008 32512
rect 9588 32496 9640 32502
rect 9588 32438 9640 32444
rect 9600 31754 9628 32438
rect 9588 31748 9640 31754
rect 9588 31690 9640 31696
rect 9968 30938 9996 32506
rect 10060 31822 10088 33186
rect 10416 33176 10468 33182
rect 10416 33118 10468 33124
rect 10140 32292 10192 32298
rect 10140 32234 10192 32240
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 10152 31414 10180 32234
rect 10428 31822 10456 33118
rect 12532 32972 12584 32978
rect 12532 32914 12584 32920
rect 11704 32768 11756 32774
rect 11704 32710 11756 32716
rect 11612 32496 11664 32502
rect 11612 32438 11664 32444
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 10600 31952 10652 31958
rect 10506 31920 10562 31929
rect 10600 31894 10652 31900
rect 10506 31855 10508 31864
rect 10560 31855 10562 31864
rect 10508 31826 10560 31832
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10508 31680 10560 31686
rect 10508 31622 10560 31628
rect 10140 31408 10192 31414
rect 10140 31350 10192 31356
rect 9956 30932 10008 30938
rect 9956 30874 10008 30880
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9600 27402 9628 29990
rect 9692 28694 9720 30670
rect 9968 30394 9996 30874
rect 10152 30734 10180 31350
rect 10232 31136 10284 31142
rect 10232 31078 10284 31084
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10138 30424 10194 30433
rect 9956 30388 10008 30394
rect 10138 30359 10194 30368
rect 9956 30330 10008 30336
rect 10152 30326 10180 30359
rect 10140 30320 10192 30326
rect 10140 30262 10192 30268
rect 9772 30184 9824 30190
rect 9772 30126 9824 30132
rect 9680 28688 9732 28694
rect 9680 28630 9732 28636
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9586 26616 9642 26625
rect 9586 26551 9588 26560
rect 9640 26551 9642 26560
rect 9588 26522 9640 26528
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9508 25294 9536 25774
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9402 22128 9458 22137
rect 9402 22063 9458 22072
rect 9508 22094 9536 24754
rect 9600 24410 9628 25774
rect 9692 25702 9720 28426
rect 9784 27878 9812 30126
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9784 27674 9812 27814
rect 9772 27668 9824 27674
rect 9772 27610 9824 27616
rect 9876 27538 9904 28494
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9864 27532 9916 27538
rect 9864 27474 9916 27480
rect 9876 26450 9904 27474
rect 9864 26444 9916 26450
rect 9864 26386 9916 26392
rect 9968 26382 9996 27814
rect 10048 27668 10100 27674
rect 10048 27610 10100 27616
rect 10060 27470 10088 27610
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9784 25809 9812 25978
rect 9770 25800 9826 25809
rect 9770 25735 9826 25744
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9586 24168 9642 24177
rect 9586 24103 9588 24112
rect 9640 24103 9642 24112
rect 9588 24074 9640 24080
rect 9692 24018 9720 25162
rect 9600 23990 9720 24018
rect 9600 23526 9628 23990
rect 9784 23730 9812 25298
rect 9876 23866 9904 25978
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9772 23588 9824 23594
rect 9772 23530 9824 23536
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9600 22982 9628 23462
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9692 22642 9720 23258
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9508 22066 9628 22094
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9324 21010 9352 21830
rect 9402 21448 9458 21457
rect 9402 21383 9404 21392
rect 9456 21383 9458 21392
rect 9404 21354 9456 21360
rect 9508 21350 9536 21830
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9496 21072 9548 21078
rect 9600 21060 9628 22066
rect 9692 21418 9720 22578
rect 9784 21962 9812 23530
rect 9876 22030 9904 23598
rect 9968 22438 9996 26318
rect 10060 25294 10088 27406
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 23905 10088 24686
rect 10046 23896 10102 23905
rect 10046 23831 10102 23840
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9680 21072 9732 21078
rect 9600 21032 9680 21060
rect 9496 21014 9548 21020
rect 9680 21014 9732 21020
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9034 18864 9090 18873
rect 9034 18799 9090 18808
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 9034 18320 9090 18329
rect 8852 18284 8904 18290
rect 9034 18255 9090 18264
rect 8852 18226 8904 18232
rect 8864 18086 8892 18226
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8864 17542 8892 18022
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8864 16250 8892 16594
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8956 15978 8984 17138
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8850 15464 8906 15473
rect 8850 15399 8906 15408
rect 8864 15162 8892 15399
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13841 8800 13874
rect 8758 13832 8814 13841
rect 8758 13767 8814 13776
rect 8666 13560 8722 13569
rect 8666 13495 8722 13504
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12782 8708 13262
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12850 8800 13126
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8864 12646 8892 14758
rect 8956 12986 8984 15302
rect 9048 15162 9076 18255
rect 9140 18057 9168 19314
rect 9232 18766 9260 19314
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9126 18048 9182 18057
rect 9126 17983 9182 17992
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9140 16590 9168 17138
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9232 16402 9260 17274
rect 9140 16374 9260 16402
rect 9140 16114 9168 16374
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 13297 9076 14418
rect 9232 14278 9260 14826
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9034 13288 9090 13297
rect 9034 13223 9090 13232
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12640 8904 12646
rect 8666 12608 8722 12617
rect 8852 12582 8904 12588
rect 8666 12543 8722 12552
rect 8392 12310 8444 12316
rect 8496 12294 8616 12322
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 7760 11852 7880 11880
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 10742 7512 11494
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 9178 7328 9590
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7484 8548 7512 9862
rect 7576 8838 7604 11222
rect 7668 10062 7696 11766
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 10266 7788 11698
rect 7852 11626 7880 11852
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8220 11064 8248 11562
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11218 8340 11494
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8220 11036 8340 11064
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 8312 10792 8340 11036
rect 8220 10764 8340 10792
rect 7840 10464 7892 10470
rect 7838 10432 7840 10441
rect 7892 10432 7894 10441
rect 7838 10367 7894 10376
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7654 9888 7710 9897
rect 7654 9823 7710 9832
rect 7668 9217 7696 9823
rect 7654 9208 7710 9217
rect 7760 9178 7788 10202
rect 8220 10130 8248 10764
rect 8404 10266 8432 12174
rect 8496 11830 8524 12294
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 7930 9616 7986 9625
rect 7930 9551 7932 9560
rect 7984 9551 7986 9560
rect 7932 9522 7984 9528
rect 7654 9143 7710 9152
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8312 9110 8340 9930
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7392 8520 7512 8548
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7392 7993 7420 8520
rect 7576 8480 7604 8774
rect 7484 8452 7604 8480
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6920 7472 6972 7478
rect 6918 7440 6920 7449
rect 7288 7472 7340 7478
rect 6972 7440 6974 7449
rect 7288 7414 7340 7420
rect 6918 7375 6974 7384
rect 6918 7304 6974 7313
rect 6736 7268 6788 7274
rect 6918 7239 6974 7248
rect 6736 7210 6788 7216
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5914 6776 6258
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6734 5536 6790 5545
rect 6734 5471 6790 5480
rect 6642 5264 6698 5273
rect 6748 5234 6776 5471
rect 6642 5199 6644 5208
rect 6696 5199 6698 5208
rect 6736 5228 6788 5234
rect 6644 5170 6696 5176
rect 6736 5170 6788 5176
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6564 3126 6592 3606
rect 6656 3602 6684 5034
rect 6840 4622 6868 6598
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3670 6776 3878
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6840 3482 6868 4150
rect 6932 3534 6960 7239
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 6118 7236 6734
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7010 5944 7066 5953
rect 7010 5879 7066 5888
rect 7024 5574 7052 5879
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7024 3942 7052 4558
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6748 3454 6868 3482
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6564 2650 6592 2926
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6564 1970 6592 2586
rect 6656 2038 6684 3402
rect 6748 2854 6776 3454
rect 7024 3058 7052 3878
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6644 2032 6696 2038
rect 6644 1974 6696 1980
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6368 1556 6420 1562
rect 6368 1498 6420 1504
rect 6748 1358 6776 2790
rect 7024 2446 7052 2994
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7024 1952 7052 2382
rect 7116 2106 7144 4490
rect 7208 2378 7236 5714
rect 7300 3670 7328 7414
rect 7392 6322 7420 7686
rect 7484 7410 7512 8452
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 4729 7420 6054
rect 7378 4720 7434 4729
rect 7378 4655 7434 4664
rect 7484 4214 7512 6802
rect 7576 5710 7604 8298
rect 7668 7410 7696 8910
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 8312 8362 8340 8774
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8022 7880 8230
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6322 7696 7142
rect 7760 6798 7788 7686
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8404 7562 8432 10066
rect 8496 10062 8524 11766
rect 8588 11014 8616 12174
rect 8680 11898 8708 12543
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8680 10674 8708 11154
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9722 8616 9998
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 8362 8524 8502
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8312 7534 8432 7562
rect 8312 7528 8340 7534
rect 8220 7500 8340 7528
rect 8116 7336 8168 7342
rect 8114 7304 8116 7313
rect 8168 7304 8170 7313
rect 8114 7239 8170 7248
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7748 6656 7800 6662
rect 8220 6644 8248 7500
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7002 8432 7346
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8220 6616 8340 6644
rect 7748 6598 7800 6604
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7484 3126 7512 3878
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7104 1964 7156 1970
rect 7024 1924 7104 1952
rect 7104 1906 7156 1912
rect 7392 1834 7420 2586
rect 7668 2038 7696 5510
rect 7760 4554 7788 6598
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8312 6372 8340 6616
rect 8404 6458 8432 6666
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8220 6344 8340 6372
rect 8220 5846 8248 6344
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8220 5624 8248 5782
rect 8220 5596 8340 5624
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8312 5352 8340 5596
rect 8220 5324 8340 5352
rect 8220 4570 8248 5324
rect 7748 4548 7800 4554
rect 8220 4542 8340 4570
rect 7748 4490 7800 4496
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 7748 4208 7800 4214
rect 8312 4196 8340 4542
rect 8404 4486 8432 5782
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 7748 4150 7800 4156
rect 8220 4168 8340 4196
rect 7656 2032 7708 2038
rect 7656 1974 7708 1980
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 7760 1222 7788 4150
rect 8220 3942 8248 4168
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 8206 2544 8262 2553
rect 8206 2479 8262 2488
rect 8220 2446 8248 2479
rect 8208 2440 8260 2446
rect 8496 2394 8524 7210
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6798 8616 7142
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 4826 8616 5578
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8680 4758 8708 10610
rect 8772 9518 8800 10678
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 8090 8800 9454
rect 8864 9382 8892 12407
rect 8956 12102 8984 12922
rect 9036 12640 9088 12646
rect 9034 12608 9036 12617
rect 9088 12608 9090 12617
rect 9034 12543 9090 12552
rect 9140 12434 9168 14214
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 13977 9260 14010
rect 9218 13968 9274 13977
rect 9218 13903 9274 13912
rect 9324 13734 9352 20810
rect 9402 20088 9458 20097
rect 9402 20023 9458 20032
rect 9416 19378 9444 20023
rect 9508 19718 9536 21014
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9416 17649 9444 19178
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18290 9536 19110
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9402 17640 9458 17649
rect 9402 17575 9458 17584
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9324 13512 9352 13670
rect 9232 13484 9352 13512
rect 9232 12850 9260 13484
rect 9310 13424 9366 13433
rect 9310 13359 9366 13368
rect 9324 13326 9352 13359
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9416 12481 9444 16390
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 14618 9536 15846
rect 9600 15434 9628 20742
rect 9692 18970 9720 20878
rect 9876 20466 9904 21966
rect 9954 21720 10010 21729
rect 9954 21655 9956 21664
rect 10008 21655 10010 21664
rect 9956 21626 10008 21632
rect 9956 21412 10008 21418
rect 9956 21354 10008 21360
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9770 20360 9826 20369
rect 9770 20295 9772 20304
rect 9824 20295 9826 20304
rect 9772 20266 9824 20272
rect 9968 19922 9996 21354
rect 10060 21146 10088 23598
rect 10152 22710 10180 29446
rect 10244 27130 10272 31078
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10336 26466 10364 26862
rect 10244 26438 10364 26466
rect 10244 23662 10272 26438
rect 10428 26382 10456 31078
rect 10520 29034 10548 31622
rect 10612 31142 10640 31894
rect 10692 31816 10744 31822
rect 10692 31758 10744 31764
rect 10600 31136 10652 31142
rect 10600 31078 10652 31084
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10508 29028 10560 29034
rect 10508 28970 10560 28976
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10336 23100 10364 26250
rect 10520 26217 10548 28970
rect 10506 26208 10562 26217
rect 10506 26143 10562 26152
rect 10508 25900 10560 25906
rect 10508 25842 10560 25848
rect 10520 25673 10548 25842
rect 10506 25664 10562 25673
rect 10506 25599 10562 25608
rect 10612 25498 10640 30670
rect 10704 30326 10732 31758
rect 10692 30320 10744 30326
rect 10692 30262 10744 30268
rect 11164 30054 11192 32370
rect 11624 32230 11652 32438
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11369 32124 11677 32133
rect 11369 32122 11375 32124
rect 11431 32122 11455 32124
rect 11511 32122 11535 32124
rect 11591 32122 11615 32124
rect 11671 32122 11677 32124
rect 11431 32070 11433 32122
rect 11613 32070 11615 32122
rect 11369 32068 11375 32070
rect 11431 32068 11455 32070
rect 11511 32068 11535 32070
rect 11591 32068 11615 32070
rect 11671 32068 11677 32070
rect 11369 32059 11677 32068
rect 11716 31482 11744 32710
rect 12544 32298 12572 32914
rect 12440 32292 12492 32298
rect 12440 32234 12492 32240
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 11978 32192 12034 32201
rect 11978 32127 12034 32136
rect 11794 31512 11850 31521
rect 11704 31476 11756 31482
rect 11794 31447 11850 31456
rect 11704 31418 11756 31424
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 11808 30977 11836 31447
rect 11794 30968 11850 30977
rect 11794 30903 11850 30912
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11716 30190 11744 30534
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11992 30122 12020 32127
rect 12452 31346 12480 32234
rect 12820 32230 12848 33526
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13176 32904 13228 32910
rect 13176 32846 13228 32852
rect 12808 32224 12860 32230
rect 12808 32166 12860 32172
rect 13188 31958 13216 32846
rect 13636 32428 13688 32434
rect 13636 32370 13688 32376
rect 13268 32360 13320 32366
rect 13268 32302 13320 32308
rect 13176 31952 13228 31958
rect 13176 31894 13228 31900
rect 13280 31754 13308 32302
rect 13544 32292 13596 32298
rect 13544 32234 13596 32240
rect 13452 31816 13504 31822
rect 13452 31758 13504 31764
rect 13268 31748 13320 31754
rect 13268 31690 13320 31696
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 13096 30870 13124 31214
rect 13084 30864 13136 30870
rect 13084 30806 13136 30812
rect 12728 30666 12940 30682
rect 12716 30660 12952 30666
rect 12768 30654 12900 30660
rect 12716 30602 12768 30608
rect 12900 30602 12952 30608
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 12164 30388 12216 30394
rect 12164 30330 12216 30336
rect 12084 30258 12112 30330
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12176 30138 12204 30330
rect 13096 30326 13124 30806
rect 13084 30320 13136 30326
rect 13084 30262 13136 30268
rect 11980 30116 12032 30122
rect 11980 30058 12032 30064
rect 12084 30110 12204 30138
rect 10692 30048 10744 30054
rect 10690 30016 10692 30025
rect 11152 30048 11204 30054
rect 10744 30016 10746 30025
rect 11152 29990 11204 29996
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 10690 29951 10746 29960
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 10692 29028 10744 29034
rect 10692 28970 10744 28976
rect 10704 28121 10732 28970
rect 10968 28688 11020 28694
rect 10968 28630 11020 28636
rect 10980 28422 11008 28630
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10690 28112 10746 28121
rect 10690 28047 10746 28056
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10796 26586 10824 27338
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10416 25424 10468 25430
rect 10468 25384 10548 25412
rect 10416 25366 10468 25372
rect 10520 25158 10548 25384
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10428 24954 10456 25094
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10520 24342 10548 24754
rect 10612 24342 10640 24754
rect 10508 24336 10560 24342
rect 10508 24278 10560 24284
rect 10600 24336 10652 24342
rect 10600 24278 10652 24284
rect 10508 24200 10560 24206
rect 10612 24188 10640 24278
rect 10560 24160 10640 24188
rect 10508 24142 10560 24148
rect 10506 24032 10562 24041
rect 10506 23967 10562 23976
rect 10520 23526 10548 23967
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10506 23216 10562 23225
rect 10506 23151 10562 23160
rect 10416 23112 10468 23118
rect 10336 23072 10416 23100
rect 10416 23054 10468 23060
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10336 22778 10364 22918
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10152 22094 10180 22646
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10152 22066 10272 22094
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19514 9996 19858
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9784 19145 9812 19382
rect 9770 19136 9826 19145
rect 9770 19071 9826 19080
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9770 18592 9826 18601
rect 9770 18527 9826 18536
rect 9784 18290 9812 18527
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17066 9720 17614
rect 9784 17338 9812 18226
rect 9876 17814 9904 18770
rect 9864 17808 9916 17814
rect 9862 17776 9864 17785
rect 9916 17776 9918 17785
rect 9862 17711 9918 17720
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9876 17542 9904 17614
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16590 9720 17002
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 15502 9720 16526
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 14006 9536 14214
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9600 13938 9628 15263
rect 9692 14890 9720 15438
rect 9784 15026 9812 17138
rect 9876 16425 9904 17478
rect 9968 17202 9996 17546
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9968 16522 9996 17138
rect 10060 17134 10088 20742
rect 10152 20466 10180 21966
rect 10244 21350 10272 22066
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10336 21128 10364 22102
rect 10244 21100 10364 21128
rect 10244 20534 10272 21100
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 18290 10180 18566
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10152 16998 10180 18226
rect 10244 17241 10272 20198
rect 10336 19310 10364 20946
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18290 10364 18906
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10322 17776 10378 17785
rect 10428 17746 10456 23054
rect 10520 22982 10548 23151
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10612 20913 10640 23802
rect 10704 23118 10732 26318
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 10796 24954 10824 26182
rect 10980 25906 11008 27950
rect 11072 27441 11100 29786
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11164 27577 11192 28562
rect 11256 28014 11284 29582
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11716 27674 11744 28086
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 11150 27568 11206 27577
rect 11150 27503 11206 27512
rect 11244 27464 11296 27470
rect 11058 27432 11114 27441
rect 11244 27406 11296 27412
rect 11058 27367 11114 27376
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 10968 25900 11020 25906
rect 10888 25860 10968 25888
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10796 24206 10824 24686
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10796 23254 10824 23734
rect 10888 23322 10916 25860
rect 10968 25842 11020 25848
rect 10968 25696 11020 25702
rect 11072 25673 11100 26250
rect 11164 26042 11192 26930
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 11152 25764 11204 25770
rect 11152 25706 11204 25712
rect 10968 25638 11020 25644
rect 11058 25664 11114 25673
rect 10980 25430 11008 25638
rect 11058 25599 11114 25608
rect 11058 25528 11114 25537
rect 11058 25463 11114 25472
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 11072 25226 11100 25463
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10980 24818 11008 25162
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10704 22710 10732 23054
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10692 22500 10744 22506
rect 10692 22442 10744 22448
rect 10704 21690 10732 22442
rect 10796 22234 10824 23190
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10782 21720 10838 21729
rect 10692 21684 10744 21690
rect 10782 21655 10784 21664
rect 10692 21626 10744 21632
rect 10836 21655 10838 21664
rect 10784 21626 10836 21632
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10704 21350 10732 21490
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10796 21010 10824 21490
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10598 20904 10654 20913
rect 10598 20839 10654 20848
rect 10612 18834 10640 20839
rect 10796 20806 10824 20946
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10704 19378 10732 20266
rect 10796 19514 10824 20266
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10784 19304 10836 19310
rect 10782 19272 10784 19281
rect 10836 19272 10838 19281
rect 10782 19207 10838 19216
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10520 17814 10548 18702
rect 10704 18630 10732 19110
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10322 17711 10324 17720
rect 10376 17711 10378 17720
rect 10416 17740 10468 17746
rect 10324 17682 10376 17688
rect 10416 17682 10468 17688
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10230 17232 10286 17241
rect 10230 17167 10286 17176
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 10048 16448 10100 16454
rect 9862 16416 9918 16425
rect 9862 16351 9918 16360
rect 10046 16416 10048 16425
rect 10100 16416 10102 16425
rect 10046 16351 10102 16360
rect 10046 16144 10102 16153
rect 10046 16079 10102 16088
rect 10060 16046 10088 16079
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9784 14770 9812 14962
rect 9692 14742 9812 14770
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9494 13560 9550 13569
rect 9494 13495 9550 13504
rect 9508 13462 9536 13495
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9048 12406 9168 12434
rect 9402 12472 9458 12481
rect 9402 12407 9458 12416
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8942 11792 8998 11801
rect 8942 11727 8944 11736
rect 8996 11727 8998 11736
rect 8944 11698 8996 11704
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11393 8984 11494
rect 8942 11384 8998 11393
rect 8942 11319 8998 11328
rect 8956 9994 8984 11319
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8864 8362 8892 9046
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8772 7818 8800 8026
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8772 5710 8800 6938
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8772 4146 8800 5646
rect 8864 5302 8892 8298
rect 8956 6390 8984 9687
rect 9048 8974 9076 12406
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11121 9168 12038
rect 9126 11112 9182 11121
rect 9126 11047 9182 11056
rect 9232 10577 9260 12242
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11665 9352 11698
rect 9310 11656 9366 11665
rect 9310 11591 9366 11600
rect 9218 10568 9274 10577
rect 9218 10503 9274 10512
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8566 9076 8910
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4146 8892 4966
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8680 3602 8708 3878
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8208 2382 8260 2388
rect 8404 2366 8524 2394
rect 8404 2310 8432 2366
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 8956 1970 8984 6054
rect 9048 3534 9076 7482
rect 9140 7342 9168 8026
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6254 9168 7278
rect 9232 7002 9260 10134
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6458 9260 6734
rect 9324 6730 9352 11591
rect 9402 11248 9458 11257
rect 9402 11183 9458 11192
rect 9416 11082 9444 11183
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9404 9648 9456 9654
rect 9402 9616 9404 9625
rect 9456 9616 9458 9625
rect 9402 9551 9458 9560
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 8566 9444 8842
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5846 9168 6190
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9140 5710 9168 5782
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 5234 9168 5646
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9324 5098 9352 6394
rect 9416 6089 9444 7822
rect 9508 7206 9536 13262
rect 9600 12170 9628 13398
rect 9692 12850 9720 14742
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9784 12073 9812 13806
rect 9876 13530 9904 15302
rect 9968 13705 9996 15506
rect 10152 14074 10180 16934
rect 10336 16794 10364 17274
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10230 16552 10286 16561
rect 10230 16487 10232 16496
rect 10284 16487 10286 16496
rect 10232 16458 10284 16464
rect 10244 16250 10272 16458
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10244 15026 10272 16186
rect 10336 15910 10364 16730
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10428 15570 10456 16186
rect 10520 16114 10548 17750
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10612 14822 10640 18362
rect 10704 18086 10732 18566
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 17814 10732 18022
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10704 16658 10732 17750
rect 10796 17066 10824 18634
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10704 16454 10732 16594
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10782 16416 10838 16425
rect 10704 16046 10732 16390
rect 10782 16351 10838 16360
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10796 15858 10824 16351
rect 10888 16250 10916 22578
rect 10980 22166 11008 24346
rect 11072 23662 11100 24822
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 11072 23186 11100 23598
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10980 22030 11008 22102
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11164 21622 11192 25706
rect 11256 23866 11284 27406
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11440 26042 11468 26182
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11348 24614 11376 24890
rect 11518 24712 11574 24721
rect 11518 24647 11574 24656
rect 11532 24614 11560 24647
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11348 23746 11376 24142
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11624 24041 11652 24074
rect 11610 24032 11666 24041
rect 11610 23967 11666 23976
rect 11256 23718 11376 23746
rect 11256 23254 11284 23718
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11244 23248 11296 23254
rect 11244 23190 11296 23196
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11072 21350 11100 21558
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 11060 21344 11112 21350
rect 11348 21332 11376 22170
rect 11716 21554 11744 27270
rect 11808 24070 11836 29990
rect 11886 29880 11942 29889
rect 11886 29815 11942 29824
rect 11980 29844 12032 29850
rect 11900 29510 11928 29815
rect 11980 29786 12032 29792
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11992 28994 12020 29786
rect 12084 29238 12112 30110
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 11992 28966 12112 28994
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11900 28218 11928 28494
rect 11888 28212 11940 28218
rect 11888 28154 11940 28160
rect 12084 27826 12112 28966
rect 12176 28626 12204 29106
rect 12268 28937 12296 29514
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12254 28928 12310 28937
rect 12254 28863 12310 28872
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12360 28558 12388 29038
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12254 27840 12310 27849
rect 12084 27798 12204 27826
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11992 26586 12020 26794
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11900 24206 11928 26454
rect 12084 24698 12112 27610
rect 12176 24954 12204 27798
rect 12254 27775 12310 27784
rect 12268 25770 12296 27775
rect 12360 27470 12388 28494
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12360 26994 12388 27406
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12256 25764 12308 25770
rect 12256 25706 12308 25712
rect 12164 24948 12216 24954
rect 12216 24908 12296 24936
rect 12164 24890 12216 24896
rect 12084 24670 12204 24698
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 11794 23352 11850 23361
rect 11794 23287 11796 23296
rect 11848 23287 11850 23296
rect 11796 23258 11848 23264
rect 11900 23202 11928 23598
rect 11808 23174 11928 23202
rect 11808 22778 11836 23174
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11796 21548 11848 21554
rect 11900 21536 11928 22918
rect 11848 21508 11928 21536
rect 11796 21490 11848 21496
rect 11060 21286 11112 21292
rect 11256 21304 11376 21332
rect 10980 17678 11008 21286
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11072 19417 11100 20334
rect 11058 19408 11114 19417
rect 11058 19343 11114 19352
rect 11072 19145 11100 19343
rect 11164 19310 11192 20402
rect 11256 19786 11284 21304
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 20777 11468 20810
rect 11426 20768 11482 20777
rect 11426 20703 11482 20712
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11716 20058 11744 21490
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11808 19938 11836 21490
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11716 19910 11836 19938
rect 11900 19922 11928 20470
rect 11992 20058 12020 23734
rect 12084 22982 12112 24210
rect 12176 23610 12204 24670
rect 12268 24206 12296 24908
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12176 23582 12296 23610
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12176 23118 12204 23258
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12268 23066 12296 23582
rect 12360 23186 12388 26386
rect 12544 25906 12572 29990
rect 12714 29336 12770 29345
rect 12714 29271 12770 29280
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 27606 12664 28358
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 12636 27470 12664 27542
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12728 27316 12756 29271
rect 13372 28801 13400 31282
rect 13464 30394 13492 31758
rect 13556 31686 13584 32234
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13648 30802 13676 32370
rect 13740 32230 13768 32982
rect 13728 32224 13780 32230
rect 13728 32166 13780 32172
rect 13832 31482 13860 33050
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13728 31136 13780 31142
rect 13726 31104 13728 31113
rect 13780 31104 13782 31113
rect 13726 31039 13782 31048
rect 13740 30938 13768 31039
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 13740 30802 13768 30874
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13452 30388 13504 30394
rect 13740 30376 13768 30738
rect 13452 30330 13504 30336
rect 13648 30348 13768 30376
rect 13648 29306 13676 30348
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13740 29753 13768 30194
rect 13726 29744 13782 29753
rect 13726 29679 13782 29688
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13636 29300 13688 29306
rect 13636 29242 13688 29248
rect 13648 29170 13676 29242
rect 13740 29170 13768 29582
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13358 28792 13414 28801
rect 13358 28727 13414 28736
rect 13648 28558 13676 29106
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13268 27940 13320 27946
rect 13268 27882 13320 27888
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12636 27288 12756 27316
rect 12808 27328 12860 27334
rect 12636 27130 12664 27288
rect 12808 27270 12860 27276
rect 12820 27130 12848 27270
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12820 26858 12848 27066
rect 12898 27024 12954 27033
rect 13188 26994 13216 27406
rect 12898 26959 12954 26968
rect 13176 26988 13228 26994
rect 12808 26852 12860 26858
rect 12808 26794 12860 26800
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12452 25294 12480 25774
rect 12544 25498 12572 25842
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12452 24954 12480 25094
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12452 23662 12480 24890
rect 12636 24818 12664 25230
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12440 23112 12492 23118
rect 12268 23050 12388 23066
rect 12440 23054 12492 23060
rect 12268 23044 12400 23050
rect 12268 23038 12348 23044
rect 12348 22986 12400 22992
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11888 19916 11940 19922
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11256 19310 11284 19450
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11256 19156 11284 19246
rect 11348 19174 11376 19858
rect 11610 19408 11666 19417
rect 11610 19343 11612 19352
rect 11664 19343 11666 19352
rect 11612 19314 11664 19320
rect 11058 19136 11114 19145
rect 11058 19071 11114 19080
rect 11164 19128 11284 19156
rect 11336 19168 11388 19174
rect 11072 18834 11100 19071
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18465 11100 18770
rect 11164 18630 11192 19128
rect 11336 19110 11388 19116
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11612 18896 11664 18902
rect 11518 18864 11574 18873
rect 11612 18838 11664 18844
rect 11518 18799 11520 18808
rect 11572 18799 11574 18808
rect 11520 18770 11572 18776
rect 11624 18766 11652 18838
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11152 18624 11204 18630
rect 11150 18592 11152 18601
rect 11428 18624 11480 18630
rect 11204 18592 11206 18601
rect 11428 18566 11480 18572
rect 11610 18592 11666 18601
rect 11150 18527 11206 18536
rect 11058 18456 11114 18465
rect 11058 18391 11114 18400
rect 11072 17678 11100 18391
rect 11440 18290 11468 18566
rect 11610 18527 11666 18536
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11624 18222 11652 18527
rect 11612 18216 11664 18222
rect 11610 18184 11612 18193
rect 11664 18184 11666 18193
rect 11610 18119 11666 18128
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10980 17270 11008 17614
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 11072 17202 11100 17614
rect 11440 17610 11468 17682
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11164 17270 11192 17546
rect 11716 17542 11744 19910
rect 11888 19858 11940 19864
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11426 17232 11482 17241
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 11072 16250 11100 16458
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10704 15830 10824 15858
rect 10704 15026 10732 15830
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 14074 10272 14350
rect 10796 14278 10824 15030
rect 10888 14482 10916 16050
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10874 14376 10930 14385
rect 10874 14311 10876 14320
rect 10928 14311 10930 14320
rect 10876 14282 10928 14288
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9876 12102 9904 12718
rect 9968 12646 9996 13631
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12481 9996 12582
rect 9954 12472 10010 12481
rect 9954 12407 10010 12416
rect 9864 12096 9916 12102
rect 9770 12064 9826 12073
rect 9864 12038 9916 12044
rect 9770 11999 9826 12008
rect 9678 11928 9734 11937
rect 9678 11863 9680 11872
rect 9732 11863 9734 11872
rect 9680 11834 9732 11840
rect 9968 11354 9996 12407
rect 10060 12306 10088 12718
rect 10152 12442 10180 13330
rect 10244 12753 10272 14010
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10428 13172 10456 13738
rect 10520 13326 10548 14214
rect 10980 13954 11008 15506
rect 11164 15502 11192 17206
rect 11426 17167 11428 17176
rect 11480 17167 11482 17176
rect 11428 17138 11480 17144
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11426 16552 11482 16561
rect 11426 16487 11428 16496
rect 11480 16487 11482 16496
rect 11520 16516 11572 16522
rect 11428 16458 11480 16464
rect 11520 16458 11572 16464
rect 11532 16425 11560 16458
rect 11518 16416 11574 16425
rect 11518 16351 11574 16360
rect 11242 16144 11298 16153
rect 11242 16079 11244 16088
rect 11296 16079 11298 16088
rect 11244 16050 11296 16056
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11150 15192 11206 15201
rect 11150 15127 11206 15136
rect 11164 14346 11192 15127
rect 11716 14890 11744 17478
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11808 14822 11836 19654
rect 11992 18902 12020 19994
rect 12084 19825 12112 21286
rect 12070 19816 12126 19825
rect 12070 19751 12126 19760
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11900 18057 11928 18770
rect 11980 18352 12032 18358
rect 11978 18320 11980 18329
rect 12032 18320 12034 18329
rect 12084 18290 12112 19654
rect 11978 18255 12034 18264
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11978 18184 12034 18193
rect 11978 18119 12034 18128
rect 11886 18048 11942 18057
rect 11886 17983 11942 17992
rect 11992 17746 12020 18119
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12084 17338 12112 18226
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12176 17218 12204 21898
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 18834 12296 21286
rect 12360 19922 12388 22714
rect 12452 21554 12480 23054
rect 12544 22642 12572 23530
rect 12636 23118 12664 24142
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12440 20936 12492 20942
rect 12438 20904 12440 20913
rect 12492 20904 12494 20913
rect 12438 20839 12494 20848
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12452 19334 12480 20334
rect 12544 20058 12572 22374
rect 12728 21690 12756 25842
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12820 24682 12848 25638
rect 12912 24886 12940 26959
rect 13176 26930 13228 26936
rect 13280 26450 13308 27882
rect 13636 26852 13688 26858
rect 13636 26794 13688 26800
rect 13648 26518 13676 26794
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12820 23322 12848 24618
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12912 23730 12940 24550
rect 13004 23730 13032 26250
rect 13648 26246 13676 26454
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 23588 12952 23594
rect 12900 23530 12952 23536
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12912 23254 12940 23530
rect 12900 23248 12952 23254
rect 12900 23190 12952 23196
rect 13004 22030 13032 23666
rect 13096 22234 13124 25434
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13188 24993 13216 25094
rect 13174 24984 13230 24993
rect 13174 24919 13230 24928
rect 13358 24440 13414 24449
rect 13358 24375 13414 24384
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13280 23905 13308 24074
rect 13266 23896 13322 23905
rect 13266 23831 13322 23840
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12820 21570 12848 21898
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12728 21542 12848 21570
rect 12636 21078 12664 21490
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12728 20913 12756 21542
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12714 20904 12770 20913
rect 12714 20839 12770 20848
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12624 19984 12676 19990
rect 12544 19932 12624 19938
rect 12544 19926 12676 19932
rect 12544 19910 12664 19926
rect 12544 19854 12572 19910
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12360 19310 12480 19334
rect 12348 19306 12480 19310
rect 12348 19304 12400 19306
rect 12348 19246 12400 19252
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12360 18698 12388 19246
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18358 12388 18634
rect 12438 18456 12494 18465
rect 12438 18391 12494 18400
rect 12452 18358 12480 18391
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12268 17678 12296 18294
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12360 17610 12388 18294
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12084 17190 12204 17218
rect 11978 17096 12034 17105
rect 11978 17031 12034 17040
rect 11992 16726 12020 17031
rect 12084 16998 12112 17190
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12176 16522 12204 16662
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11886 15600 11942 15609
rect 11886 15535 11888 15544
rect 11940 15535 11942 15544
rect 11888 15506 11940 15512
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11808 14550 11836 14758
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 10796 13938 11008 13954
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10796 13932 11020 13938
rect 10796 13926 10968 13932
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10322 13152 10378 13161
rect 10428 13144 10548 13172
rect 10322 13087 10378 13096
rect 10336 12986 10364 13087
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10230 12744 10286 12753
rect 10230 12679 10286 12688
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10244 12238 10272 12582
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10138 11928 10194 11937
rect 10138 11863 10194 11872
rect 10152 11694 10180 11863
rect 10140 11688 10192 11694
rect 10232 11688 10284 11694
rect 10140 11630 10192 11636
rect 10230 11656 10232 11665
rect 10284 11656 10286 11665
rect 10230 11591 10286 11600
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10138 11248 10194 11257
rect 10138 11183 10194 11192
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10674 9720 10950
rect 9862 10840 9918 10849
rect 9862 10775 9918 10784
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9876 10198 9904 10775
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 10060 10470 10088 10639
rect 10048 10464 10100 10470
rect 9968 10424 10048 10452
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9586 9752 9642 9761
rect 9586 9687 9588 9696
rect 9640 9687 9642 9696
rect 9588 9658 9640 9664
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9600 8906 9628 9318
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8673 9628 8842
rect 9586 8664 9642 8673
rect 9586 8599 9642 8608
rect 9588 8424 9640 8430
rect 9586 8392 9588 8401
rect 9640 8392 9642 8401
rect 9586 8327 9642 8336
rect 9600 8090 9628 8327
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9402 6080 9458 6089
rect 9402 6015 9458 6024
rect 9600 5302 9628 7686
rect 9692 7478 9720 9318
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9784 6866 9812 9114
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9770 6760 9826 6769
rect 9770 6695 9826 6704
rect 9784 6662 9812 6695
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6390 9812 6598
rect 9772 6384 9824 6390
rect 9692 6344 9772 6372
rect 9692 5574 9720 6344
rect 9772 6326 9824 6332
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9784 5642 9812 5850
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9692 5250 9720 5510
rect 9876 5370 9904 9998
rect 9968 9654 9996 10424
rect 10048 10406 10100 10412
rect 10046 10296 10102 10305
rect 10046 10231 10048 10240
rect 10100 10231 10102 10240
rect 10048 10202 10100 10208
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9692 5234 9904 5250
rect 9692 5228 9916 5234
rect 9692 5222 9864 5228
rect 9864 5170 9916 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9140 2106 9168 5034
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9232 2378 9260 4014
rect 9324 3466 9352 4082
rect 9508 3534 9536 4490
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9600 3126 9628 4082
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3126 9720 3878
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 2922 9812 5102
rect 9968 4010 9996 6938
rect 10060 6390 10088 9862
rect 10152 9654 10180 11183
rect 10244 11150 10272 11494
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10336 10588 10364 12310
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11762 10456 12106
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 11393 10456 11698
rect 10414 11384 10470 11393
rect 10414 11319 10416 11328
rect 10468 11319 10470 11328
rect 10416 11290 10468 11296
rect 10244 10560 10364 10588
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 9178 10180 9590
rect 10244 9450 10272 10560
rect 10520 10266 10548 13144
rect 10704 12832 10732 13874
rect 10796 12986 10824 13926
rect 10968 13874 11020 13880
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10612 12804 10732 12832
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9772 2916 9824 2922
rect 9692 2876 9772 2904
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9508 2038 9536 2790
rect 9692 2530 9720 2876
rect 9772 2858 9824 2864
rect 9956 2644 10008 2650
rect 10060 2632 10088 5850
rect 10244 5846 10272 9386
rect 10336 6730 10364 9930
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10428 8838 10456 9590
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8090 10456 8434
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10520 7274 10548 9046
rect 10612 8974 10640 12804
rect 10782 12472 10838 12481
rect 10782 12407 10838 12416
rect 10796 12306 10824 12407
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10888 12238 10916 13806
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 13394 11008 13670
rect 11058 13560 11114 13569
rect 11164 13530 11192 13874
rect 11058 13495 11114 13504
rect 11152 13524 11204 13530
rect 10968 13388 11020 13394
rect 11072 13376 11100 13495
rect 11152 13466 11204 13472
rect 11152 13388 11204 13394
rect 11072 13348 11152 13376
rect 10968 13330 11020 13336
rect 11152 13330 11204 13336
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12986 11192 13126
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10704 9110 10732 12174
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10796 9518 10824 12106
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11354 10916 12038
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10888 10538 10916 10678
rect 10980 10674 11008 12922
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12374 11100 12582
rect 11164 12442 11192 12786
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11256 12186 11284 14418
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11348 14113 11376 14282
rect 11334 14104 11390 14113
rect 11334 14039 11390 14048
rect 11532 13802 11560 14418
rect 11900 14226 11928 15506
rect 11992 14550 12020 16186
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12084 14657 12112 15846
rect 12070 14648 12126 14657
rect 12070 14583 12126 14592
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11716 14198 11928 14226
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11716 13870 11744 14198
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11348 13258 11376 13466
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12782 11468 13126
rect 11612 12980 11664 12986
rect 11716 12968 11744 13806
rect 11808 13705 11836 14010
rect 11794 13696 11850 13705
rect 11794 13631 11850 13640
rect 11808 13258 11836 13631
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11664 12940 11744 12968
rect 11612 12922 11664 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11428 12776 11480 12782
rect 11624 12753 11652 12786
rect 11428 12718 11480 12724
rect 11610 12744 11666 12753
rect 11610 12679 11666 12688
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11164 12158 11284 12186
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 11072 10266 11100 11018
rect 11164 10606 11192 12158
rect 11244 12096 11296 12102
rect 11716 12050 11744 12940
rect 11244 12038 11296 12044
rect 11256 11830 11284 12038
rect 11624 12022 11744 12050
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11624 11762 11652 12022
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 11665 11652 11698
rect 11610 11656 11666 11665
rect 11610 11591 11666 11600
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10784 8900 10836 8906
rect 10888 8888 10916 9862
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10836 8860 10916 8888
rect 10784 8842 10836 8848
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 7886 10640 8774
rect 10784 8424 10836 8430
rect 10782 8392 10784 8401
rect 10836 8392 10838 8401
rect 10782 8327 10838 8336
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10232 5228 10284 5234
rect 10336 5216 10364 6258
rect 10284 5188 10364 5216
rect 10232 5170 10284 5176
rect 10152 4282 10180 5170
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10008 2604 10088 2632
rect 9956 2586 10008 2592
rect 9692 2502 9812 2530
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 9692 1970 9720 2382
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 9680 1964 9732 1970
rect 9680 1906 9732 1912
rect 9784 1494 9812 2502
rect 10152 2446 10180 3470
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9772 1488 9824 1494
rect 9772 1430 9824 1436
rect 10336 1358 10364 3402
rect 10428 3398 10456 7142
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10520 4010 10548 6938
rect 10704 6882 10732 8026
rect 10612 6854 10732 6882
rect 10612 5642 10640 6854
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10612 4826 10640 5578
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10520 2774 10548 3946
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3058 10640 3878
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10428 2746 10548 2774
rect 10428 2632 10456 2746
rect 10508 2644 10560 2650
rect 10428 2604 10508 2632
rect 10508 2586 10560 2592
rect 10704 1358 10732 6734
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6254 10824 6666
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5302 10824 6190
rect 10888 6186 10916 8860
rect 10980 8498 11008 9522
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 6934 11008 8434
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11072 6746 11100 8570
rect 11164 8294 11192 9930
rect 11256 9625 11284 10950
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11610 10160 11666 10169
rect 11610 10095 11666 10104
rect 11624 10062 11652 10095
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11624 9654 11652 9998
rect 11612 9648 11664 9654
rect 11242 9616 11298 9625
rect 11612 9590 11664 9596
rect 11242 9551 11298 9560
rect 11624 9489 11652 9590
rect 11716 9586 11744 11863
rect 11808 11150 11836 12038
rect 11900 11354 11928 14010
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11992 11218 12020 14214
rect 12084 13734 12112 14583
rect 12176 14113 12204 16458
rect 12268 15094 12296 17070
rect 12360 16590 12388 17546
rect 12452 16590 12480 18294
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12544 17338 12572 17682
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12532 16108 12584 16114
rect 12636 16096 12664 19790
rect 12728 17626 12756 20839
rect 12820 18630 12848 21014
rect 12912 19990 12940 21626
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13004 21146 13032 21490
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13096 21026 13124 21082
rect 13004 20998 13124 21026
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12912 19417 12940 19926
rect 13004 19718 13032 20998
rect 13188 20874 13216 22986
rect 13280 22098 13308 23666
rect 13372 22710 13400 24375
rect 13464 23866 13492 25842
rect 13740 25344 13768 28358
rect 13832 27674 13860 30874
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13924 27470 13952 32166
rect 14016 28694 14044 33594
rect 19156 33584 19208 33590
rect 19156 33526 19208 33532
rect 16764 33516 16816 33522
rect 16764 33458 16816 33464
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 14464 33448 14516 33454
rect 14464 33390 14516 33396
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 14108 31890 14136 33050
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14384 32434 14412 32506
rect 14476 32434 14504 33390
rect 16488 33380 16540 33386
rect 16488 33322 16540 33328
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14660 32434 14688 32710
rect 14842 32668 15150 32677
rect 14842 32666 14848 32668
rect 14904 32666 14928 32668
rect 14984 32666 15008 32668
rect 15064 32666 15088 32668
rect 15144 32666 15150 32668
rect 14904 32614 14906 32666
rect 15086 32614 15088 32666
rect 14842 32612 14848 32614
rect 14904 32612 14928 32614
rect 14984 32612 15008 32614
rect 15064 32612 15088 32614
rect 15144 32612 15150 32614
rect 14842 32603 15150 32612
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 14188 32360 14240 32366
rect 14556 32360 14608 32366
rect 14240 32308 14320 32314
rect 14188 32302 14320 32308
rect 14556 32302 14608 32308
rect 14200 32286 14320 32302
rect 14096 31884 14148 31890
rect 14096 31826 14148 31832
rect 14292 31754 14320 32286
rect 14188 31748 14240 31754
rect 14292 31726 14412 31754
rect 14188 31690 14240 31696
rect 14200 30546 14228 31690
rect 14200 30518 14320 30546
rect 14188 30388 14240 30394
rect 14188 30330 14240 30336
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14108 29345 14136 29650
rect 14094 29336 14150 29345
rect 14094 29271 14150 29280
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14004 28688 14056 28694
rect 14004 28630 14056 28636
rect 14108 28626 14136 29174
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14200 28218 14228 30330
rect 14292 29646 14320 30518
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14384 29306 14412 31726
rect 14568 31278 14596 32302
rect 14844 32298 15332 32314
rect 14832 32292 15332 32298
rect 14884 32286 15332 32292
rect 14832 32234 14884 32240
rect 15304 31754 15332 32286
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 15304 31726 15516 31754
rect 15292 31680 15344 31686
rect 15290 31648 15292 31657
rect 15344 31648 15346 31657
rect 14842 31580 15150 31589
rect 15290 31583 15346 31592
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 14740 31408 14792 31414
rect 14740 31350 14792 31356
rect 14556 31272 14608 31278
rect 14556 31214 14608 31220
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14476 30394 14504 31078
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14476 29102 14504 30126
rect 14568 29782 14596 31214
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14660 30433 14688 30534
rect 14646 30424 14702 30433
rect 14646 30359 14702 30368
rect 14752 30190 14780 31350
rect 15488 31346 15516 31726
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15200 31136 15252 31142
rect 15200 31078 15252 31084
rect 15474 31104 15530 31113
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 14832 30388 14884 30394
rect 14832 30330 14884 30336
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 14556 29776 14608 29782
rect 14556 29718 14608 29724
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14280 28960 14332 28966
rect 14280 28902 14332 28908
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 14108 27130 14136 28018
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14108 26994 14136 27066
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14002 26616 14058 26625
rect 14002 26551 14004 26560
rect 14056 26551 14058 26560
rect 14004 26522 14056 26528
rect 13910 25528 13966 25537
rect 13910 25463 13966 25472
rect 13820 25424 13872 25430
rect 13820 25366 13872 25372
rect 13648 25316 13768 25344
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13556 23798 13584 24754
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13372 21978 13400 22510
rect 13280 21950 13400 21978
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13280 20754 13308 21950
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 20942 13400 21830
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13280 20726 13400 20754
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13084 20392 13136 20398
rect 13082 20360 13084 20369
rect 13136 20360 13138 20369
rect 13082 20295 13138 20304
rect 13082 20224 13138 20233
rect 13082 20159 13138 20168
rect 13096 20058 13124 20159
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12898 19408 12954 19417
rect 12898 19343 12954 19352
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12806 18320 12862 18329
rect 12806 18255 12862 18264
rect 12820 17882 12848 18255
rect 12912 18222 12940 19178
rect 13004 18698 13032 19654
rect 13188 19446 13216 19790
rect 13280 19446 13308 20402
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 13266 19272 13322 19281
rect 13266 19207 13322 19216
rect 13280 19174 13308 19207
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12728 17598 12940 17626
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12728 16590 12756 16730
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 16114 12756 16186
rect 12584 16068 12664 16096
rect 12716 16108 12768 16114
rect 12532 16050 12584 16056
rect 12716 16050 12768 16056
rect 12820 16046 12848 17478
rect 12912 16998 12940 17598
rect 13004 17134 13032 18634
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12900 16992 12952 16998
rect 13096 16980 13124 18566
rect 13372 18358 13400 20726
rect 13464 20534 13492 22918
rect 13556 22030 13584 22918
rect 13648 22794 13676 25316
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13740 24138 13768 25162
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13832 23866 13860 25366
rect 13924 24206 13952 25463
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 14016 23186 14044 25230
rect 14108 25158 14136 26930
rect 14200 26761 14228 26930
rect 14186 26752 14242 26761
rect 14186 26687 14242 26696
rect 14292 25752 14320 28902
rect 14384 28150 14412 28902
rect 14568 28234 14596 29582
rect 14844 29560 14872 30330
rect 15014 30016 15070 30025
rect 15014 29951 15070 29960
rect 14924 29776 14976 29782
rect 15028 29764 15056 29951
rect 14976 29736 15056 29764
rect 14924 29718 14976 29724
rect 15028 29646 15056 29736
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14752 29532 14872 29560
rect 14646 29472 14702 29481
rect 14646 29407 14702 29416
rect 14660 29073 14688 29407
rect 14646 29064 14702 29073
rect 14646 28999 14702 29008
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14476 28206 14596 28234
rect 14372 28144 14424 28150
rect 14372 28086 14424 28092
rect 14476 28082 14504 28206
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14384 27713 14412 27950
rect 14370 27704 14426 27713
rect 14370 27639 14372 27648
rect 14424 27639 14426 27648
rect 14372 27610 14424 27616
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14200 25724 14320 25752
rect 14200 25294 14228 25724
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14188 25152 14240 25158
rect 14188 25094 14240 25100
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 13648 22778 13768 22794
rect 14108 22778 14136 24006
rect 13648 22772 13780 22778
rect 13648 22766 13728 22772
rect 13728 22714 13780 22720
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14200 22710 14228 25094
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14292 23633 14320 24006
rect 14278 23624 14334 23633
rect 14278 23559 14334 23568
rect 14384 23254 14412 27406
rect 14556 27396 14608 27402
rect 14556 27338 14608 27344
rect 14568 27130 14596 27338
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14476 25922 14504 26454
rect 14660 26450 14688 28630
rect 14752 27849 14780 29532
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 15212 29238 15240 31078
rect 15474 31039 15530 31048
rect 15384 30796 15436 30802
rect 15384 30738 15436 30744
rect 15292 30592 15344 30598
rect 15290 30560 15292 30569
rect 15344 30560 15346 30569
rect 15290 30495 15346 30504
rect 15396 30326 15424 30738
rect 15488 30598 15516 31039
rect 15580 30734 15608 31622
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15384 30320 15436 30326
rect 15384 30262 15436 30268
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 14832 29232 14884 29238
rect 14832 29174 14884 29180
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 14844 29034 14872 29174
rect 14832 29028 14884 29034
rect 14832 28970 14884 28976
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 14844 28422 14872 28970
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 15212 28082 15240 28970
rect 15108 28076 15160 28082
rect 15108 28018 15160 28024
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15120 27946 15148 28018
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 14738 27840 14794 27849
rect 14738 27775 14794 27784
rect 15304 27606 15332 30194
rect 15488 30190 15516 30534
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15580 30138 15608 30670
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15672 30240 15700 30534
rect 15764 30394 15792 31758
rect 15936 30660 15988 30666
rect 15936 30602 15988 30608
rect 15948 30433 15976 30602
rect 15934 30424 15990 30433
rect 15752 30388 15804 30394
rect 15934 30359 15990 30368
rect 15752 30330 15804 30336
rect 15936 30320 15988 30326
rect 15936 30262 15988 30268
rect 15672 30212 15792 30240
rect 15580 30110 15700 30138
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15382 29336 15438 29345
rect 15382 29271 15384 29280
rect 15436 29271 15438 29280
rect 15384 29242 15436 29248
rect 15384 29164 15436 29170
rect 15384 29106 15436 29112
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14648 26240 14700 26246
rect 14646 26208 14648 26217
rect 14700 26208 14702 26217
rect 14646 26143 14702 26152
rect 14476 25894 14688 25922
rect 14554 25800 14610 25809
rect 14554 25735 14610 25744
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 24138 14504 25638
rect 14568 25265 14596 25735
rect 14554 25256 14610 25265
rect 14554 25191 14610 25200
rect 14554 25120 14610 25129
rect 14554 25055 14610 25064
rect 14568 24682 14596 25055
rect 14660 24936 14688 25894
rect 14752 25809 14780 26998
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15120 26790 15148 26930
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 14830 26616 14886 26625
rect 14830 26551 14886 26560
rect 14844 26382 14872 26551
rect 15120 26518 15148 26726
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14738 25800 14794 25809
rect 14738 25735 14794 25744
rect 15014 25528 15070 25537
rect 15014 25463 15016 25472
rect 15068 25463 15070 25472
rect 15016 25434 15068 25440
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14660 24908 14872 24936
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 14844 24206 14872 24908
rect 15014 24440 15070 24449
rect 15014 24375 15070 24384
rect 15028 24206 15056 24375
rect 15212 24342 15240 27338
rect 15290 27296 15346 27305
rect 15290 27231 15346 27240
rect 15304 26625 15332 27231
rect 15396 27130 15424 29106
rect 15488 29102 15516 29446
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15488 27470 15516 27950
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15474 27160 15530 27169
rect 15384 27124 15436 27130
rect 15474 27095 15530 27104
rect 15384 27066 15436 27072
rect 15488 27062 15516 27095
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15290 26616 15346 26625
rect 15290 26551 15346 26560
rect 15292 26240 15344 26246
rect 15290 26208 15292 26217
rect 15344 26208 15346 26217
rect 15290 26143 15346 26152
rect 15396 25294 15424 26930
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15304 24886 15332 25162
rect 15292 24880 15344 24886
rect 15292 24822 15344 24828
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14464 23656 14516 23662
rect 14462 23624 14464 23633
rect 14516 23624 14518 23633
rect 14462 23559 14518 23568
rect 14568 23322 14596 24142
rect 14752 23866 14780 24142
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15200 23792 15252 23798
rect 15304 23780 15332 24822
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15252 23752 15332 23780
rect 15200 23734 15252 23740
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 13636 22704 13688 22710
rect 14188 22704 14240 22710
rect 13636 22646 13688 22652
rect 13910 22672 13966 22681
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13556 20602 13584 21966
rect 13648 21146 13676 22646
rect 14188 22646 14240 22652
rect 13910 22607 13966 22616
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13726 22128 13782 22137
rect 13726 22063 13782 22072
rect 13740 21706 13768 22063
rect 13832 21894 13860 22510
rect 13924 22438 13952 22607
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13740 21678 13860 21706
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13634 20496 13690 20505
rect 13634 20431 13690 20440
rect 13648 20058 13676 20431
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13452 19848 13504 19854
rect 13504 19808 13584 19836
rect 13452 19790 13504 19796
rect 13556 19446 13584 19808
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13280 17678 13308 18226
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13268 17672 13320 17678
rect 13266 17640 13268 17649
rect 13320 17640 13322 17649
rect 13266 17575 13322 17584
rect 13372 17270 13400 18158
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 12900 16934 12952 16940
rect 13004 16952 13124 16980
rect 13004 16726 13032 16952
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12440 15904 12492 15910
rect 12492 15864 12572 15892
rect 12440 15846 12492 15852
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12256 15088 12308 15094
rect 12308 15048 12388 15076
rect 12256 15030 12308 15036
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 14550 12296 14758
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12256 14408 12308 14414
rect 12254 14376 12256 14385
rect 12308 14376 12310 14385
rect 12254 14311 12310 14320
rect 12162 14104 12218 14113
rect 12162 14039 12218 14048
rect 12360 13938 12388 15048
rect 12452 14929 12480 15098
rect 12438 14920 12494 14929
rect 12438 14855 12494 14864
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 12306 12112 13670
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 12764 12204 13398
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12360 13190 12388 13262
rect 12348 13184 12400 13190
rect 12452 13161 12480 13262
rect 12348 13126 12400 13132
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12176 12736 12296 12764
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11898 12112 12106
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12070 11520 12126 11529
rect 12070 11455 12126 11464
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11610 9480 11666 9489
rect 11610 9415 11666 9424
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11612 9172 11664 9178
rect 11664 9132 11744 9160
rect 11612 9114 11664 9120
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 8809 11376 8842
rect 11334 8800 11390 8809
rect 11334 8735 11390 8744
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10980 6718 11100 6746
rect 10980 6202 11008 6718
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6322 11100 6598
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10876 6180 10928 6186
rect 10980 6174 11100 6202
rect 10876 6122 10928 6128
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10888 5710 10916 5782
rect 11072 5710 11100 6174
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11164 5352 11192 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 6882 11284 7686
rect 11716 7290 11744 9132
rect 11808 8566 11836 10406
rect 11900 9178 11928 11086
rect 11978 10296 12034 10305
rect 11978 10231 11980 10240
rect 12032 10231 12034 10240
rect 11980 10202 12032 10208
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11992 9897 12020 9998
rect 11978 9888 12034 9897
rect 11978 9823 12034 9832
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11992 8022 12020 9522
rect 12084 9466 12112 11455
rect 12176 10169 12204 12582
rect 12268 11937 12296 12736
rect 12348 12368 12400 12374
rect 12544 12345 12572 15864
rect 12636 15026 12664 15914
rect 12820 15434 12848 15982
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12728 14618 12756 15302
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 14006 12756 14554
rect 12912 14482 12940 16050
rect 13004 15162 13032 16390
rect 13096 15609 13124 16526
rect 13188 16114 13216 17206
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13280 16969 13308 17070
rect 13266 16960 13322 16969
rect 13266 16895 13322 16904
rect 13280 16182 13308 16895
rect 13372 16522 13400 17206
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13280 15978 13308 16118
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13082 15600 13138 15609
rect 13082 15535 13138 15544
rect 13372 15502 13400 16458
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13096 15162 13124 15438
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13096 14498 13124 15098
rect 13360 15020 13412 15026
rect 13464 15008 13492 19110
rect 13556 18290 13584 19382
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18426 13676 18566
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13556 17270 13584 18022
rect 13648 17882 13676 18022
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13740 17338 13768 21286
rect 13832 18970 13860 21678
rect 13924 21010 13952 22374
rect 14094 21448 14150 21457
rect 14094 21383 14150 21392
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 19446 13952 20742
rect 14016 20398 14044 20810
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 14016 19446 14044 20198
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14016 18766 14044 19382
rect 14108 19174 14136 21383
rect 14200 20262 14228 22646
rect 14292 21622 14320 22986
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14476 20602 14504 22578
rect 14568 21146 14596 23122
rect 14660 22030 14688 23190
rect 14752 22166 14780 23598
rect 14832 23520 14884 23526
rect 14830 23488 14832 23497
rect 14884 23488 14886 23497
rect 14830 23423 14886 23432
rect 15028 23322 15056 23666
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 15212 22760 15240 23734
rect 15396 23254 15424 24210
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15120 22732 15240 22760
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 15028 22273 15056 22374
rect 15014 22264 15070 22273
rect 15014 22199 15070 22208
rect 15120 22166 15148 22732
rect 14740 22160 14792 22166
rect 14740 22102 14792 22108
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14292 19334 14320 19722
rect 14200 19306 14320 19334
rect 14096 19168 14148 19174
rect 14200 19145 14228 19306
rect 14096 19110 14148 19116
rect 14186 19136 14242 19145
rect 14186 19071 14242 19080
rect 14004 18760 14056 18766
rect 13910 18728 13966 18737
rect 14004 18702 14056 18708
rect 13910 18663 13966 18672
rect 13818 17912 13874 17921
rect 13818 17847 13820 17856
rect 13872 17847 13874 17856
rect 13820 17818 13872 17824
rect 13924 17728 13952 18663
rect 14016 18057 14044 18702
rect 14200 18290 14228 19071
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14002 18048 14058 18057
rect 14002 17983 14058 17992
rect 14002 17912 14058 17921
rect 14002 17847 14058 17856
rect 13832 17700 13952 17728
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13832 17270 13860 17700
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13924 17513 13952 17546
rect 13910 17504 13966 17513
rect 13910 17439 13966 17448
rect 13924 17270 13952 17439
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13556 16454 13584 17206
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13542 16008 13598 16017
rect 13542 15943 13598 15952
rect 13556 15910 13584 15943
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13544 15020 13596 15026
rect 13464 14980 13544 15008
rect 13360 14962 13412 14968
rect 13544 14962 13596 14968
rect 13372 14634 13400 14962
rect 13372 14606 13492 14634
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13004 14470 13124 14498
rect 13358 14512 13414 14521
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12348 12310 12400 12316
rect 12530 12336 12586 12345
rect 12254 11928 12310 11937
rect 12254 11863 12256 11872
rect 12308 11863 12310 11872
rect 12256 11834 12308 11840
rect 12254 11656 12310 11665
rect 12254 11591 12310 11600
rect 12268 10849 12296 11591
rect 12254 10840 12310 10849
rect 12254 10775 12310 10784
rect 12268 10674 12296 10775
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12360 10470 12388 12310
rect 12530 12271 12586 12280
rect 12636 11354 12664 13670
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12256 10056 12308 10062
rect 12360 10044 12388 10406
rect 12452 10130 12480 10950
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12308 10016 12388 10044
rect 12256 9998 12308 10004
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12176 9654 12204 9930
rect 12452 9926 12480 10066
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12084 9438 12296 9466
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12162 9344 12218 9353
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7313 12020 7958
rect 11978 7304 12034 7313
rect 11716 7262 11928 7290
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11256 6854 11376 6882
rect 11244 6792 11296 6798
rect 11242 6760 11244 6769
rect 11296 6760 11298 6769
rect 11242 6695 11298 6704
rect 11348 6202 11376 6854
rect 11072 5324 11192 5352
rect 11256 6174 11376 6202
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10324 1352 10376 1358
rect 8206 1320 8262 1329
rect 10324 1294 10376 1300
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 10888 1290 10916 2790
rect 10980 2514 11008 4966
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 8206 1255 8208 1264
rect 8260 1255 8262 1264
rect 10876 1284 10928 1290
rect 8208 1226 8260 1232
rect 10876 1226 10928 1232
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 9956 1216 10008 1222
rect 9956 1158 10008 1164
rect 4068 876 4120 882
rect 4068 818 4120 824
rect 5920 814 5948 1158
rect 7896 1116 8204 1125
rect 7896 1114 7902 1116
rect 7958 1114 7982 1116
rect 8038 1114 8062 1116
rect 8118 1114 8142 1116
rect 8198 1114 8204 1116
rect 7958 1062 7960 1114
rect 8140 1062 8142 1114
rect 7896 1060 7902 1062
rect 7958 1060 7982 1062
rect 8038 1060 8062 1062
rect 8118 1060 8142 1062
rect 8198 1060 8204 1062
rect 7896 1051 8204 1060
rect 9968 950 9996 1158
rect 10980 1018 11008 1906
rect 11072 1358 11100 5324
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4826 11192 5170
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11164 2106 11192 4626
rect 11256 2990 11284 6174
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11256 2446 11284 2586
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11256 1426 11284 2382
rect 11716 2310 11744 7142
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 4758 11836 6258
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11900 4622 11928 7262
rect 11978 7239 12034 7248
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11369 1660 11677 1669
rect 11369 1658 11375 1660
rect 11431 1658 11455 1660
rect 11511 1658 11535 1660
rect 11591 1658 11615 1660
rect 11671 1658 11677 1660
rect 11431 1606 11433 1658
rect 11613 1606 11615 1658
rect 11369 1604 11375 1606
rect 11431 1604 11455 1606
rect 11511 1604 11535 1606
rect 11591 1604 11615 1606
rect 11671 1604 11677 1606
rect 11369 1595 11677 1604
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11808 1358 11836 4490
rect 12084 3670 12112 9318
rect 12162 9279 12218 9288
rect 12176 7818 12204 9279
rect 12268 8906 12296 9438
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12360 7993 12388 9114
rect 12346 7984 12402 7993
rect 12346 7919 12402 7928
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6905 12204 6938
rect 12162 6896 12218 6905
rect 12162 6831 12218 6840
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12176 6118 12204 6394
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12176 3058 12204 4422
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12268 1834 12296 7346
rect 12452 6769 12480 9862
rect 12544 9178 12572 11222
rect 12728 10130 12756 13767
rect 12912 12918 12940 13874
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12442 12848 12786
rect 12898 12744 12954 12753
rect 12898 12679 12954 12688
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12912 10810 12940 12679
rect 13004 11150 13032 14470
rect 13358 14447 13414 14456
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13096 12102 13124 14350
rect 13280 13734 13308 14350
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13372 13530 13400 14447
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13464 13326 13492 14606
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13556 13841 13584 14010
rect 13542 13832 13598 13841
rect 13542 13767 13598 13776
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13542 13288 13598 13297
rect 13542 13223 13598 13232
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13372 11354 13400 13126
rect 13464 12170 13492 13126
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 11014 13032 11086
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12636 8974 12664 9318
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12452 6474 12480 6695
rect 12360 6446 12480 6474
rect 12360 6322 12388 6446
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12452 6202 12480 6326
rect 12360 6174 12480 6202
rect 12360 4554 12388 6174
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12544 4214 12572 7919
rect 12636 5370 12664 8230
rect 12728 7002 12756 9930
rect 12820 9654 12848 10746
rect 13082 10704 13138 10713
rect 13082 10639 13138 10648
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12820 7818 12848 9590
rect 12898 9480 12954 9489
rect 12898 9415 12954 9424
rect 12912 9382 12940 9415
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 13004 9178 13032 10202
rect 13096 9466 13124 10639
rect 13174 10568 13230 10577
rect 13174 10503 13230 10512
rect 13188 10266 13216 10503
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13174 10024 13230 10033
rect 13174 9959 13230 9968
rect 13188 9654 13216 9959
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13096 9438 13216 9466
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12898 8800 12954 8809
rect 12898 8735 12954 8744
rect 12912 8294 12940 8735
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12820 7546 12848 7754
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7478 12940 8230
rect 13096 7886 13124 9318
rect 13188 8838 13216 9438
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8362 13216 8774
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12912 6934 12940 7414
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 4622 12756 6122
rect 12912 5914 12940 6734
rect 13004 5914 13032 6734
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 13004 5545 13032 5578
rect 12990 5536 13046 5545
rect 12990 5471 13046 5480
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12348 4072 12400 4078
rect 12728 4060 12756 4558
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12400 4032 12756 4060
rect 12348 4014 12400 4020
rect 12360 2038 12388 4014
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12544 2038 12572 2858
rect 12636 2582 12664 2926
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12348 2032 12400 2038
rect 12348 1974 12400 1980
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 12728 1834 12756 3130
rect 12820 2650 12848 3606
rect 12912 3534 12940 4422
rect 13096 3670 13124 7142
rect 13280 6798 13308 11290
rect 13556 11218 13584 13223
rect 13648 12782 13676 16934
rect 13832 16454 13860 17002
rect 13924 16674 13952 17206
rect 14016 16794 14044 17847
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13924 16646 14044 16674
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13740 14618 13768 16390
rect 13910 15464 13966 15473
rect 13910 15399 13966 15408
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13832 14618 13860 15030
rect 13924 14890 13952 15399
rect 14016 15201 14044 16646
rect 14002 15192 14058 15201
rect 14002 15127 14058 15136
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13726 13968 13782 13977
rect 13726 13903 13728 13912
rect 13780 13903 13782 13912
rect 13728 13874 13780 13880
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13740 11801 13768 13670
rect 13832 13462 13860 14010
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13832 12850 13860 12922
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13924 12434 13952 14486
rect 14016 13258 14044 14962
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14016 12986 14044 13194
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13832 12406 13952 12434
rect 13726 11792 13782 11801
rect 13636 11756 13688 11762
rect 13726 11727 13782 11736
rect 13636 11698 13688 11704
rect 13648 11626 13676 11698
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13648 11150 13676 11562
rect 13636 11144 13688 11150
rect 13450 11112 13506 11121
rect 13636 11086 13688 11092
rect 13450 11047 13506 11056
rect 13728 11076 13780 11082
rect 13464 10062 13492 11047
rect 13728 11018 13780 11024
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13372 6458 13400 9522
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13464 9178 13492 9386
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13450 8664 13506 8673
rect 13450 8599 13506 8608
rect 13464 8498 13492 8599
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13450 8392 13506 8401
rect 13450 8327 13506 8336
rect 13464 7002 13492 8327
rect 13556 8294 13584 10678
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10130 13676 10610
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 8974 13676 9862
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13740 8838 13768 11018
rect 13832 9178 13860 12406
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13924 11558 13952 12135
rect 14108 11830 14136 18158
rect 14200 16794 14228 18226
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14292 15858 14320 18634
rect 14384 16998 14412 19790
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 19514 14504 19654
rect 14660 19553 14688 21830
rect 14752 20584 14780 22102
rect 15120 21894 15148 22102
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15212 21672 15240 21830
rect 15120 21644 15240 21672
rect 15120 20874 15148 21644
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14752 20556 14964 20584
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14844 20210 14872 20402
rect 14752 20182 14872 20210
rect 14646 19544 14702 19553
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14556 19508 14608 19514
rect 14646 19479 14702 19488
rect 14556 19450 14608 19456
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14476 16182 14504 18634
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14292 15830 14504 15858
rect 14476 15638 14504 15830
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14200 14906 14228 15506
rect 14200 14878 14320 14906
rect 14292 14822 14320 14878
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14278 14648 14334 14657
rect 14278 14583 14334 14592
rect 14292 14482 14320 14583
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13938 14228 14214
rect 14384 14090 14412 15506
rect 14568 14890 14596 19450
rect 14660 19446 14688 19479
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14752 19394 14780 20182
rect 14936 19854 14964 20556
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 15106 19816 15162 19825
rect 14936 19718 14964 19790
rect 15106 19751 15162 19760
rect 15120 19718 15148 19751
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14832 19440 14884 19446
rect 14752 19388 14832 19394
rect 14752 19382 14884 19388
rect 14922 19408 14978 19417
rect 14752 19366 14872 19382
rect 14922 19343 14978 19352
rect 14936 19174 14964 19343
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15212 18698 15240 21286
rect 15304 21146 15332 22918
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15304 18986 15332 20334
rect 15396 19854 15424 22714
rect 15488 20058 15516 26182
rect 15580 24698 15608 29990
rect 15672 28558 15700 30110
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15764 28218 15792 30212
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15856 28529 15884 30058
rect 15948 30054 15976 30262
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 15948 28966 15976 29514
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15842 28520 15898 28529
rect 15842 28455 15898 28464
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15660 27872 15712 27878
rect 15660 27814 15712 27820
rect 15672 24818 15700 27814
rect 15764 27538 15792 28154
rect 15948 27962 15976 28902
rect 16040 28762 16068 32370
rect 16212 32292 16264 32298
rect 16212 32234 16264 32240
rect 16120 30048 16172 30054
rect 16118 30016 16120 30025
rect 16172 30016 16174 30025
rect 16118 29951 16174 29960
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 15948 27946 16068 27962
rect 15948 27940 16080 27946
rect 15948 27934 16028 27940
rect 16028 27882 16080 27888
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15764 27334 15792 27474
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15844 27056 15896 27062
rect 15764 27016 15844 27044
rect 15764 24818 15792 27016
rect 15844 26998 15896 27004
rect 16132 26518 16160 29514
rect 16224 29345 16252 32234
rect 16304 31748 16356 31754
rect 16304 31690 16356 31696
rect 16316 31521 16344 31690
rect 16302 31512 16358 31521
rect 16302 31447 16358 31456
rect 16302 30016 16358 30025
rect 16302 29951 16358 29960
rect 16210 29336 16266 29345
rect 16210 29271 16266 29280
rect 16224 29034 16252 29271
rect 16212 29028 16264 29034
rect 16212 28970 16264 28976
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16224 28014 16252 28154
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16316 26858 16344 29951
rect 16408 29646 16436 32914
rect 16500 32774 16528 33322
rect 16776 32978 16804 33458
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 16764 32972 16816 32978
rect 16764 32914 16816 32920
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16868 32552 16896 33322
rect 17144 33182 17172 33458
rect 17316 33244 17368 33250
rect 17316 33186 17368 33192
rect 17132 33176 17184 33182
rect 17132 33118 17184 33124
rect 16960 32966 17264 32994
rect 16960 32910 16988 32966
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 16868 32524 16988 32552
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16580 31748 16632 31754
rect 16684 31736 16712 32302
rect 16632 31708 16712 31736
rect 16580 31690 16632 31696
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 16500 30870 16528 31418
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16488 30864 16540 30870
rect 16488 30806 16540 30812
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16500 29306 16528 29786
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 16500 26382 16528 27882
rect 16592 27130 16620 31282
rect 16684 31210 16712 31708
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16672 31204 16724 31210
rect 16672 31146 16724 31152
rect 16670 29880 16726 29889
rect 16670 29815 16726 29824
rect 16684 29306 16712 29815
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16776 29238 16804 29718
rect 16764 29232 16816 29238
rect 16764 29174 16816 29180
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24993 15884 25230
rect 15842 24984 15898 24993
rect 15842 24919 15898 24928
rect 15948 24818 15976 26250
rect 16040 25430 16068 26250
rect 16132 25430 16160 26318
rect 16500 25906 16528 26318
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16488 25900 16540 25906
rect 16488 25842 16540 25848
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 16120 25424 16172 25430
rect 16120 25366 16172 25372
rect 16132 24818 16160 25366
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16040 24721 16068 24754
rect 16026 24712 16082 24721
rect 15580 24670 15700 24698
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 20262 15608 24550
rect 15672 23526 15700 24670
rect 16026 24647 16082 24656
rect 16224 24206 16252 25842
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16316 25129 16344 25638
rect 16488 25152 16540 25158
rect 16302 25120 16358 25129
rect 16488 25094 16540 25100
rect 16302 25055 16358 25064
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15948 23633 15976 23666
rect 15934 23624 15990 23633
rect 15934 23559 15990 23568
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15764 23050 15792 23258
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15672 22438 15700 22578
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15764 21962 15792 22986
rect 15948 22094 15976 23559
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 16040 22817 16068 23258
rect 16026 22808 16082 22817
rect 16026 22743 16082 22752
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16040 22098 16068 22578
rect 15856 22066 15976 22094
rect 16028 22092 16080 22098
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15764 21622 15792 21898
rect 15856 21690 15884 22066
rect 16028 22034 16080 22040
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15672 19786 15700 21082
rect 15764 20942 15792 21558
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15764 20398 15792 20878
rect 16040 20874 16068 21830
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19961 15792 20198
rect 15948 20074 15976 20810
rect 16028 20256 16080 20262
rect 16026 20224 16028 20233
rect 16080 20224 16082 20233
rect 16026 20159 16082 20168
rect 15948 20046 16068 20074
rect 15750 19952 15806 19961
rect 15750 19887 15806 19896
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15304 18958 15424 18986
rect 15396 18766 15424 18958
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15292 18624 15344 18630
rect 15212 18572 15292 18578
rect 15212 18566 15344 18572
rect 15212 18550 15332 18566
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14646 18320 14702 18329
rect 14646 18255 14702 18264
rect 14660 17134 14688 18255
rect 14844 18086 14872 18362
rect 15014 18184 15070 18193
rect 15014 18119 15016 18128
rect 15068 18119 15070 18128
rect 15016 18090 15068 18096
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 15212 17746 15240 18550
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15290 18048 15346 18057
rect 15290 17983 15346 17992
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15016 17672 15068 17678
rect 15068 17620 15240 17626
rect 15016 17614 15240 17620
rect 15028 17598 15240 17614
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14660 16250 14688 17070
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14660 14482 14688 15846
rect 14752 15162 14780 16934
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14936 15706 14964 16186
rect 15212 16114 15240 17598
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14646 14376 14702 14385
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14292 14062 14412 14090
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14200 13433 14228 13738
rect 14186 13424 14242 13433
rect 14186 13359 14242 13368
rect 14292 12850 14320 14062
rect 14370 13968 14426 13977
rect 14370 13903 14426 13912
rect 14384 13394 14412 13903
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14476 13274 14504 14214
rect 14568 13433 14596 14350
rect 14646 14311 14702 14320
rect 14554 13424 14610 13433
rect 14554 13359 14610 13368
rect 14476 13246 14596 13274
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14200 11830 14228 12310
rect 14384 12238 14412 12854
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13924 10674 13952 11290
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14016 9704 14044 11698
rect 14292 11336 14320 12174
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14200 11308 14320 11336
rect 14016 9676 14136 9704
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13648 8090 13676 8434
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 6202 13400 6394
rect 13464 6322 13492 6938
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13372 6174 13492 6202
rect 13174 6080 13230 6089
rect 13174 6015 13230 6024
rect 13188 5778 13216 6015
rect 13358 5944 13414 5953
rect 13358 5879 13414 5888
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13268 5636 13320 5642
rect 13372 5624 13400 5879
rect 13320 5596 13400 5624
rect 13268 5578 13320 5584
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13188 3534 13216 5578
rect 13372 5234 13400 5596
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13280 3058 13308 4014
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13280 2582 13308 2994
rect 13464 2961 13492 6174
rect 13556 5930 13584 7686
rect 13648 6798 13676 7686
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6254 13676 6734
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13556 5902 13676 5930
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13556 3618 13584 5714
rect 13648 5302 13676 5902
rect 13740 5545 13768 6666
rect 13832 6089 13860 8978
rect 13818 6080 13874 6089
rect 13818 6015 13874 6024
rect 13726 5536 13782 5545
rect 13726 5471 13782 5480
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13556 3590 13676 3618
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13450 2952 13506 2961
rect 13450 2887 13506 2896
rect 13556 2854 13584 3470
rect 13648 3194 13676 3590
rect 13740 3534 13768 4490
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4214 13860 4422
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13924 4010 13952 9318
rect 14016 6934 14044 9522
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 14016 5574 14044 6870
rect 14108 6118 14136 9676
rect 14200 9654 14228 11308
rect 14278 11248 14334 11257
rect 14278 11183 14334 11192
rect 14292 11150 14320 11183
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14384 10996 14412 11766
rect 14292 10968 14412 10996
rect 14292 9654 14320 10968
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 9761 14412 10610
rect 14370 9752 14426 9761
rect 14370 9687 14426 9696
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14280 9648 14332 9654
rect 14476 9602 14504 12378
rect 14280 9590 14332 9596
rect 14200 8566 14228 9590
rect 14384 9574 14504 9602
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 7886 14228 8366
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14108 5370 14136 5578
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14200 5166 14228 7278
rect 14292 6089 14320 8842
rect 14384 7206 14412 9574
rect 14568 9518 14596 13246
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14476 9364 14504 9454
rect 14476 9336 14596 9364
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 8945 14504 9114
rect 14568 8974 14596 9336
rect 14660 9178 14688 14311
rect 14752 12986 14780 14962
rect 15028 14521 15056 15098
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15014 14512 15070 14521
rect 15014 14447 15070 14456
rect 15120 14414 15148 14826
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 15106 12880 15162 12889
rect 14740 12844 14792 12850
rect 15106 12815 15108 12824
rect 14740 12786 14792 12792
rect 15160 12815 15162 12824
rect 15108 12786 15160 12792
rect 14752 11218 14780 12786
rect 15108 12368 15160 12374
rect 15106 12336 15108 12345
rect 15160 12336 15162 12345
rect 15106 12271 15162 12280
rect 15108 12232 15160 12238
rect 14936 12192 15108 12220
rect 14832 12164 14884 12170
rect 14936 12152 14964 12192
rect 15108 12174 15160 12180
rect 15212 12170 15240 16050
rect 15304 15366 15332 17983
rect 15396 17882 15424 18158
rect 15488 17921 15516 19382
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15474 17912 15530 17921
rect 15384 17876 15436 17882
rect 15474 17847 15530 17856
rect 15384 17818 15436 17824
rect 15396 17626 15424 17818
rect 15396 17598 15516 17626
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15396 16726 15424 17478
rect 15488 17066 15516 17598
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15396 16153 15424 16662
rect 15382 16144 15438 16153
rect 15382 16079 15438 16088
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 13734 15332 14758
rect 15396 14346 15424 16079
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15488 13870 15516 16730
rect 15580 16114 15608 19110
rect 15672 19009 15700 19314
rect 15658 19000 15714 19009
rect 15658 18935 15714 18944
rect 15658 18456 15714 18465
rect 15658 18391 15714 18400
rect 15672 18290 15700 18391
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15672 18057 15700 18226
rect 15658 18048 15714 18057
rect 15658 17983 15714 17992
rect 15660 17808 15712 17814
rect 15658 17776 15660 17785
rect 15712 17776 15714 17785
rect 15658 17711 15714 17720
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15672 15502 15700 17478
rect 15764 16114 15792 19722
rect 15856 19281 15884 19790
rect 15948 19310 15976 19790
rect 15936 19304 15988 19310
rect 15842 19272 15898 19281
rect 15936 19246 15988 19252
rect 15842 19207 15898 19216
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 13938 15608 15302
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15658 14784 15714 14793
rect 15658 14719 15714 14728
rect 15672 14006 15700 14719
rect 15764 14618 15792 14962
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15856 14074 15884 19110
rect 16040 18057 16068 20046
rect 16132 18154 16160 24074
rect 16224 23526 16252 24142
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16316 23633 16344 23734
rect 16302 23624 16358 23633
rect 16302 23559 16358 23568
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16408 23322 16436 24686
rect 16500 24206 16528 25094
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16486 24032 16542 24041
rect 16486 23967 16542 23976
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16224 21690 16252 23054
rect 16408 22642 16436 23258
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16500 21554 16528 23967
rect 16592 23497 16620 26794
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16578 23488 16634 23497
rect 16578 23423 16634 23432
rect 16684 23066 16712 25842
rect 16776 23186 16804 28018
rect 16868 27130 16896 31690
rect 16960 29578 16988 32524
rect 17144 32450 17172 32846
rect 17052 32422 17172 32450
rect 17052 30954 17080 32422
rect 17130 31920 17186 31929
rect 17130 31855 17186 31864
rect 17144 31822 17172 31855
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17236 31142 17264 32966
rect 17328 32842 17356 33186
rect 19168 33114 19196 33526
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 17316 32836 17368 32842
rect 17316 32778 17368 32784
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17052 30926 17172 30954
rect 17144 30326 17172 30926
rect 17328 30784 17356 32370
rect 17408 32292 17460 32298
rect 17408 32234 17460 32240
rect 17420 31929 17448 32234
rect 17590 32192 17646 32201
rect 17590 32127 17646 32136
rect 17498 32056 17554 32065
rect 17498 31991 17554 32000
rect 17406 31920 17462 31929
rect 17406 31855 17462 31864
rect 17512 31736 17540 31991
rect 17604 31958 17632 32127
rect 18064 32065 18092 32370
rect 18315 32124 18623 32133
rect 18315 32122 18321 32124
rect 18377 32122 18401 32124
rect 18457 32122 18481 32124
rect 18537 32122 18561 32124
rect 18617 32122 18623 32124
rect 18377 32070 18379 32122
rect 18559 32070 18561 32122
rect 18315 32068 18321 32070
rect 18377 32068 18401 32070
rect 18457 32068 18481 32070
rect 18537 32068 18561 32070
rect 18617 32068 18623 32070
rect 18050 32056 18106 32065
rect 18315 32059 18623 32068
rect 18050 31991 18106 32000
rect 17592 31952 17644 31958
rect 17592 31894 17644 31900
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18418 31920 18474 31929
rect 17420 31708 17540 31736
rect 17684 31748 17736 31754
rect 17420 31482 17448 31708
rect 17684 31690 17736 31696
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17236 30756 17356 30784
rect 17236 30410 17264 30756
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17236 30382 17356 30410
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29646 17172 29990
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 17144 29170 17172 29582
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17052 28558 17080 29106
rect 17236 29102 17264 29582
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 17328 27418 17356 30382
rect 17420 28694 17448 30534
rect 17512 30054 17540 31214
rect 17696 30802 17724 31690
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17788 30734 17816 31622
rect 18248 30938 18276 31894
rect 18418 31855 18474 31864
rect 18432 31822 18460 31855
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 18696 31136 18748 31142
rect 18696 31078 18748 31084
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 18236 30932 18288 30938
rect 18236 30874 18288 30880
rect 18052 30796 18104 30802
rect 18052 30738 18104 30744
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17684 30388 17736 30394
rect 17684 30330 17736 30336
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17408 28688 17460 28694
rect 17408 28630 17460 28636
rect 17408 28144 17460 28150
rect 17408 28086 17460 28092
rect 17144 27390 17356 27418
rect 17038 27160 17094 27169
rect 16856 27124 16908 27130
rect 17038 27095 17094 27104
rect 16856 27066 16908 27072
rect 17052 26994 17080 27095
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 16948 25968 17000 25974
rect 17052 25956 17080 26930
rect 17000 25928 17080 25956
rect 16948 25910 17000 25916
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16868 23798 16896 25230
rect 16946 24984 17002 24993
rect 16946 24919 17002 24928
rect 16960 24682 16988 24919
rect 16948 24676 17000 24682
rect 16948 24618 17000 24624
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16960 24070 16988 24210
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 17144 23361 17172 27390
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26858 17264 26930
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17328 26382 17356 27270
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17130 23352 17186 23361
rect 17130 23287 17186 23296
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 17132 23112 17184 23118
rect 16580 23044 16632 23050
rect 16684 23038 16804 23066
rect 17132 23054 17184 23060
rect 16580 22986 16632 22992
rect 16592 22710 16620 22986
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16776 22094 16804 23038
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16868 22642 16896 22918
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16684 22066 16804 22094
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 21146 16528 21490
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16210 20088 16266 20097
rect 16210 20023 16212 20032
rect 16264 20023 16266 20032
rect 16212 19994 16264 20000
rect 16316 19854 16344 20742
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16304 19848 16356 19854
rect 16210 19816 16266 19825
rect 16304 19790 16356 19796
rect 16210 19751 16266 19760
rect 16224 19514 16252 19751
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16396 19440 16448 19446
rect 16210 19408 16266 19417
rect 16210 19343 16212 19352
rect 16264 19343 16266 19352
rect 16316 19388 16396 19394
rect 16316 19382 16448 19388
rect 16316 19366 16436 19382
rect 16212 19314 16264 19320
rect 16210 19000 16266 19009
rect 16210 18935 16266 18944
rect 16224 18902 16252 18935
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16212 18080 16264 18086
rect 16026 18048 16082 18057
rect 16212 18022 16264 18028
rect 16026 17983 16082 17992
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 16794 15976 17614
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 16040 16969 16068 17546
rect 16026 16960 16082 16969
rect 16026 16895 16082 16904
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16040 15706 16068 16895
rect 16132 16590 16160 17711
rect 16224 17202 16252 18022
rect 16316 17610 16344 19366
rect 16394 18864 16450 18873
rect 16394 18799 16450 18808
rect 16408 18766 16436 18799
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16408 18193 16436 18226
rect 16394 18184 16450 18193
rect 16394 18119 16450 18128
rect 16394 17912 16450 17921
rect 16394 17847 16396 17856
rect 16448 17847 16450 17856
rect 16396 17818 16448 17824
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16302 17368 16358 17377
rect 16302 17303 16304 17312
rect 16356 17303 16358 17312
rect 16304 17274 16356 17280
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16408 17105 16436 17478
rect 16500 17338 16528 20402
rect 16592 17626 16620 21966
rect 16684 19990 16712 22066
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16684 19417 16712 19450
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16776 18970 16804 21830
rect 16868 20466 16896 22578
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16960 20924 16988 21558
rect 17052 21350 17080 22578
rect 17144 21962 17172 23054
rect 17236 22234 17264 25094
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17328 24313 17356 24346
rect 17420 24342 17448 28086
rect 17604 27962 17632 29990
rect 17512 27934 17632 27962
rect 17512 25906 17540 27934
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17408 24336 17460 24342
rect 17314 24304 17370 24313
rect 17408 24278 17460 24284
rect 17314 24239 17370 24248
rect 17420 24154 17448 24278
rect 17328 24126 17448 24154
rect 17328 24041 17356 24126
rect 17408 24064 17460 24070
rect 17314 24032 17370 24041
rect 17408 24006 17460 24012
rect 17314 23967 17370 23976
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17328 23662 17356 23734
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 17420 23474 17448 24006
rect 17328 23446 17448 23474
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17328 22137 17356 23446
rect 17604 23322 17632 27814
rect 17696 26790 17724 30330
rect 17880 29850 17908 30602
rect 17972 30025 18000 30670
rect 18064 30433 18092 30738
rect 18050 30424 18106 30433
rect 18708 30394 18736 31078
rect 18800 30938 18828 31622
rect 18878 31512 18934 31521
rect 19076 31482 19104 33050
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 18878 31447 18934 31456
rect 19064 31476 19116 31482
rect 18892 30938 18920 31447
rect 19064 31418 19116 31424
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 18970 30832 19026 30841
rect 18970 30767 19026 30776
rect 18984 30569 19012 30767
rect 18970 30560 19026 30569
rect 18970 30495 19026 30504
rect 18050 30359 18106 30368
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 18156 30054 18184 30262
rect 18236 30184 18288 30190
rect 18236 30126 18288 30132
rect 18144 30048 18196 30054
rect 17958 30016 18014 30025
rect 18144 29990 18196 29996
rect 17958 29951 18014 29960
rect 17868 29844 17920 29850
rect 17868 29786 17920 29792
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 17958 28792 18014 28801
rect 17958 28727 18014 28736
rect 17972 28694 18000 28727
rect 17960 28688 18012 28694
rect 17960 28630 18012 28636
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 17880 27470 17908 28494
rect 18064 27674 18092 29786
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17868 27464 17920 27470
rect 17788 27424 17868 27452
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17696 25226 17724 26386
rect 17788 25838 17816 27424
rect 17868 27406 17920 27412
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 17972 26994 18000 27066
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17880 26790 17908 26862
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17960 26512 18012 26518
rect 17960 26454 18012 26460
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17696 23633 17724 24754
rect 17788 24750 17816 25774
rect 17880 25498 17908 25842
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17972 24682 18000 26454
rect 18064 25362 18092 26930
rect 18156 26761 18184 29174
rect 18248 28966 18276 30126
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 18604 29232 18656 29238
rect 18604 29174 18656 29180
rect 18972 29232 19024 29238
rect 18972 29174 19024 29180
rect 18616 28966 18644 29174
rect 18984 28994 19012 29174
rect 18892 28966 19012 28994
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 18236 28960 18288 28966
rect 18236 28902 18288 28908
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18694 28928 18750 28937
rect 18248 28608 18276 28902
rect 18315 28860 18623 28869
rect 18694 28863 18750 28872
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18708 28694 18736 28863
rect 18696 28688 18748 28694
rect 18696 28630 18748 28636
rect 18248 28580 18368 28608
rect 18340 28490 18368 28580
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18142 26752 18198 26761
rect 18142 26687 18198 26696
rect 18248 25838 18276 28426
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18326 28248 18382 28257
rect 18326 28183 18382 28192
rect 18510 28248 18566 28257
rect 18510 28183 18566 28192
rect 18340 27946 18368 28183
rect 18524 28150 18552 28183
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18328 27940 18380 27946
rect 18328 27882 18380 27888
rect 18708 27826 18736 28358
rect 18892 28132 18920 28966
rect 18972 28688 19024 28694
rect 18972 28630 19024 28636
rect 18984 28218 19012 28630
rect 19062 28248 19118 28257
rect 18972 28212 19024 28218
rect 19062 28183 19118 28192
rect 18972 28154 19024 28160
rect 18800 28104 18920 28132
rect 18800 27928 18828 28104
rect 19076 28082 19104 28183
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 18800 27900 19012 27928
rect 18708 27798 18828 27826
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 18694 27704 18750 27713
rect 18694 27639 18750 27648
rect 18420 27396 18472 27402
rect 18420 27338 18472 27344
rect 18432 26926 18460 27338
rect 18708 27305 18736 27639
rect 18694 27296 18750 27305
rect 18694 27231 18750 27240
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18696 26920 18748 26926
rect 18800 26908 18828 27798
rect 18984 27169 19012 27900
rect 19064 27872 19116 27878
rect 19062 27840 19064 27849
rect 19116 27840 19118 27849
rect 19062 27775 19118 27784
rect 19062 27704 19118 27713
rect 19062 27639 19118 27648
rect 18970 27160 19026 27169
rect 19076 27130 19104 27639
rect 18970 27095 19026 27104
rect 19064 27124 19116 27130
rect 18748 26880 18828 26908
rect 18696 26862 18748 26868
rect 18432 26772 18460 26862
rect 18432 26744 18736 26772
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18616 25838 18644 25910
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 18052 25220 18104 25226
rect 18052 25162 18104 25168
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24410 17816 24550
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17972 23866 18000 24142
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18064 23798 18092 25162
rect 18156 24206 18184 25706
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18236 24336 18288 24342
rect 18236 24278 18288 24284
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18248 24206 18276 24278
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17682 23624 17738 23633
rect 17682 23559 17738 23568
rect 17592 23316 17644 23322
rect 17420 23276 17592 23304
rect 17420 22574 17448 23276
rect 17592 23258 17644 23264
rect 17696 23118 17724 23559
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17314 22128 17370 22137
rect 17314 22063 17370 22072
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17040 20936 17092 20942
rect 16960 20896 17040 20924
rect 17040 20878 17092 20884
rect 16946 20768 17002 20777
rect 16946 20703 17002 20712
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16868 18222 16896 18838
rect 16960 18426 16988 20703
rect 17052 18737 17080 20878
rect 17144 19446 17172 21898
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17224 21616 17276 21622
rect 17420 21570 17448 21830
rect 17224 21558 17276 21564
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17236 19334 17264 21558
rect 17328 21554 17448 21570
rect 17316 21548 17448 21554
rect 17368 21542 17448 21548
rect 17316 21490 17368 21496
rect 17328 20777 17356 21490
rect 17512 20874 17540 22646
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17604 22234 17632 22442
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17696 20874 17724 23054
rect 17788 22778 17816 23666
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 17776 22636 17828 22642
rect 17880 22624 17908 23054
rect 18064 22794 18092 23734
rect 17972 22778 18092 22794
rect 17960 22772 18092 22778
rect 18012 22766 18092 22772
rect 17960 22714 18012 22720
rect 18052 22704 18104 22710
rect 17828 22596 17908 22624
rect 17972 22652 18052 22658
rect 17972 22646 18104 22652
rect 17972 22630 18092 22646
rect 17776 22578 17828 22584
rect 17774 22128 17830 22137
rect 17774 22063 17830 22072
rect 17788 21078 17816 22063
rect 17972 21146 18000 22630
rect 18156 22438 18184 23802
rect 18340 23508 18368 24278
rect 18708 23866 18736 26744
rect 18800 26246 18828 26880
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 18800 24682 18828 26182
rect 18984 25226 19012 27095
rect 19064 27066 19116 27072
rect 18972 25220 19024 25226
rect 18892 25180 18972 25208
rect 18788 24676 18840 24682
rect 18788 24618 18840 24624
rect 18892 24342 18920 25180
rect 18972 25162 19024 25168
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18984 24274 19012 24550
rect 19076 24342 19104 24754
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18248 23480 18368 23508
rect 18248 22642 18276 23480
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18694 23352 18750 23361
rect 18616 23296 18694 23304
rect 18616 23287 18750 23296
rect 18616 23276 18736 23287
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17776 21072 17828 21078
rect 17776 21014 17828 21020
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17776 20800 17828 20806
rect 17314 20768 17370 20777
rect 17776 20742 17828 20748
rect 17314 20703 17370 20712
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17512 20369 17540 20402
rect 17592 20392 17644 20398
rect 17498 20360 17554 20369
rect 17644 20352 17724 20380
rect 17592 20334 17644 20340
rect 17498 20295 17554 20304
rect 17512 19854 17540 20295
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17144 19306 17264 19334
rect 17038 18728 17094 18737
rect 17038 18663 17094 18672
rect 17144 18630 17172 19306
rect 17328 18766 17356 19722
rect 17316 18760 17368 18766
rect 17236 18720 17316 18748
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 16592 17598 16712 17626
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16394 17096 16450 17105
rect 16316 17054 16394 17082
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16040 15065 16068 15098
rect 16026 15056 16082 15065
rect 16026 14991 16082 15000
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14884 12124 14964 12152
rect 15200 12164 15252 12170
rect 14832 12106 14884 12112
rect 15200 12106 15252 12112
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14844 11393 14872 11698
rect 14830 11384 14886 11393
rect 14936 11354 14964 11698
rect 14830 11319 14886 11328
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14844 10996 14872 11154
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 14752 10968 14872 10996
rect 14752 9178 14780 10968
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 15212 10810 15240 11018
rect 15304 10810 15332 12582
rect 15382 11928 15438 11937
rect 15488 11898 15516 13194
rect 15672 13161 15700 13670
rect 15658 13152 15714 13161
rect 15658 13087 15714 13096
rect 15764 13002 15792 13806
rect 15672 12974 15792 13002
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12753 15608 12786
rect 15566 12744 15622 12753
rect 15566 12679 15622 12688
rect 15672 12628 15700 12974
rect 15580 12600 15700 12628
rect 15752 12640 15804 12646
rect 15580 12238 15608 12600
rect 15752 12582 15804 12588
rect 15568 12232 15620 12238
rect 15566 12200 15568 12209
rect 15660 12232 15712 12238
rect 15620 12200 15622 12209
rect 15660 12174 15712 12180
rect 15566 12135 15622 12144
rect 15566 12064 15622 12073
rect 15566 11999 15622 12008
rect 15382 11863 15438 11872
rect 15476 11892 15528 11898
rect 15396 11830 15424 11863
rect 15476 11834 15528 11840
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15580 11762 15608 11999
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15672 11642 15700 12174
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15580 11614 15700 11642
rect 15396 11257 15424 11562
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15212 10690 15240 10746
rect 15212 10674 15424 10690
rect 15108 10668 15160 10674
rect 15212 10668 15436 10674
rect 15212 10662 15384 10668
rect 15108 10610 15160 10616
rect 15384 10610 15436 10616
rect 15120 10305 15148 10610
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15106 10296 15162 10305
rect 15106 10231 15162 10240
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14844 9058 14872 9658
rect 15108 9648 15160 9654
rect 15106 9616 15108 9625
rect 15160 9616 15162 9625
rect 15106 9551 15162 9560
rect 15108 9512 15160 9518
rect 15014 9480 15070 9489
rect 15108 9454 15160 9460
rect 15014 9415 15070 9424
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14660 9030 14872 9058
rect 14556 8968 14608 8974
rect 14462 8936 14518 8945
rect 14556 8910 14608 8916
rect 14462 8871 14518 8880
rect 14476 8498 14504 8871
rect 14660 8786 14688 9030
rect 14936 8888 14964 9114
rect 15028 9042 15056 9415
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14568 8758 14688 8786
rect 14752 8860 14964 8888
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 7886 14504 8298
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14278 6080 14334 6089
rect 14278 6015 14334 6024
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14292 5545 14320 5578
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14384 4622 14412 6598
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 1970 13308 2518
rect 13740 2446 13768 3334
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 14292 1834 14320 3946
rect 14384 3194 14412 4558
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14476 2774 14504 6938
rect 14568 6118 14596 8758
rect 14752 8634 14780 8860
rect 15120 8838 15148 9454
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 8401 14688 8434
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 15120 8090 15148 8191
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14660 6662 14688 7414
rect 14738 7304 14794 7313
rect 14738 7239 14794 7248
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6186 14688 6598
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14568 4622 14596 5714
rect 14752 5352 14780 7239
rect 14844 7002 14872 7414
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 15028 6934 15056 7346
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15120 6798 15148 6870
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 15212 6458 15240 10406
rect 15304 10266 15332 10406
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15292 9512 15344 9518
rect 15290 9480 15292 9489
rect 15344 9480 15346 9489
rect 15290 9415 15346 9424
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8498 15332 9318
rect 15396 8566 15424 10610
rect 15488 9722 15516 11290
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15474 9208 15530 9217
rect 15474 9143 15476 9152
rect 15528 9143 15530 9152
rect 15476 9114 15528 9120
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15488 8412 15516 8910
rect 15580 8634 15608 11614
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15672 10266 15700 11222
rect 15764 10606 15792 12582
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11286 15884 12038
rect 15948 11354 15976 14758
rect 16132 14618 16160 14826
rect 16224 14618 16252 16050
rect 16316 15570 16344 17054
rect 16394 17031 16450 17040
rect 16396 16584 16448 16590
rect 16394 16552 16396 16561
rect 16448 16552 16450 16561
rect 16394 16487 16450 16496
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16302 15328 16358 15337
rect 16302 15263 16358 15272
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16040 14056 16068 14486
rect 16040 14028 16252 14056
rect 16118 13968 16174 13977
rect 16028 13932 16080 13938
rect 16118 13903 16174 13912
rect 16028 13874 16080 13880
rect 16040 13326 16068 13874
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12073 16068 13126
rect 16026 12064 16082 12073
rect 16026 11999 16082 12008
rect 16026 11928 16082 11937
rect 16026 11863 16082 11872
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15934 11248 15990 11257
rect 15934 11183 15990 11192
rect 15948 11082 15976 11183
rect 16040 11082 16068 11863
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15856 9674 15884 10950
rect 15948 10713 15976 11018
rect 16132 11014 16160 13903
rect 16224 13274 16252 14028
rect 16316 13705 16344 15263
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16302 13696 16358 13705
rect 16302 13631 16358 13640
rect 16224 13246 16344 13274
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16224 12850 16252 13126
rect 16316 12918 16344 13246
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16224 12594 16252 12786
rect 16224 12566 16344 12594
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16118 10840 16174 10849
rect 16118 10775 16174 10784
rect 16132 10742 16160 10775
rect 16120 10736 16172 10742
rect 15934 10704 15990 10713
rect 15934 10639 15990 10648
rect 16040 10696 16120 10724
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15672 9646 15884 9674
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15396 8384 15516 8412
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15304 6390 15332 7210
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14832 6248 14884 6254
rect 15212 6225 15240 6258
rect 15292 6248 15344 6254
rect 14832 6190 14884 6196
rect 15198 6216 15254 6225
rect 14844 5778 14872 6190
rect 15292 6190 15344 6196
rect 15198 6151 15254 6160
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 15200 5704 15252 5710
rect 15198 5672 15200 5681
rect 15252 5672 15254 5681
rect 15198 5607 15254 5616
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14832 5364 14884 5370
rect 14752 5324 14832 5352
rect 14832 5306 14884 5312
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 15304 4536 15332 6190
rect 15396 5012 15424 8384
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15474 7032 15530 7041
rect 15474 6967 15476 6976
rect 15528 6967 15530 6976
rect 15476 6938 15528 6944
rect 15474 6760 15530 6769
rect 15474 6695 15476 6704
rect 15528 6695 15530 6704
rect 15476 6666 15528 6672
rect 15474 6488 15530 6497
rect 15474 6423 15530 6432
rect 15488 6322 15516 6423
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5574 15516 6258
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5166 15516 5510
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15396 4984 15516 5012
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15212 4508 15332 4536
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14476 2746 14596 2774
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 12256 1828 12308 1834
rect 12256 1770 12308 1776
rect 12716 1828 12768 1834
rect 12716 1770 12768 1776
rect 14280 1828 14332 1834
rect 14280 1770 14332 1776
rect 14476 1426 14504 1974
rect 14568 1494 14596 2746
rect 14660 2446 14688 4422
rect 14752 4214 14780 4422
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 15212 2514 15240 4508
rect 15396 4282 15424 4626
rect 15488 4554 15516 4984
rect 15580 4758 15608 8230
rect 15672 6746 15700 9646
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 9382 15792 9522
rect 15948 9518 15976 9862
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15752 9376 15804 9382
rect 15750 9344 15752 9353
rect 15804 9344 15806 9353
rect 15750 9279 15806 9288
rect 15856 8634 15884 9386
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15948 8430 15976 9454
rect 16040 8838 16068 10696
rect 16120 10678 16172 10684
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 9489 16160 9998
rect 16118 9480 16174 9489
rect 16118 9415 16174 9424
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16028 8560 16080 8566
rect 16132 8537 16160 9318
rect 16028 8502 16080 8508
rect 16118 8528 16174 8537
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15948 7954 15976 8366
rect 16040 8022 16068 8502
rect 16118 8463 16174 8472
rect 16224 8022 16252 11494
rect 16316 10248 16344 12566
rect 16408 12374 16436 14350
rect 16500 12986 16528 15574
rect 16592 15026 16620 17478
rect 16684 17134 16712 17598
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16590 16712 17070
rect 16776 16998 16804 17750
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16580 14408 16632 14414
rect 16684 14385 16712 16390
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16580 14350 16632 14356
rect 16670 14376 16726 14385
rect 16592 14074 16620 14350
rect 16670 14311 16726 14320
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16776 13546 16804 15506
rect 16868 15366 16896 17478
rect 16960 17105 16988 18362
rect 17052 18329 17080 18362
rect 17038 18320 17094 18329
rect 17038 18255 17094 18264
rect 17130 17912 17186 17921
rect 17130 17847 17186 17856
rect 17144 17610 17172 17847
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17144 17241 17172 17546
rect 17130 17232 17186 17241
rect 17040 17196 17092 17202
rect 17130 17167 17186 17176
rect 17040 17138 17092 17144
rect 16946 17096 17002 17105
rect 16946 17031 17002 17040
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16960 16658 16988 16730
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16856 15088 16908 15094
rect 16856 15030 16908 15036
rect 16868 13938 16896 15030
rect 16960 14657 16988 16390
rect 17052 15094 17080 17138
rect 17144 16697 17172 17167
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17236 15978 17264 18720
rect 17316 18702 17368 18708
rect 17314 17640 17370 17649
rect 17314 17575 17370 17584
rect 17328 17270 17356 17575
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17314 17096 17370 17105
rect 17314 17031 17370 17040
rect 17328 16590 17356 17031
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 17236 15570 17264 15914
rect 17224 15564 17276 15570
rect 17144 15524 17224 15552
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16946 14648 17002 14657
rect 16946 14583 17002 14592
rect 17052 14482 17080 14894
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17144 14414 17172 15524
rect 17224 15506 17276 15512
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17130 13968 17186 13977
rect 16856 13932 16908 13938
rect 17130 13903 17186 13912
rect 16856 13874 16908 13880
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16592 13518 16804 13546
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16592 12102 16620 13518
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16854 13424 16910 13433
rect 16684 12442 16712 13398
rect 16854 13359 16910 13368
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 10674 16528 11834
rect 16592 11529 16620 12038
rect 16776 11762 16804 13126
rect 16868 12442 16896 13359
rect 16960 13258 16988 13738
rect 17144 13734 17172 13903
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17038 13424 17094 13433
rect 17038 13359 17094 13368
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 17052 12850 17080 13359
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16578 11520 16634 11529
rect 16578 11455 16634 11464
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16580 10260 16632 10266
rect 16316 10220 16436 10248
rect 16302 10160 16358 10169
rect 16302 10095 16358 10104
rect 16316 10062 16344 10095
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16302 8936 16358 8945
rect 16302 8871 16358 8880
rect 16316 8838 16344 8871
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15856 7750 15884 7890
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16120 7880 16172 7886
rect 16316 7834 16344 8570
rect 16120 7822 16172 7828
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 16040 7546 16068 7822
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16132 7290 16160 7822
rect 16040 7262 16160 7290
rect 16224 7806 16344 7834
rect 15844 6792 15896 6798
rect 15672 6718 15792 6746
rect 15844 6734 15896 6740
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 5234 15700 6598
rect 15764 6497 15792 6718
rect 15750 6488 15806 6497
rect 15750 6423 15806 6432
rect 15752 6316 15804 6322
rect 15856 6304 15884 6734
rect 15804 6276 15884 6304
rect 15752 6258 15804 6264
rect 16040 6225 16068 7262
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6730 16160 7142
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16224 6322 16252 7806
rect 16408 7478 16436 10220
rect 16580 10202 16632 10208
rect 16486 9616 16542 9625
rect 16486 9551 16488 9560
rect 16540 9551 16542 9560
rect 16488 9522 16540 9528
rect 16486 9208 16542 9217
rect 16486 9143 16542 9152
rect 16500 7886 16528 9143
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16488 6928 16540 6934
rect 16486 6896 16488 6905
rect 16540 6896 16542 6905
rect 16486 6831 16542 6840
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15842 6216 15898 6225
rect 15842 6151 15898 6160
rect 16026 6216 16082 6225
rect 16224 6186 16252 6258
rect 16026 6151 16082 6160
rect 16212 6180 16264 6186
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15304 2446 15332 3334
rect 15396 2650 15424 4014
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3602 15608 3878
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15488 3126 15516 3470
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15488 2582 15516 2926
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15580 2446 15608 3538
rect 15672 3534 15700 4966
rect 15764 4690 15792 5782
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 15108 1760 15160 1766
rect 15108 1702 15160 1708
rect 14556 1488 14608 1494
rect 14556 1430 14608 1436
rect 14464 1420 14516 1426
rect 14464 1362 14516 1368
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 15120 1222 15148 1702
rect 15212 1358 15240 2314
rect 15488 1816 15516 2382
rect 15568 1828 15620 1834
rect 15488 1788 15568 1816
rect 15568 1770 15620 1776
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15108 1216 15160 1222
rect 15108 1158 15160 1164
rect 14842 1116 15150 1125
rect 14842 1114 14848 1116
rect 14904 1114 14928 1116
rect 14984 1114 15008 1116
rect 15064 1114 15088 1116
rect 15144 1114 15150 1116
rect 14904 1062 14906 1114
rect 15086 1062 15088 1114
rect 14842 1060 14848 1062
rect 14904 1060 14928 1062
rect 14984 1060 15008 1062
rect 15064 1060 15088 1062
rect 15144 1060 15150 1062
rect 14842 1051 15150 1060
rect 10968 1012 11020 1018
rect 10968 954 11020 960
rect 9956 944 10008 950
rect 9956 886 10008 892
rect 5908 808 5960 814
rect 5908 750 5960 756
rect 3976 672 4028 678
rect 3976 614 4028 620
rect 15580 610 15608 1770
rect 15672 1426 15700 3062
rect 15856 2854 15884 6151
rect 16212 6122 16264 6128
rect 16026 6080 16082 6089
rect 16026 6015 16082 6024
rect 16040 5574 16068 6015
rect 16224 5778 16252 6122
rect 16592 5953 16620 10202
rect 16684 8430 16712 11290
rect 16868 11082 16896 12174
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16960 10742 16988 12106
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10810 17080 10950
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16960 10554 16988 10678
rect 16960 10526 17080 10554
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 10130 16988 10406
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 17052 10062 17080 10526
rect 17040 10056 17092 10062
rect 16762 10024 16818 10033
rect 17040 9998 17092 10004
rect 16762 9959 16818 9968
rect 16948 9988 17000 9994
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16776 8378 16804 9959
rect 16948 9930 17000 9936
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 8566 16896 9862
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16776 8350 16896 8378
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 6390 16712 7890
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16578 5944 16634 5953
rect 16578 5879 16634 5888
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16592 5642 16620 5879
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16132 4282 16160 5578
rect 16684 5302 16712 6326
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 15856 1358 15884 2790
rect 15948 2038 15976 3402
rect 16408 2650 16436 4694
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16500 2038 16528 3674
rect 16776 3398 16804 8230
rect 16868 6798 16896 8350
rect 16960 7546 16988 9930
rect 17038 9480 17094 9489
rect 17038 9415 17094 9424
rect 17052 9382 17080 9415
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17052 7002 17080 9318
rect 17144 9024 17172 13262
rect 17236 10810 17264 14962
rect 17328 14006 17356 15302
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17328 11937 17356 13942
rect 17420 13705 17448 19790
rect 17592 19372 17644 19378
rect 17696 19360 17724 20352
rect 17788 20058 17816 20742
rect 17880 20466 17908 20878
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17972 20398 18000 20742
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17880 19446 17908 19994
rect 17972 19689 18000 20334
rect 18064 19990 18092 22374
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18156 21622 18184 22170
rect 18248 22137 18276 22578
rect 18524 22506 18552 23190
rect 18616 23050 18644 23276
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22953 18644 22986
rect 18602 22944 18658 22953
rect 18602 22879 18658 22888
rect 18708 22710 18736 23122
rect 18800 22982 18828 23666
rect 18892 23322 18920 24142
rect 19076 24041 19104 24278
rect 19062 24032 19118 24041
rect 19062 23967 19118 23976
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18984 23633 19012 23666
rect 18970 23624 19026 23633
rect 18970 23559 19026 23568
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18984 22760 19012 23559
rect 19168 23254 19196 28970
rect 19260 28014 19288 32846
rect 20444 32496 20496 32502
rect 20444 32438 20496 32444
rect 19432 32360 19484 32366
rect 19432 32302 19484 32308
rect 19444 31822 19472 32302
rect 20456 32230 20484 32438
rect 21192 32230 21220 33594
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 23388 33380 23440 33386
rect 23388 33322 23440 33328
rect 22928 32904 22980 32910
rect 22928 32846 22980 32852
rect 21272 32836 21324 32842
rect 21272 32778 21324 32784
rect 21284 32230 21312 32778
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 21788 32668 22096 32677
rect 21788 32666 21794 32668
rect 21850 32666 21874 32668
rect 21930 32666 21954 32668
rect 22010 32666 22034 32668
rect 22090 32666 22096 32668
rect 21850 32614 21852 32666
rect 22032 32614 22034 32666
rect 21788 32612 21794 32614
rect 21850 32612 21874 32614
rect 21930 32612 21954 32614
rect 22010 32612 22034 32614
rect 22090 32612 22096 32614
rect 21788 32603 22096 32612
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22112 32434 22140 32506
rect 22204 32434 22232 32710
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 19616 32224 19668 32230
rect 19616 32166 19668 32172
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 21180 32224 21232 32230
rect 21180 32166 21232 32172
rect 21272 32224 21324 32230
rect 21272 32166 21324 32172
rect 19432 31816 19484 31822
rect 19352 31764 19432 31770
rect 19352 31758 19484 31764
rect 19352 31742 19472 31758
rect 19352 31278 19380 31742
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19352 30818 19380 31214
rect 19524 30864 19576 30870
rect 19352 30790 19472 30818
rect 19524 30806 19576 30812
rect 19444 30734 19472 30790
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 30190 19472 30670
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19444 29646 19472 30126
rect 19536 29646 19564 30806
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19352 29306 19380 29446
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19444 29170 19472 29582
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19628 28994 19656 32166
rect 20812 31952 20864 31958
rect 20812 31894 20864 31900
rect 20824 31793 20852 31894
rect 21548 31816 21600 31822
rect 20810 31784 20866 31793
rect 21548 31758 21600 31764
rect 20810 31719 20866 31728
rect 21560 31686 21588 31758
rect 22112 31754 22140 32370
rect 22940 31958 22968 32846
rect 22928 31952 22980 31958
rect 22928 31894 22980 31900
rect 22112 31726 22232 31754
rect 21548 31680 21600 31686
rect 20718 31648 20774 31657
rect 21548 31622 21600 31628
rect 20718 31583 20774 31592
rect 20732 31210 20760 31583
rect 21560 31278 21588 31622
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 20720 31204 20772 31210
rect 20720 31146 20772 31152
rect 20996 31204 21048 31210
rect 20996 31146 21048 31152
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20732 30394 20760 30602
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20720 30184 20772 30190
rect 20720 30126 20772 30132
rect 19352 28966 19656 28994
rect 20272 29566 20668 29594
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19260 27606 19288 27950
rect 19248 27600 19300 27606
rect 19248 27542 19300 27548
rect 19352 27452 19380 28966
rect 19708 28960 19760 28966
rect 19708 28902 19760 28908
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19260 27424 19380 27452
rect 19260 26518 19288 27424
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 27130 19380 27270
rect 19444 27130 19472 28018
rect 19536 28014 19564 28494
rect 19720 28490 19748 28902
rect 19708 28484 19760 28490
rect 19708 28426 19760 28432
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19616 27328 19668 27334
rect 19616 27270 19668 27276
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19432 26988 19484 26994
rect 19536 26976 19564 27066
rect 19628 26994 19656 27270
rect 19484 26948 19564 26976
rect 19616 26988 19668 26994
rect 19432 26930 19484 26936
rect 19616 26930 19668 26936
rect 19340 26784 19392 26790
rect 19616 26784 19668 26790
rect 19392 26744 19616 26772
rect 19340 26726 19392 26732
rect 19616 26726 19668 26732
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19432 26376 19484 26382
rect 19484 26324 19564 26330
rect 19432 26318 19564 26324
rect 19444 26302 19564 26318
rect 19812 26314 19840 27950
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19536 26296 19564 26302
rect 19800 26308 19852 26314
rect 19536 26268 19800 26296
rect 19800 26250 19852 26256
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 19260 25498 19288 25774
rect 19340 25696 19392 25702
rect 19444 25650 19472 26182
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19392 25644 19472 25650
rect 19340 25638 19472 25644
rect 19352 25622 19472 25638
rect 19812 25498 19840 25842
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 18800 22732 19012 22760
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18800 22522 18828 22732
rect 19168 22642 19196 22918
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18708 22494 18828 22522
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18234 22128 18290 22137
rect 18234 22063 18290 22072
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 17958 19680 18014 19689
rect 17958 19615 18014 19624
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17776 19372 17828 19378
rect 17696 19332 17776 19360
rect 17592 19314 17644 19320
rect 17776 19314 17828 19320
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18737 17540 19110
rect 17498 18728 17554 18737
rect 17498 18663 17554 18672
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 17377 17540 18226
rect 17604 17610 17632 19314
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17498 17368 17554 17377
rect 17498 17303 17554 17312
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16114 17540 16934
rect 17604 16658 17632 17070
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17512 13802 17540 15642
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17406 13696 17462 13705
rect 17406 13631 17462 13640
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17314 11928 17370 11937
rect 17314 11863 17370 11872
rect 17314 11384 17370 11393
rect 17314 11319 17316 11328
rect 17368 11319 17370 11328
rect 17316 11290 17368 11296
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17236 10033 17264 10134
rect 17222 10024 17278 10033
rect 17222 9959 17224 9968
rect 17276 9959 17278 9968
rect 17224 9930 17276 9936
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 9178 17264 9522
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17144 8996 17264 9024
rect 17236 8634 17264 8996
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17144 7002 17172 7754
rect 17222 7168 17278 7177
rect 17222 7103 17278 7112
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17236 6934 17264 7103
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 6254 16896 6734
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16960 5642 16988 6598
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4214 16896 4966
rect 16960 4690 16988 5578
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5234 17080 5510
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17144 5098 17172 6190
rect 17328 6186 17356 10406
rect 17420 9654 17448 13466
rect 17512 12918 17540 13738
rect 17604 13326 17632 16594
rect 17696 16046 17724 18566
rect 17788 17882 17816 19314
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17788 16658 17816 16730
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17880 16522 17908 18702
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17880 16114 17908 16458
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17684 15904 17736 15910
rect 17776 15904 17828 15910
rect 17684 15846 17736 15852
rect 17774 15872 17776 15881
rect 17828 15872 17830 15881
rect 17696 15638 17724 15846
rect 17774 15807 17830 15816
rect 17880 15706 17908 16050
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 14929 17724 15438
rect 17866 15192 17922 15201
rect 17866 15127 17868 15136
rect 17920 15127 17922 15136
rect 17868 15098 17920 15104
rect 17682 14920 17738 14929
rect 17682 14855 17738 14864
rect 17972 14618 18000 19450
rect 18156 19446 18184 21558
rect 18248 20602 18276 21966
rect 18616 21962 18644 22170
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18328 21888 18380 21894
rect 18326 21856 18328 21865
rect 18380 21856 18382 21865
rect 18326 21791 18382 21800
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18432 21457 18460 21626
rect 18418 21448 18474 21457
rect 18418 21383 18474 21392
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18340 20482 18368 20810
rect 18248 20454 18368 20482
rect 18248 19553 18276 20454
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18234 19544 18290 19553
rect 18234 19479 18290 19488
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18064 19174 18092 19314
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18766 18092 19110
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18064 16658 18092 17546
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 18064 15026 18092 16594
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18156 14958 18184 19246
rect 18248 17490 18276 19479
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18616 19174 18644 19314
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18326 18456 18382 18465
rect 18326 18391 18328 18400
rect 18380 18391 18382 18400
rect 18328 18362 18380 18368
rect 18616 18222 18644 18838
rect 18708 18630 18736 22494
rect 18892 22030 18920 22578
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 19064 22432 19116 22438
rect 19062 22400 19064 22409
rect 19116 22400 19118 22409
rect 19062 22335 19118 22344
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18984 22098 19012 22170
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18878 21720 18934 21729
rect 18878 21655 18934 21664
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18800 17882 18828 21286
rect 18892 21146 18920 21655
rect 19168 21418 19196 22442
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 19062 21040 19118 21049
rect 19062 20975 19118 20984
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18326 17776 18382 17785
rect 18326 17711 18382 17720
rect 18340 17678 18368 17711
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17490 18644 17546
rect 18248 17462 18644 17490
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18142 14512 18198 14521
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 13728 17828 13734
rect 17774 13696 17776 13705
rect 17828 13696 17830 13705
rect 17774 13631 17830 13640
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17597 13320 17649 13326
rect 17597 13262 17649 13268
rect 17604 12918 17632 13262
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17498 12472 17554 12481
rect 17498 12407 17500 12416
rect 17552 12407 17554 12416
rect 17500 12378 17552 12384
rect 17498 11792 17554 11801
rect 17498 11727 17500 11736
rect 17552 11727 17554 11736
rect 17500 11698 17552 11704
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 17236 4758 17264 5850
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 15936 2032 15988 2038
rect 15936 1974 15988 1980
rect 16488 2032 16540 2038
rect 16488 1974 16540 1980
rect 15844 1352 15896 1358
rect 15844 1294 15896 1300
rect 16776 746 16804 3334
rect 16868 3126 16896 4150
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 3738 16988 4082
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 17052 1358 17080 3334
rect 17236 2774 17264 4694
rect 17328 3126 17356 5238
rect 17420 3194 17448 8230
rect 17512 5234 17540 11154
rect 17604 7290 17632 12718
rect 17696 10266 17724 12786
rect 17788 11150 17816 13398
rect 17880 12889 17908 14350
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17972 14006 18000 14282
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17972 13326 18000 13942
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17972 12918 18000 13262
rect 17960 12912 18012 12918
rect 17866 12880 17922 12889
rect 17960 12854 18012 12860
rect 17866 12815 17922 12824
rect 17972 12170 18000 12854
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17866 11928 17922 11937
rect 17866 11863 17922 11872
rect 17960 11892 18012 11898
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10538 17816 10950
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17880 9674 17908 11863
rect 17960 11834 18012 11840
rect 17788 9646 17908 9674
rect 17788 8566 17816 9646
rect 17972 9586 18000 11834
rect 18064 9586 18092 14486
rect 18142 14447 18198 14456
rect 18156 12918 18184 14447
rect 18248 13190 18276 17206
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18602 16688 18658 16697
rect 18708 16674 18736 17138
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18800 16794 18828 17002
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18708 16646 18828 16674
rect 18602 16623 18658 16632
rect 18616 16114 18644 16623
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 16425 18736 16526
rect 18694 16416 18750 16425
rect 18694 16351 18750 16360
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 15434 18460 15506
rect 18708 15434 18736 16351
rect 18800 15434 18828 16646
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18340 15026 18368 15370
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18708 14006 18736 15370
rect 18696 14000 18748 14006
rect 18510 13968 18566 13977
rect 18328 13932 18380 13938
rect 18696 13942 18748 13948
rect 18510 13903 18566 13912
rect 18328 13874 18380 13880
rect 18340 13841 18368 13874
rect 18326 13832 18382 13841
rect 18326 13767 18382 13776
rect 18524 13734 18552 13903
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18708 12968 18736 13942
rect 18786 13832 18842 13841
rect 18786 13767 18842 13776
rect 18800 13326 18828 13767
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18616 12940 18736 12968
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18156 12442 18184 12854
rect 18616 12646 18644 12940
rect 18800 12866 18828 13262
rect 18892 12986 18920 20402
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18984 19446 19012 19994
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17202 19012 17478
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18984 16726 19012 17138
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 19076 16250 19104 20975
rect 19260 20942 19288 25298
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19352 24750 19380 25230
rect 19904 25226 19932 27814
rect 19892 25220 19944 25226
rect 19892 25162 19944 25168
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19524 24744 19576 24750
rect 19524 24686 19576 24692
rect 19338 24576 19394 24585
rect 19338 24511 19394 24520
rect 19352 23118 19380 24511
rect 19536 24410 19564 24686
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19524 24404 19576 24410
rect 19524 24346 19576 24352
rect 19628 24290 19656 24618
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19536 24262 19656 24290
rect 19800 24336 19852 24342
rect 19800 24278 19852 24284
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19444 23050 19472 24210
rect 19536 24138 19564 24262
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19352 22778 19380 22918
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19444 22658 19472 22986
rect 19352 22630 19472 22658
rect 19352 22094 19380 22630
rect 19430 22264 19486 22273
rect 19536 22234 19564 24074
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19628 22710 19656 23666
rect 19706 23488 19762 23497
rect 19706 23423 19762 23432
rect 19720 23254 19748 23423
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19720 22953 19748 23190
rect 19706 22944 19762 22953
rect 19706 22879 19762 22888
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19720 22234 19748 22578
rect 19430 22199 19432 22208
rect 19484 22199 19486 22208
rect 19524 22228 19576 22234
rect 19432 22170 19484 22176
rect 19524 22170 19576 22176
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19720 22094 19748 22170
rect 19352 22066 19564 22094
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 20466 19196 20810
rect 19246 20632 19302 20641
rect 19246 20567 19302 20576
rect 19260 20466 19288 20567
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19168 18272 19196 20402
rect 19246 19680 19302 19689
rect 19246 19615 19302 19624
rect 19260 18970 19288 19615
rect 19352 19310 19380 21966
rect 19536 20398 19564 22066
rect 19628 22066 19748 22094
rect 19628 20942 19656 22066
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19720 21690 19748 21966
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19444 19145 19472 19926
rect 19536 19922 19564 20198
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19430 19136 19486 19145
rect 19430 19071 19486 19080
rect 19338 19000 19394 19009
rect 19248 18964 19300 18970
rect 19338 18935 19394 18944
rect 19248 18906 19300 18912
rect 19352 18766 19380 18935
rect 19536 18816 19564 19722
rect 19628 19009 19656 20742
rect 19614 19000 19670 19009
rect 19614 18935 19670 18944
rect 19536 18788 19656 18816
rect 19340 18760 19392 18766
rect 19628 18748 19656 18788
rect 19628 18720 19672 18748
rect 19340 18702 19392 18708
rect 19432 18624 19484 18630
rect 19644 18578 19672 18720
rect 19432 18566 19484 18572
rect 19444 18358 19472 18566
rect 19536 18550 19672 18578
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18284 19392 18290
rect 19168 18244 19340 18272
rect 19260 17678 19288 18244
rect 19340 18226 19392 18232
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19260 16658 19288 17478
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16504 19288 16594
rect 19168 16476 19288 16504
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 15337 19012 15438
rect 18970 15328 19026 15337
rect 18970 15263 19026 15272
rect 18972 14408 19024 14414
rect 19168 14362 19196 16476
rect 19246 16416 19302 16425
rect 19246 16351 19302 16360
rect 18972 14350 19024 14356
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18708 12838 18828 12866
rect 18878 12880 18934 12889
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18248 12170 18276 12310
rect 18340 12306 18368 12378
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 10826 18184 12038
rect 18418 11928 18474 11937
rect 18418 11863 18474 11872
rect 18432 11694 18460 11863
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18248 11286 18276 11630
rect 18524 11608 18552 12378
rect 18708 12102 18736 12838
rect 18878 12815 18934 12824
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11898 18736 12038
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18800 11626 18828 12718
rect 18788 11620 18840 11626
rect 18524 11580 18736 11608
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18156 10810 18276 10826
rect 18156 10804 18288 10810
rect 18156 10798 18236 10804
rect 18236 10746 18288 10752
rect 18144 10736 18196 10742
rect 18340 10690 18368 10950
rect 18196 10684 18368 10690
rect 18144 10678 18368 10684
rect 18156 10662 18368 10678
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18156 9489 18184 10662
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18142 9480 18198 9489
rect 18142 9415 18198 9424
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17880 7834 17908 8366
rect 17972 8022 18000 9318
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 8090 18092 8230
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17880 7806 18092 7834
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 7313 17908 7346
rect 17866 7304 17922 7313
rect 17604 7262 17724 7290
rect 17696 6474 17724 7262
rect 17866 7239 17922 7248
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17604 6458 17724 6474
rect 17880 6458 17908 6666
rect 17592 6452 17724 6458
rect 17644 6446 17724 6452
rect 17868 6452 17920 6458
rect 17592 6394 17644 6400
rect 17868 6394 17920 6400
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 17604 5846 17632 6122
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17604 4826 17632 5782
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17696 3670 17724 6326
rect 17972 6322 18000 7414
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 4214 17908 6054
rect 17972 5710 18000 6258
rect 18064 6186 18092 7806
rect 18156 7546 18184 8570
rect 18340 8378 18368 8774
rect 18708 8537 18736 11580
rect 18788 11562 18840 11568
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18800 10198 18828 10678
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18892 9654 18920 12815
rect 18984 11898 19012 14350
rect 19076 14346 19196 14362
rect 19064 14340 19196 14346
rect 19116 14334 19196 14340
rect 19064 14282 19116 14288
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19076 13297 19104 14010
rect 19168 13938 19196 14214
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 19168 13138 19196 13874
rect 19260 13258 19288 16351
rect 19352 16250 19380 18022
rect 19536 17678 19564 18550
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19338 16144 19394 16153
rect 19338 16079 19394 16088
rect 19432 16108 19484 16114
rect 19352 13394 19380 16079
rect 19536 16096 19564 17614
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19628 17513 19656 17546
rect 19614 17504 19670 17513
rect 19614 17439 19670 17448
rect 19484 16068 19564 16096
rect 19432 16050 19484 16056
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19168 13110 19288 13138
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19168 12782 19196 12922
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19076 12170 19104 12718
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18892 9489 18920 9590
rect 18878 9480 18934 9489
rect 18878 9415 18934 9424
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18694 8528 18750 8537
rect 18694 8463 18750 8472
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18248 8350 18368 8378
rect 18694 8392 18750 8401
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18248 7342 18276 8350
rect 18694 8327 18750 8336
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18524 7818 18552 8026
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18616 7206 18644 7346
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18248 6390 18276 7142
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18708 6866 18736 8327
rect 18800 8090 18828 8434
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18892 7936 18920 8910
rect 18800 7908 18920 7936
rect 18800 7478 18828 7908
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17972 5302 18000 5646
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 18064 4758 18092 6122
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18708 5817 18736 6258
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18432 5030 18460 5578
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 3120 17368 3126
rect 17368 3068 17540 3074
rect 17316 3062 17540 3068
rect 17328 3046 17540 3062
rect 17236 2746 17448 2774
rect 17420 2650 17448 2746
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17512 2582 17540 3046
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17408 2440 17460 2446
rect 17604 2394 17632 2926
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17460 2388 17632 2394
rect 17408 2382 17632 2388
rect 17420 2366 17632 2382
rect 17420 1970 17448 2366
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17512 2038 17540 2246
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17696 1970 17724 2586
rect 17788 2446 17816 3878
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17880 2514 17908 3606
rect 18248 3534 18276 4422
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18800 3097 18828 6054
rect 18892 5234 18920 7686
rect 18984 6458 19012 10406
rect 19076 8838 19104 11698
rect 19168 8906 19196 12582
rect 19260 11830 19288 13110
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19352 11286 19380 12718
rect 19444 12442 19472 15914
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19628 13870 19656 14350
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19340 11280 19392 11286
rect 19246 11248 19302 11257
rect 19340 11222 19392 11228
rect 19246 11183 19302 11192
rect 19260 11014 19288 11183
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19444 10742 19472 12106
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19352 10470 19380 10610
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19260 10266 19288 10406
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19168 7410 19196 8026
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19260 6866 19288 10066
rect 19444 10062 19472 10678
rect 19536 10606 19564 13126
rect 19628 11121 19656 13670
rect 19720 12986 19748 20946
rect 19812 20942 19840 24278
rect 19904 22982 19932 25162
rect 19996 23866 20024 28154
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20076 27328 20128 27334
rect 20076 27270 20128 27276
rect 20088 26042 20116 27270
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 24954 20116 25842
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 20088 23322 20116 24754
rect 20180 23866 20208 27474
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20272 23730 20300 29566
rect 20640 29510 20668 29566
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20444 28960 20496 28966
rect 20444 28902 20496 28908
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20364 26246 20392 28494
rect 20456 26790 20484 28902
rect 20548 26790 20576 29446
rect 20628 28416 20680 28422
rect 20628 28358 20680 28364
rect 20640 28218 20668 28358
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20640 27334 20668 28018
rect 20732 27606 20760 30126
rect 20916 29306 20944 30194
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20904 27668 20956 27674
rect 20824 27628 20904 27656
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20824 27470 20852 27628
rect 20904 27610 20956 27616
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20442 26616 20498 26625
rect 20442 26551 20498 26560
rect 20352 26240 20404 26246
rect 20352 26182 20404 26188
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19996 22681 20024 23190
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 19982 22672 20038 22681
rect 19982 22607 20038 22616
rect 19890 22128 19946 22137
rect 19890 22063 19946 22072
rect 19904 21622 19932 22063
rect 20088 21865 20116 22986
rect 20180 22001 20208 23054
rect 20272 22817 20300 23666
rect 20456 23594 20484 26551
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20258 22808 20314 22817
rect 20258 22743 20314 22752
rect 20548 22710 20576 25842
rect 20732 25673 20760 26930
rect 20916 26586 20944 27406
rect 21008 27130 21036 31146
rect 21456 31136 21508 31142
rect 21456 31078 21508 31084
rect 21468 30734 21496 31078
rect 21560 30938 21588 31214
rect 21548 30932 21600 30938
rect 21548 30874 21600 30880
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21560 29850 21588 30874
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21088 29096 21140 29102
rect 21088 29038 21140 29044
rect 21100 28762 21128 29038
rect 21468 28762 21496 29106
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 20996 27124 21048 27130
rect 20996 27066 21048 27072
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 20904 26308 20956 26314
rect 20904 26250 20956 26256
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20718 25664 20774 25673
rect 20718 25599 20774 25608
rect 20718 25528 20774 25537
rect 20718 25463 20774 25472
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20640 24410 20668 25298
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20640 22778 20668 23666
rect 20732 23526 20760 25463
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20166 21992 20222 22001
rect 20456 21962 20484 22646
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20534 22128 20590 22137
rect 20534 22063 20590 22072
rect 20166 21927 20222 21936
rect 20444 21956 20496 21962
rect 20074 21856 20130 21865
rect 20074 21791 20130 21800
rect 19892 21616 19944 21622
rect 19892 21558 19944 21564
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19904 20466 19932 20878
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20088 20602 20116 20742
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19812 19854 19840 20334
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 18465 19840 19790
rect 19904 19446 19932 20266
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19798 18456 19854 18465
rect 19798 18391 19854 18400
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19812 17882 19840 18226
rect 19904 18057 19932 18702
rect 19890 18048 19946 18057
rect 19890 17983 19946 17992
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19996 17814 20024 20334
rect 20180 19360 20208 21927
rect 20444 21898 20496 21904
rect 20456 21842 20484 21898
rect 20364 21814 20484 21842
rect 20364 21554 20392 21814
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20364 20856 20392 21490
rect 20456 21457 20484 21490
rect 20442 21448 20498 21457
rect 20442 21383 20498 21392
rect 20456 21350 20484 21383
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20444 20868 20496 20874
rect 20364 20828 20444 20856
rect 20444 20810 20496 20816
rect 20456 20466 20484 20810
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 19786 20484 20402
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20088 19332 20208 19360
rect 20088 18222 20116 19332
rect 20442 19272 20498 19281
rect 20168 19236 20220 19242
rect 20442 19207 20498 19216
rect 20168 19178 20220 19184
rect 20180 19145 20208 19178
rect 20166 19136 20222 19145
rect 20222 19094 20392 19122
rect 20166 19071 20222 19080
rect 20364 18766 20392 19094
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20180 18358 20208 18702
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 17202 20024 17614
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19982 17096 20038 17105
rect 19982 17031 20038 17040
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19904 16289 19932 16594
rect 19890 16280 19946 16289
rect 19890 16215 19946 16224
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 15094 19840 15302
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19708 12436 19760 12442
rect 19812 12434 19840 14758
rect 19904 13938 19932 15030
rect 19996 14958 20024 17031
rect 20088 15570 20116 17546
rect 20180 15638 20208 17682
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19996 14521 20024 14894
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19982 14512 20038 14521
rect 20088 14482 20116 14758
rect 19982 14447 20038 14456
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19982 14376 20038 14385
rect 19982 14311 20038 14320
rect 19996 13938 20024 14311
rect 20180 14278 20208 15438
rect 20272 14822 20300 18634
rect 20350 18456 20406 18465
rect 20350 18391 20406 18400
rect 20364 16454 20392 18391
rect 20456 17338 20484 19207
rect 20548 17785 20576 22063
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 20330 20668 20402
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20640 20233 20668 20266
rect 20626 20224 20682 20233
rect 20626 20159 20682 20168
rect 20732 20058 20760 22578
rect 20824 22098 20852 26182
rect 20916 25498 20944 26250
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21008 25974 21036 26182
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 21100 25650 21128 26522
rect 21192 25838 21220 26930
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 21008 25622 21128 25650
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 21008 24614 21036 25622
rect 21284 25430 21312 28494
rect 21456 28212 21508 28218
rect 21456 28154 21508 28160
rect 21362 27568 21418 27577
rect 21362 27503 21418 27512
rect 21376 27470 21404 27503
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21468 26874 21496 28154
rect 21560 27606 21588 29174
rect 21548 27600 21600 27606
rect 21548 27542 21600 27548
rect 21546 27432 21602 27441
rect 21652 27402 21680 31282
rect 21744 30666 21772 31418
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 22204 30394 22232 31726
rect 23400 31686 23428 33322
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 23492 32434 23520 33050
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 21916 30048 21968 30054
rect 21916 29990 21968 29996
rect 21928 29646 21956 29990
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 22296 29306 22324 30874
rect 23584 30734 23612 32302
rect 23676 31890 23704 32982
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23940 31748 23992 31754
rect 23940 31690 23992 31696
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22112 28490 22140 29106
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 22388 28150 22416 30534
rect 23216 30394 23244 30670
rect 23204 30388 23256 30394
rect 23204 30330 23256 30336
rect 22560 30184 22612 30190
rect 22560 30126 22612 30132
rect 22572 29850 22600 30126
rect 22744 30116 22796 30122
rect 22744 30058 22796 30064
rect 22756 29850 22784 30058
rect 23020 30048 23072 30054
rect 23020 29990 23072 29996
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 22020 27470 22048 27542
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 21546 27367 21602 27376
rect 21640 27396 21692 27402
rect 21560 27334 21588 27367
rect 21640 27338 21692 27344
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 21376 26846 21496 26874
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21272 25424 21324 25430
rect 21272 25366 21324 25372
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20916 24274 20944 24550
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20902 21992 20958 22001
rect 20902 21927 20904 21936
rect 20956 21927 20958 21936
rect 20904 21898 20956 21904
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20640 18426 20668 19246
rect 20732 18834 20760 19790
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20824 18630 20852 20810
rect 20916 19174 20944 21898
rect 21008 21486 21036 24278
rect 21100 22098 21128 25230
rect 21376 24936 21404 26846
rect 21454 26752 21510 26761
rect 21454 26687 21510 26696
rect 21192 24908 21404 24936
rect 21192 23905 21220 24908
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21376 24070 21404 24754
rect 21468 24342 21496 26687
rect 21560 25838 21588 26862
rect 21652 26625 21680 26998
rect 21638 26616 21694 26625
rect 21638 26551 21694 26560
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 26217 21680 26250
rect 22204 26217 22232 27270
rect 22296 26382 22324 27270
rect 22388 27062 22416 27338
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22468 26376 22520 26382
rect 22468 26318 22520 26324
rect 21638 26208 21694 26217
rect 21638 26143 21694 26152
rect 22190 26208 22246 26217
rect 21788 26140 22096 26149
rect 22190 26143 22246 26152
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 21560 24750 21588 25774
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22020 25498 22048 25638
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 21456 24336 21508 24342
rect 21456 24278 21508 24284
rect 22020 24274 22048 24686
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21178 23896 21234 23905
rect 21178 23831 21234 23840
rect 21284 23594 21312 24006
rect 21272 23588 21324 23594
rect 21272 23530 21324 23536
rect 21088 22092 21140 22098
rect 21560 22094 21588 24210
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22296 23866 22324 25910
rect 22480 25786 22508 26318
rect 22388 25758 22508 25786
rect 22388 25702 22416 25758
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22572 25498 22600 29786
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22848 29170 22876 29242
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22664 27470 22692 27814
rect 22652 27464 22704 27470
rect 22704 27424 22784 27452
rect 22652 27406 22704 27412
rect 22756 26382 22784 27424
rect 22834 27296 22890 27305
rect 22834 27231 22890 27240
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22652 26240 22704 26246
rect 22652 26182 22704 26188
rect 22560 25492 22612 25498
rect 22480 25452 22560 25480
rect 22480 25294 22508 25452
rect 22560 25434 22612 25440
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22664 24585 22692 26182
rect 22756 25906 22784 26318
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22744 25696 22796 25702
rect 22744 25638 22796 25644
rect 22650 24576 22706 24585
rect 22650 24511 22706 24520
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 22388 23866 22416 24074
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21652 22166 21680 22646
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21088 22034 21140 22040
rect 21468 22066 21588 22094
rect 21468 21962 21496 22066
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21284 20058 21312 21490
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21100 19378 21128 19858
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20812 18148 20864 18154
rect 20916 18136 20944 18702
rect 20864 18108 20944 18136
rect 20812 18090 20864 18096
rect 20534 17776 20590 17785
rect 20534 17711 20590 17720
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16114 20484 16390
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15706 20392 15914
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20364 14618 20392 14826
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20350 14512 20406 14521
rect 20350 14447 20406 14456
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19890 13696 19946 13705
rect 20180 13682 20208 13942
rect 20180 13654 20300 13682
rect 19890 13631 19946 13640
rect 19904 13258 19932 13631
rect 20272 13326 20300 13654
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20088 12850 20116 12922
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19996 12617 20024 12650
rect 19982 12608 20038 12617
rect 19982 12543 20038 12552
rect 19892 12436 19944 12442
rect 19812 12406 19892 12434
rect 19708 12378 19760 12384
rect 19892 12378 19944 12384
rect 19614 11112 19670 11121
rect 19614 11047 19616 11056
rect 19668 11047 19670 11056
rect 19616 11018 19668 11024
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19352 8888 19380 9522
rect 19444 9042 19472 9998
rect 19720 9926 19748 12378
rect 19798 12336 19854 12345
rect 19798 12271 19854 12280
rect 19812 12102 19840 12271
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19904 11778 19932 12378
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 19996 12170 20024 12310
rect 20088 12306 20116 12786
rect 20260 12776 20312 12782
rect 20364 12764 20392 14447
rect 20456 14362 20484 15846
rect 20548 15026 20576 17070
rect 20640 16046 20668 17478
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 16726 20760 17138
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 16114 20760 16662
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20732 14929 20760 15098
rect 20718 14920 20774 14929
rect 20718 14855 20774 14864
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 14618 20668 14758
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20824 14385 20852 18090
rect 20902 17096 20958 17105
rect 20902 17031 20958 17040
rect 20916 16590 20944 17031
rect 20904 16584 20956 16590
rect 21008 16561 21036 19110
rect 21100 16998 21128 19314
rect 21192 19310 21220 19722
rect 21468 19446 21496 21898
rect 21546 21040 21602 21049
rect 21546 20975 21602 20984
rect 21560 20874 21588 20975
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21560 20534 21588 20810
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21456 19440 21508 19446
rect 21362 19408 21418 19417
rect 21456 19382 21508 19388
rect 21362 19343 21418 19352
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21192 18698 21220 18906
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21192 16658 21220 17138
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20904 16526 20956 16532
rect 20994 16552 21050 16561
rect 20994 16487 21050 16496
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20810 14376 20866 14385
rect 20456 14334 20576 14362
rect 20548 14090 20576 14334
rect 20720 14340 20772 14346
rect 20810 14311 20866 14320
rect 20720 14282 20772 14288
rect 20312 12736 20392 12764
rect 20456 14062 20576 14090
rect 20260 12718 20312 12724
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19800 11756 19852 11762
rect 19904 11750 20024 11778
rect 19800 11698 19852 11704
rect 19812 11370 19840 11698
rect 19996 11694 20024 11750
rect 19984 11688 20036 11694
rect 19890 11656 19946 11665
rect 19984 11630 20036 11636
rect 19890 11591 19892 11600
rect 19944 11591 19946 11600
rect 19892 11562 19944 11568
rect 19812 11342 19932 11370
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19812 10606 19840 11086
rect 19904 11014 19932 11342
rect 20088 11150 20116 12242
rect 20180 12102 20208 12650
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20168 11824 20220 11830
rect 20272 11801 20300 11834
rect 20168 11766 20220 11772
rect 20258 11792 20314 11801
rect 20180 11354 20208 11766
rect 20258 11727 20314 11736
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20364 11082 20392 11834
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19982 10840 20038 10849
rect 19982 10775 20038 10784
rect 19996 10742 20024 10775
rect 19984 10736 20036 10742
rect 19904 10696 19984 10724
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 9450 19748 9862
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19524 8900 19576 8906
rect 19352 8860 19524 8888
rect 19352 8498 19380 8860
rect 19524 8842 19576 8848
rect 19522 8528 19578 8537
rect 19340 8492 19392 8498
rect 19522 8463 19524 8472
rect 19340 8434 19392 8440
rect 19576 8463 19578 8472
rect 19524 8434 19576 8440
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18984 5710 19012 6394
rect 19062 6352 19118 6361
rect 19062 6287 19064 6296
rect 19116 6287 19118 6296
rect 19064 6258 19116 6264
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18786 3088 18842 3097
rect 18786 3023 18842 3032
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17408 1964 17460 1970
rect 17408 1906 17460 1912
rect 17684 1964 17736 1970
rect 17684 1906 17736 1912
rect 17224 1760 17276 1766
rect 17224 1702 17276 1708
rect 17040 1352 17092 1358
rect 17040 1294 17092 1300
rect 17236 1170 17264 1702
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 17328 1494 17356 1527
rect 17316 1488 17368 1494
rect 17316 1430 17368 1436
rect 17420 1358 17448 1906
rect 17868 1828 17920 1834
rect 17868 1770 17920 1776
rect 17880 1601 17908 1770
rect 17972 1766 18000 2858
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 17866 1592 17922 1601
rect 18156 1562 18184 2382
rect 18616 1970 18644 2382
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18315 1660 18623 1669
rect 18315 1658 18321 1660
rect 18377 1658 18401 1660
rect 18457 1658 18481 1660
rect 18537 1658 18561 1660
rect 18617 1658 18623 1660
rect 18377 1606 18379 1658
rect 18559 1606 18561 1658
rect 18315 1604 18321 1606
rect 18377 1604 18401 1606
rect 18457 1604 18481 1606
rect 18537 1604 18561 1606
rect 18617 1604 18623 1606
rect 18315 1595 18623 1604
rect 18708 1562 18736 2518
rect 18892 2446 18920 4558
rect 19168 2774 19196 6802
rect 19260 6322 19288 6802
rect 19352 6730 19380 8298
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19444 7818 19472 8230
rect 19536 8090 19564 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19628 7886 19656 9114
rect 19812 8362 19840 9590
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19904 7970 19932 10696
rect 19984 10678 20036 10684
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 10062 20024 10406
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19720 7942 19932 7970
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19616 7744 19668 7750
rect 19720 7732 19748 7942
rect 19892 7880 19944 7886
rect 19890 7848 19892 7857
rect 19984 7880 20036 7886
rect 19944 7848 19946 7857
rect 19984 7822 20036 7828
rect 19890 7783 19946 7792
rect 19668 7704 19748 7732
rect 19616 7686 19668 7692
rect 19628 7546 19656 7686
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19444 5710 19472 7346
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 5302 19380 5578
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 4622 19472 5646
rect 19536 5234 19564 6598
rect 19628 6390 19656 7278
rect 19904 6866 19932 7414
rect 19996 7410 20024 7822
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19982 7304 20038 7313
rect 19982 7239 19984 7248
rect 20036 7239 20038 7248
rect 19984 7210 20036 7216
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19996 6390 20024 6802
rect 19616 6384 19668 6390
rect 19616 6326 19668 6332
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 3738 19380 4490
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19536 3738 19564 3878
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19720 3652 19748 6190
rect 19800 5636 19852 5642
rect 19800 5578 19852 5584
rect 19812 5370 19840 5578
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19996 4060 20024 6326
rect 20088 5098 20116 9454
rect 20272 8906 20300 10542
rect 20364 10198 20392 11018
rect 20456 10810 20484 14062
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 13326 20576 13874
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20640 13394 20668 13806
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20732 13190 20760 14282
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12986 20760 13126
rect 20824 13002 20852 14214
rect 20916 13444 20944 15846
rect 21008 14958 21036 16390
rect 21086 16280 21142 16289
rect 21086 16215 21142 16224
rect 21100 15434 21128 16215
rect 21192 15706 21220 16458
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20996 13456 21048 13462
rect 20916 13416 20996 13444
rect 20996 13398 21048 13404
rect 21100 13258 21128 15370
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20720 12980 20772 12986
rect 20824 12974 20944 13002
rect 20720 12922 20772 12928
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20548 10674 20576 12038
rect 20640 10996 20668 12786
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12238 20760 12582
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20732 11150 20760 11766
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20640 10968 20760 10996
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20456 8906 20484 10202
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20640 9654 20668 9930
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20442 8664 20498 8673
rect 20442 8599 20498 8608
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20180 6798 20208 8298
rect 20456 7426 20484 8599
rect 20640 8498 20668 9318
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20732 8090 20760 10968
rect 20824 10674 20852 12854
rect 20916 12782 20944 12974
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12374 20944 12718
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20916 11082 20944 12106
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20824 10266 20852 10610
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21008 10198 21036 13194
rect 21100 11257 21128 13194
rect 21192 11626 21220 15302
rect 21284 14822 21312 19246
rect 21376 18766 21404 19343
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 15881 21404 18566
rect 21468 18358 21496 19382
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21560 17610 21588 19654
rect 21652 18970 21680 22102
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 22204 21690 22232 22578
rect 22296 21690 22324 23666
rect 22468 23248 22520 23254
rect 22468 23190 22520 23196
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22388 22438 22416 23122
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21744 21146 21772 21490
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 22112 20874 22140 21422
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22296 21026 22324 21354
rect 22480 21026 22508 23190
rect 22572 22778 22600 24074
rect 22756 23361 22784 25638
rect 22848 24206 22876 27231
rect 22928 26512 22980 26518
rect 22928 26454 22980 26460
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22742 23352 22798 23361
rect 22742 23287 22798 23296
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22848 23202 22876 23258
rect 22756 23174 22876 23202
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22572 22273 22600 22578
rect 22756 22574 22784 23174
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22558 22264 22614 22273
rect 22558 22199 22614 22208
rect 22756 22094 22784 22510
rect 22664 22066 22784 22094
rect 22664 22030 22692 22066
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22664 21486 22692 21966
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22848 21350 22876 22714
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22296 20998 22508 21026
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 21744 20330 21772 20470
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22204 19334 22232 19926
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 21928 19306 22232 19334
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 21928 18698 21956 19306
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 22112 18686 22232 18714
rect 22112 18630 22140 18686
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21362 15872 21418 15881
rect 21362 15807 21418 15816
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21376 14521 21404 15642
rect 21362 14512 21418 14521
rect 21362 14447 21418 14456
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10606 21128 11018
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 21008 9722 21036 10134
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21100 9586 21128 10134
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20548 7970 20576 8026
rect 20548 7942 20852 7970
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7546 20668 7754
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20456 7398 20668 7426
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20272 6322 20300 7142
rect 20548 7002 20576 7210
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20640 6934 20668 7398
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20732 7002 20760 7346
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20260 6316 20312 6322
rect 20640 6304 20668 6870
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 6322 20760 6598
rect 20260 6258 20312 6264
rect 20548 6276 20668 6304
rect 20720 6316 20772 6322
rect 20548 5574 20576 6276
rect 20720 6258 20772 6264
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20640 5846 20668 6122
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20180 5234 20208 5510
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 20076 4072 20128 4078
rect 19996 4032 20076 4060
rect 20076 4014 20128 4020
rect 19800 3664 19852 3670
rect 19720 3632 19800 3652
rect 19852 3632 19854 3641
rect 19720 3624 19798 3632
rect 19798 3567 19854 3576
rect 20088 3466 20116 4014
rect 20180 3738 20208 4558
rect 20456 4010 20484 5102
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20548 4826 20576 5034
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20456 3913 20484 3946
rect 20536 3936 20588 3942
rect 20442 3904 20498 3913
rect 20536 3878 20588 3884
rect 20442 3839 20498 3848
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19076 2746 19196 2774
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 17866 1527 17922 1536
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18696 1556 18748 1562
rect 18696 1498 18748 1504
rect 17408 1352 17460 1358
rect 17408 1294 17460 1300
rect 17592 1352 17644 1358
rect 17592 1294 17644 1300
rect 17604 1170 17632 1294
rect 17236 1142 17632 1170
rect 18880 1216 18932 1222
rect 18880 1158 18932 1164
rect 16764 740 16816 746
rect 16764 682 16816 688
rect 18892 610 18920 1158
rect 19076 610 19104 2746
rect 19430 2680 19486 2689
rect 19430 2615 19486 2624
rect 19444 2582 19472 2615
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19628 2446 19656 3334
rect 20180 2446 20208 3674
rect 20442 3496 20498 3505
rect 20442 3431 20498 3440
rect 20456 3194 20484 3431
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20272 2922 20300 3130
rect 20548 3058 20576 3878
rect 20640 3670 20668 5646
rect 20732 5234 20760 6258
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4214 20760 4966
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20824 3670 20852 7942
rect 20916 7546 20944 8774
rect 21100 8294 21128 9522
rect 21192 8294 21220 11086
rect 21284 11082 21312 13874
rect 21468 12306 21496 17478
rect 21560 16425 21588 17546
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 21928 16522 21956 17070
rect 22020 16522 22048 17138
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 21546 16416 21602 16425
rect 21546 16351 21602 16360
rect 21546 15872 21602 15881
rect 21546 15807 21602 15816
rect 21560 15502 21588 15807
rect 21652 15502 21680 16458
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21836 15638 21864 15846
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21560 15366 21588 15438
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21560 15026 21588 15302
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21560 14414 21588 14962
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 13938 21588 14350
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21652 13802 21680 15030
rect 22204 14362 22232 18686
rect 22296 17338 22324 19790
rect 22388 19514 22416 20878
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22480 19394 22508 20998
rect 22940 20913 22968 26454
rect 23032 25974 23060 29990
rect 23216 27062 23244 30330
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 23492 28966 23520 30262
rect 23676 30258 23704 31282
rect 23952 30938 23980 31690
rect 24964 31346 24992 33390
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24596 30258 24624 30670
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 23676 29646 23704 30194
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 23676 29102 23704 29582
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23754 29064 23810 29073
rect 23754 28999 23810 29008
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23664 28960 23716 28966
rect 23664 28902 23716 28908
rect 23676 28558 23704 28902
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23400 26518 23428 26726
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23112 26376 23164 26382
rect 23296 26376 23348 26382
rect 23112 26318 23164 26324
rect 23202 26344 23258 26353
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23032 23662 23060 24754
rect 23124 24313 23152 26318
rect 23296 26318 23348 26324
rect 23202 26279 23204 26288
rect 23256 26279 23258 26288
rect 23204 26250 23256 26256
rect 23204 25968 23256 25974
rect 23204 25910 23256 25916
rect 23216 25498 23244 25910
rect 23308 25537 23336 26318
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23294 25528 23350 25537
rect 23204 25492 23256 25498
rect 23294 25463 23350 25472
rect 23204 25434 23256 25440
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23400 24721 23428 24890
rect 23386 24712 23442 24721
rect 23492 24682 23520 25842
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23386 24647 23442 24656
rect 23480 24676 23532 24682
rect 23480 24618 23532 24624
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23110 24304 23166 24313
rect 23110 24239 23166 24248
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23020 23656 23072 23662
rect 23020 23598 23072 23604
rect 23018 23352 23074 23361
rect 23018 23287 23074 23296
rect 23032 23118 23060 23287
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23124 22778 23152 24006
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23216 21593 23244 24074
rect 23308 23730 23336 24142
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23308 23322 23336 23666
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 23308 21672 23336 22986
rect 23400 22438 23428 24550
rect 23584 23798 23612 25162
rect 23676 25158 23704 28494
rect 23768 26790 23796 28999
rect 23860 28762 23888 29582
rect 24492 29572 24544 29578
rect 24492 29514 24544 29520
rect 23848 28756 23900 28762
rect 23848 28698 23900 28704
rect 24032 27872 24084 27878
rect 24124 27872 24176 27878
rect 24032 27814 24084 27820
rect 24122 27840 24124 27849
rect 24176 27840 24178 27849
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23940 26784 23992 26790
rect 23940 26726 23992 26732
rect 23848 26308 23900 26314
rect 23848 26250 23900 26256
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23860 24857 23888 26250
rect 23846 24848 23902 24857
rect 23846 24783 23902 24792
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23664 24336 23716 24342
rect 23664 24278 23716 24284
rect 23572 23792 23624 23798
rect 23572 23734 23624 23740
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23308 21644 23428 21672
rect 23202 21584 23258 21593
rect 23202 21519 23258 21528
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21078 23152 21286
rect 23308 21146 23336 21490
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 22926 20904 22982 20913
rect 22926 20839 22982 20848
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22388 19366 22508 19394
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22388 17270 22416 19366
rect 22572 18698 22600 19654
rect 22756 19514 22784 20402
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22848 18766 22876 20198
rect 23032 19446 23060 20810
rect 23124 19825 23152 21014
rect 23110 19816 23166 19825
rect 23110 19751 23166 19760
rect 23400 19514 23428 21644
rect 23492 21418 23520 23666
rect 23676 23633 23704 24278
rect 23662 23624 23718 23633
rect 23662 23559 23718 23568
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23480 21412 23532 21418
rect 23480 21354 23532 21360
rect 23584 21078 23612 22646
rect 23768 21894 23796 24686
rect 23952 24138 23980 26726
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23584 19922 23612 20198
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 23296 19236 23348 19242
rect 23296 19178 23348 19184
rect 23572 19236 23624 19242
rect 23572 19178 23624 19184
rect 23308 18902 23336 19178
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22480 18154 22784 18170
rect 22468 18148 22784 18154
rect 22520 18142 22784 18148
rect 22468 18090 22520 18096
rect 22756 18086 22784 18142
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22572 17814 22600 18022
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22480 17066 22508 17614
rect 22560 17604 22612 17610
rect 22560 17546 22612 17552
rect 22572 17270 22600 17546
rect 22848 17542 22876 18702
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23032 17610 23060 17750
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22848 17134 22876 17478
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22296 16250 22324 16662
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22388 16182 22416 17002
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22388 14521 22416 14962
rect 22374 14512 22430 14521
rect 22374 14447 22430 14456
rect 22204 14334 22416 14362
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22204 13977 22232 14010
rect 22190 13968 22246 13977
rect 22190 13903 22246 13912
rect 22100 13864 22152 13870
rect 22098 13832 22100 13841
rect 22152 13832 22154 13841
rect 21640 13796 21692 13802
rect 22098 13767 22154 13776
rect 21640 13738 21692 13744
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21560 12374 21588 13466
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21376 10130 21404 12106
rect 21560 11830 21588 12310
rect 21652 11898 21680 13738
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22296 12850 22324 14214
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22388 12730 22416 14334
rect 22480 14006 22508 14962
rect 22572 14346 22600 15982
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22480 12850 22508 13942
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 12918 22600 13670
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22388 12702 22508 12730
rect 22480 12646 22508 12702
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22112 12209 22140 12378
rect 22284 12232 22336 12238
rect 22098 12200 22154 12209
rect 22284 12174 22336 12180
rect 22098 12135 22154 12144
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21376 9382 21404 10066
rect 21468 9654 21496 11018
rect 21560 10198 21588 11562
rect 22020 11286 22048 11630
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21652 10146 21680 11222
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 21732 10192 21784 10198
rect 21652 10140 21732 10146
rect 21652 10134 21784 10140
rect 22112 10146 22140 10542
rect 21652 10118 21772 10134
rect 21824 10124 21876 10130
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21284 8974 21312 9318
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21376 7936 21404 9318
rect 21560 8974 21588 9862
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 8090 21588 8230
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21548 7948 21600 7954
rect 21376 7908 21548 7936
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21376 6390 21404 7908
rect 21548 7890 21600 7896
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 7274 21588 7686
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21652 6730 21680 10118
rect 22112 10118 22232 10146
rect 21824 10066 21876 10072
rect 21836 9994 21864 10066
rect 22204 10062 22232 10118
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 22112 9908 22140 9998
rect 22112 9880 22232 9908
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 8945 22048 9386
rect 22006 8936 22062 8945
rect 22006 8871 22062 8880
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 21928 8537 21956 8570
rect 22112 8537 22140 8570
rect 21914 8528 21970 8537
rect 21914 8463 21970 8472
rect 22098 8528 22154 8537
rect 22204 8514 22232 9880
rect 22296 9586 22324 12174
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22388 9042 22416 12582
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22480 11558 22508 12106
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 10062 22508 11494
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22572 10810 22600 11222
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22664 10674 22692 16050
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22756 13734 22784 15506
rect 23124 15065 23152 17138
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 16182 23336 16458
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23110 15056 23166 15065
rect 23110 14991 23166 15000
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22848 13802 22876 14486
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22756 13326 22784 13398
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22756 11665 22784 13262
rect 22940 12374 22968 14350
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23124 13870 23152 14282
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23124 13530 23152 13806
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23124 13258 23152 13466
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23124 12434 23152 13194
rect 23032 12406 23152 12434
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22926 12200 22982 12209
rect 23032 12170 23060 12406
rect 23216 12186 23244 15370
rect 23308 15026 23336 15846
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23400 14550 23428 16526
rect 23492 16454 23520 18702
rect 23584 18630 23612 19178
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23676 18426 23704 18566
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23768 18290 23796 19382
rect 23860 19174 23888 21830
rect 23952 21622 23980 23462
rect 24044 22982 24072 27814
rect 24122 27775 24178 27784
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 25498 24164 27270
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24124 25492 24176 25498
rect 24124 25434 24176 25440
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 24136 23361 24164 23462
rect 24122 23352 24178 23361
rect 24122 23287 24178 23296
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 24044 19938 24072 21558
rect 23952 19910 24072 19938
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23676 17762 23704 18158
rect 23584 17734 23704 17762
rect 23584 17542 23612 17734
rect 23768 17626 23796 18226
rect 23952 18154 23980 19910
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23676 17598 23796 17626
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23676 16266 23704 17598
rect 23860 16726 23888 17818
rect 23952 17746 23980 18090
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23848 16720 23900 16726
rect 23848 16662 23900 16668
rect 24044 16454 24072 19790
rect 24136 18290 24164 22034
rect 24228 20602 24256 23666
rect 24320 23089 24348 26930
rect 24504 24614 24532 29514
rect 24596 28558 24624 29582
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24688 28218 24716 31282
rect 24858 30968 24914 30977
rect 25148 30938 25176 32438
rect 25261 32124 25569 32133
rect 25261 32122 25267 32124
rect 25323 32122 25347 32124
rect 25403 32122 25427 32124
rect 25483 32122 25507 32124
rect 25563 32122 25569 32124
rect 25323 32070 25325 32122
rect 25505 32070 25507 32122
rect 25261 32068 25267 32070
rect 25323 32068 25347 32070
rect 25403 32068 25427 32070
rect 25483 32068 25507 32070
rect 25563 32068 25569 32070
rect 25261 32059 25569 32068
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 24858 30903 24914 30912
rect 25136 30932 25188 30938
rect 24872 30433 24900 30903
rect 25136 30874 25188 30880
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24858 30424 24914 30433
rect 24858 30359 24914 30368
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24766 28656 24822 28665
rect 24766 28591 24822 28600
rect 24780 28218 24808 28591
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24872 28082 24900 30194
rect 24964 29306 24992 30670
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 25608 29034 25636 33458
rect 27344 33312 27396 33318
rect 27344 33254 27396 33260
rect 26792 33176 26844 33182
rect 26792 33118 26844 33124
rect 26424 32836 26476 32842
rect 26424 32778 26476 32784
rect 25780 32768 25832 32774
rect 25780 32710 25832 32716
rect 25792 31210 25820 32710
rect 25872 32564 25924 32570
rect 25872 32506 25924 32512
rect 25884 31958 25912 32506
rect 25964 32428 26016 32434
rect 25964 32370 26016 32376
rect 25872 31952 25924 31958
rect 25872 31894 25924 31900
rect 25976 31346 26004 32370
rect 26436 31958 26464 32778
rect 26424 31952 26476 31958
rect 26424 31894 26476 31900
rect 26516 31952 26568 31958
rect 26516 31894 26568 31900
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26424 31816 26476 31822
rect 26424 31758 26476 31764
rect 25964 31340 26016 31346
rect 25964 31282 26016 31288
rect 25780 31204 25832 31210
rect 25780 31146 25832 31152
rect 25976 30802 26004 31282
rect 26240 31272 26292 31278
rect 26146 31240 26202 31249
rect 26240 31214 26292 31220
rect 26146 31175 26202 31184
rect 25964 30796 26016 30802
rect 25964 30738 26016 30744
rect 25870 30424 25926 30433
rect 25870 30359 25926 30368
rect 25884 29322 25912 30359
rect 25976 30258 26004 30738
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 25884 29294 26004 29322
rect 25872 29232 25924 29238
rect 25870 29200 25872 29209
rect 25924 29200 25926 29209
rect 25780 29164 25832 29170
rect 25870 29135 25926 29144
rect 25780 29106 25832 29112
rect 25792 29073 25820 29106
rect 25778 29064 25834 29073
rect 24952 29028 25004 29034
rect 24952 28970 25004 28976
rect 25596 29028 25648 29034
rect 25778 28999 25834 29008
rect 25596 28970 25648 28976
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24964 27713 24992 28970
rect 25688 28960 25740 28966
rect 25134 28928 25190 28937
rect 25688 28902 25740 28908
rect 25134 28863 25190 28872
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24950 27704 25006 27713
rect 24950 27639 25006 27648
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24688 26450 24716 27406
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24584 25696 24636 25702
rect 24688 25684 24716 26386
rect 24636 25656 24716 25684
rect 24584 25638 24636 25644
rect 24780 25430 24808 26930
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24596 24886 24624 25230
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24688 23769 24716 25094
rect 24872 24682 24900 26250
rect 24964 25974 24992 26862
rect 25056 26761 25084 28358
rect 25148 28218 25176 28863
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 25516 28626 25636 28642
rect 25516 28620 25648 28626
rect 25516 28614 25596 28620
rect 25136 28212 25188 28218
rect 25136 28154 25188 28160
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25148 27418 25176 28018
rect 25516 27962 25544 28614
rect 25596 28562 25648 28568
rect 25594 28520 25650 28529
rect 25594 28455 25650 28464
rect 25608 28082 25636 28455
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25516 27934 25636 27962
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25148 27390 25268 27418
rect 25136 27328 25188 27334
rect 25134 27296 25136 27305
rect 25188 27296 25190 27305
rect 25134 27231 25190 27240
rect 25240 26874 25268 27390
rect 25148 26846 25268 26874
rect 25042 26752 25098 26761
rect 25042 26687 25098 26696
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 24952 25968 25004 25974
rect 24952 25910 25004 25916
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24964 24410 24992 25638
rect 25056 24886 25084 25978
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25148 24290 25176 26846
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25608 25974 25636 27934
rect 25700 26489 25728 28902
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25976 28506 26004 29294
rect 26068 28762 26096 30194
rect 26160 29850 26188 31175
rect 26252 30938 26280 31214
rect 26240 30932 26292 30938
rect 26240 30874 26292 30880
rect 26240 30320 26292 30326
rect 26238 30288 26240 30297
rect 26292 30288 26294 30297
rect 26238 30223 26294 30232
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26252 28914 26280 29038
rect 26160 28886 26280 28914
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 25686 26480 25742 26489
rect 25686 26415 25742 26424
rect 25596 25968 25648 25974
rect 25596 25910 25648 25916
rect 25686 25936 25742 25945
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25608 24886 25636 25910
rect 25686 25871 25688 25880
rect 25740 25871 25742 25880
rect 25688 25842 25740 25848
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25056 24262 25176 24290
rect 25056 24177 25084 24262
rect 25136 24200 25188 24206
rect 25042 24168 25098 24177
rect 24860 24132 24912 24138
rect 25136 24142 25188 24148
rect 25042 24103 25098 24112
rect 24860 24074 24912 24080
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24674 23760 24730 23769
rect 24674 23695 24730 23704
rect 24492 23520 24544 23526
rect 24492 23462 24544 23468
rect 24306 23080 24362 23089
rect 24306 23015 24362 23024
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24320 20369 24348 22374
rect 24412 21010 24440 22986
rect 24400 21004 24452 21010
rect 24504 20992 24532 23462
rect 24582 23216 24638 23225
rect 24582 23151 24638 23160
rect 24596 22642 24624 23151
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24674 22536 24730 22545
rect 24674 22471 24676 22480
rect 24728 22471 24730 22480
rect 24676 22442 24728 22448
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24584 21004 24636 21010
rect 24504 20964 24584 20992
rect 24400 20946 24452 20952
rect 24584 20946 24636 20952
rect 24596 20466 24624 20946
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24306 20360 24362 20369
rect 24306 20295 24362 20304
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 23492 16238 23704 16266
rect 23492 15366 23520 16238
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23492 12714 23520 14962
rect 23584 14550 23612 15914
rect 23676 14890 23704 15914
rect 24044 15502 24072 15982
rect 24136 15978 24164 16390
rect 24124 15972 24176 15978
rect 24124 15914 24176 15920
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23940 14952 23992 14958
rect 24044 14940 24072 15438
rect 23992 14912 24072 14940
rect 23940 14894 23992 14900
rect 23664 14884 23716 14890
rect 23664 14826 23716 14832
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23768 14278 23796 14758
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23584 14074 23612 14214
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23584 12850 23612 13670
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23296 12640 23348 12646
rect 23294 12608 23296 12617
rect 23348 12608 23350 12617
rect 23294 12543 23350 12552
rect 22926 12135 22982 12144
rect 23020 12164 23072 12170
rect 22742 11656 22798 11665
rect 22742 11591 22798 11600
rect 22940 10674 22968 12135
rect 23020 12106 23072 12112
rect 23124 12158 23244 12186
rect 23124 11626 23152 12158
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23216 11762 23244 12038
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22572 8922 22600 10474
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22848 9761 22876 10066
rect 22834 9752 22890 9761
rect 22834 9687 22890 9696
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22388 8906 22600 8922
rect 22376 8900 22600 8906
rect 22428 8894 22600 8900
rect 22376 8842 22428 8848
rect 22388 8809 22416 8842
rect 22468 8832 22520 8838
rect 22374 8800 22430 8809
rect 22468 8774 22520 8780
rect 22374 8735 22430 8744
rect 22204 8486 22416 8514
rect 22098 8463 22154 8472
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22296 7546 22324 8366
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 21744 6866 21772 7482
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 21364 6384 21416 6390
rect 22100 6384 22152 6390
rect 21364 6326 21416 6332
rect 22020 6332 22100 6338
rect 22020 6326 22152 6332
rect 22020 6310 22140 6326
rect 22204 6322 22232 7346
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22192 6316 22244 6322
rect 22020 6254 22048 6310
rect 22192 6258 22244 6264
rect 21088 6248 21140 6254
rect 20994 6216 21050 6225
rect 21088 6190 21140 6196
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 20994 6151 20996 6160
rect 21048 6151 21050 6160
rect 20996 6122 21048 6128
rect 21008 5030 21036 6122
rect 21100 5846 21128 6190
rect 21284 5914 21312 6190
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 21652 4690 21680 5170
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19720 2258 19748 2382
rect 20456 2310 20484 2450
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 19444 2230 19748 2258
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 19444 1358 19472 2230
rect 20548 1986 20576 2382
rect 20548 1958 20668 1986
rect 20916 1970 20944 3062
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21192 2145 21220 2586
rect 21284 2378 21312 4422
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21560 3466 21588 4082
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 21178 2136 21234 2145
rect 21178 2071 21234 2080
rect 21376 1970 21404 3334
rect 20640 1902 20668 1958
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 21364 1964 21416 1970
rect 21364 1906 21416 1912
rect 20628 1896 20680 1902
rect 20628 1838 20680 1844
rect 21468 1358 21496 3334
rect 21560 3126 21588 3402
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 21652 2582 21680 4218
rect 22204 4146 22232 5578
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22296 4010 22324 7278
rect 22388 5930 22416 8486
rect 22480 7954 22508 8774
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22572 7342 22600 7822
rect 22664 7410 22692 9590
rect 22756 9382 22784 9590
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22848 9178 22876 9522
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22940 9058 22968 10610
rect 23216 10198 23244 11086
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23308 10130 23336 12543
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23400 10962 23428 12310
rect 23492 12238 23520 12378
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23400 10934 23520 10962
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23492 9466 23520 10934
rect 23584 9586 23612 12242
rect 23676 11694 23704 12786
rect 23768 12374 23796 14214
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23952 13394 23980 13466
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 24044 13326 24072 14912
rect 24228 14074 24256 19722
rect 24688 19417 24716 21830
rect 24780 20534 24808 23802
rect 24872 23322 24900 24074
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 25148 22642 25176 24142
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24872 22234 24900 22510
rect 25148 22234 25176 22578
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25148 22094 25176 22170
rect 24964 22066 25176 22094
rect 24964 22030 24992 22066
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 25056 21350 25084 21558
rect 25608 21418 25636 24006
rect 25700 23225 25728 25434
rect 25686 23216 25742 23225
rect 25686 23151 25742 23160
rect 25792 22982 25820 28494
rect 25872 28484 25924 28490
rect 25976 28478 26096 28506
rect 25872 28426 25924 28432
rect 25884 26994 25912 28426
rect 26068 28218 26096 28478
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26068 27033 26096 28018
rect 26054 27024 26110 27033
rect 25872 26988 25924 26994
rect 26054 26959 26110 26968
rect 25872 26930 25924 26936
rect 26160 26897 26188 28886
rect 26240 28688 26292 28694
rect 26240 28630 26292 28636
rect 26252 27674 26280 28630
rect 26344 28218 26372 31758
rect 26436 30784 26464 31758
rect 26528 31142 26556 31894
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26620 31090 26648 31758
rect 26804 31346 26832 33118
rect 27356 31822 27384 33254
rect 27896 33244 27948 33250
rect 27896 33186 27948 33192
rect 27712 32972 27764 32978
rect 27712 32914 27764 32920
rect 27724 31958 27752 32914
rect 27712 31952 27764 31958
rect 27712 31894 27764 31900
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 27066 31376 27122 31385
rect 26792 31340 26844 31346
rect 27066 31311 27122 31320
rect 26792 31282 26844 31288
rect 26792 31136 26844 31142
rect 26620 31062 26740 31090
rect 26792 31078 26844 31084
rect 26436 30756 26556 30784
rect 26422 30696 26478 30705
rect 26422 30631 26478 30640
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 26436 28082 26464 30631
rect 26528 29782 26556 30756
rect 26516 29776 26568 29782
rect 26516 29718 26568 29724
rect 26608 29640 26660 29646
rect 26608 29582 26660 29588
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26528 27985 26556 29106
rect 26514 27976 26570 27985
rect 26514 27911 26570 27920
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26146 26888 26202 26897
rect 26146 26823 26202 26832
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25870 25800 25926 25809
rect 25870 25735 25872 25744
rect 25924 25735 25926 25744
rect 25872 25706 25924 25712
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 20942 25176 21286
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25884 21049 25912 24550
rect 25976 22642 26004 26726
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26056 25288 26108 25294
rect 26056 25230 26108 25236
rect 26068 24274 26096 25230
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 26160 23526 26188 26318
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 23118 26188 23462
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 26252 21690 26280 24074
rect 26436 22982 26464 25162
rect 26528 24206 26556 26182
rect 26620 24954 26648 29582
rect 26712 29238 26740 31062
rect 26804 30190 26832 31078
rect 27080 30802 27108 31311
rect 27804 30864 27856 30870
rect 27802 30832 27804 30841
rect 27856 30832 27858 30841
rect 27068 30796 27120 30802
rect 27802 30767 27858 30776
rect 27068 30738 27120 30744
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 26792 30184 26844 30190
rect 26792 30126 26844 30132
rect 26700 29232 26752 29238
rect 26700 29174 26752 29180
rect 27080 29170 27108 30194
rect 27618 30152 27674 30161
rect 27618 30087 27674 30096
rect 27632 29646 27660 30087
rect 27804 30048 27856 30054
rect 27804 29990 27856 29996
rect 27816 29753 27844 29990
rect 27802 29744 27858 29753
rect 27802 29679 27858 29688
rect 27620 29640 27672 29646
rect 27158 29608 27214 29617
rect 27620 29582 27672 29588
rect 27158 29543 27214 29552
rect 27172 29306 27200 29543
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27908 29170 27936 33186
rect 28734 32668 29042 32677
rect 28734 32666 28740 32668
rect 28796 32666 28820 32668
rect 28876 32666 28900 32668
rect 28956 32666 28980 32668
rect 29036 32666 29042 32668
rect 28796 32614 28798 32666
rect 28978 32614 28980 32666
rect 28734 32612 28740 32614
rect 28796 32612 28820 32614
rect 28876 32612 28900 32614
rect 28956 32612 28980 32614
rect 29036 32612 29042 32614
rect 28734 32603 29042 32612
rect 28080 32292 28132 32298
rect 28080 32234 28132 32240
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 28000 32026 28028 32166
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 27988 30252 28040 30258
rect 27988 30194 28040 30200
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27896 29164 27948 29170
rect 27896 29106 27948 29112
rect 27618 28112 27674 28121
rect 27618 28047 27620 28056
rect 27672 28047 27674 28056
rect 27620 28018 27672 28024
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 25498 27660 27270
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 28000 25401 28028 30194
rect 28092 26994 28120 32234
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 28356 26240 28408 26246
rect 28356 26182 28408 26188
rect 27986 25392 28042 25401
rect 27986 25327 28042 25336
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26516 23044 26568 23050
rect 26516 22986 26568 22992
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 25870 21040 25926 21049
rect 25870 20975 25926 20984
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24768 20528 24820 20534
rect 24768 20470 24820 20476
rect 24964 20058 24992 20810
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 24674 19408 24730 19417
rect 24308 19372 24360 19378
rect 24674 19343 24730 19352
rect 24308 19314 24360 19320
rect 24320 17814 24348 19314
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 24952 18964 25004 18970
rect 25056 18952 25084 19110
rect 25004 18924 25084 18952
rect 24952 18906 25004 18912
rect 25148 18834 25176 20402
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 24412 18222 24440 18770
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 24320 14929 24348 17546
rect 25056 17202 25084 18022
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24596 16969 24624 17002
rect 24582 16960 24638 16969
rect 24582 16895 24638 16904
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25700 16794 25728 20538
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24596 15502 24624 16594
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24872 15162 24900 16458
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25608 15706 25636 16050
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24306 14920 24362 14929
rect 24306 14855 24362 14864
rect 24964 14414 24992 15642
rect 25792 15502 25820 18022
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25884 15094 25912 20742
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26068 16522 26096 19654
rect 26252 18426 26280 20402
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26344 17882 26372 20742
rect 26528 20482 26556 22986
rect 26620 22137 26648 23462
rect 26606 22128 26662 22137
rect 26606 22063 26662 22072
rect 27448 22001 27476 25094
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27434 21992 27490 22001
rect 27434 21927 27490 21936
rect 27816 21146 27844 24006
rect 28368 23866 28396 26182
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26436 20454 26556 20482
rect 26436 19990 26464 20454
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26424 19984 26476 19990
rect 26424 19926 26476 19932
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26528 17678 26556 20198
rect 26804 19922 26832 20878
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26804 19446 26832 19858
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26804 17882 26832 19382
rect 28184 19242 28212 21830
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28172 19236 28224 19242
rect 28172 19178 28224 19184
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17338 26188 17478
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26252 16250 26280 17138
rect 26804 16998 26832 17818
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 26804 16794 26832 16934
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25976 14890 26004 15574
rect 27080 15502 27108 16934
rect 27448 16250 27476 18158
rect 27804 17808 27856 17814
rect 27802 17776 27804 17785
rect 27856 17776 27858 17785
rect 27802 17711 27858 17720
rect 28368 17542 28396 19654
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27528 16992 27580 16998
rect 27528 16934 27580 16940
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27540 16114 27568 16934
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27632 15994 27660 17070
rect 27804 17060 27856 17066
rect 27804 17002 27856 17008
rect 27540 15966 27660 15994
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 25964 14884 26016 14890
rect 25964 14826 26016 14832
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25976 14618 26004 14826
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 26332 14408 26384 14414
rect 26436 14396 26464 15438
rect 27540 15366 27568 15966
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 14958 27568 15302
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 26384 14368 26464 14396
rect 26332 14350 26384 14356
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24504 14074 24532 14214
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 25504 14000 25556 14006
rect 25502 13968 25504 13977
rect 25556 13968 25558 13977
rect 24216 13932 24268 13938
rect 25502 13903 25558 13912
rect 24216 13874 24268 13880
rect 24228 13530 24256 13874
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 24964 13530 24992 13806
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 23848 13252 23900 13258
rect 23848 13194 23900 13200
rect 23860 12442 23888 13194
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23756 12368 23808 12374
rect 23756 12310 23808 12316
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23676 10810 23704 11630
rect 24044 11354 24072 12922
rect 24596 12918 24624 13262
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24398 12744 24454 12753
rect 24398 12679 24454 12688
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23676 10606 23704 10746
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23676 9586 23704 10542
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23492 9438 23796 9466
rect 23768 9382 23796 9438
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 22848 9030 22968 9058
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22756 7546 22784 8842
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22848 6390 22876 9030
rect 23112 8900 23164 8906
rect 23112 8842 23164 8848
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23124 8430 23152 8842
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 22926 7984 22982 7993
rect 22926 7919 22982 7928
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22388 5902 22784 5930
rect 22756 5846 22784 5902
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22940 5778 22968 7919
rect 23124 7002 23152 8026
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23216 7410 23244 7686
rect 23492 7478 23520 8230
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23584 7274 23612 8842
rect 23860 7886 23888 10406
rect 24044 10198 24072 11290
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23952 7886 23980 9862
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24044 9178 24072 9658
rect 24412 9450 24440 12679
rect 24688 12238 24716 13126
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24872 11898 24900 13466
rect 25056 12442 25084 13670
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 25148 12209 25176 13806
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25332 12753 25360 12786
rect 25318 12744 25374 12753
rect 26160 12730 26188 13466
rect 26436 13326 26464 14368
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 13326 26740 14214
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 27172 13530 27200 13806
rect 27448 13802 27476 14758
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26436 12918 26464 13262
rect 27172 12918 27200 13466
rect 26424 12912 26476 12918
rect 26424 12854 26476 12860
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 26160 12714 26280 12730
rect 26160 12708 26292 12714
rect 26160 12702 26240 12708
rect 25318 12679 25374 12688
rect 26240 12650 26292 12656
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 26436 12306 26464 12854
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24688 11082 24716 11562
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 25042 11112 25098 11121
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24872 10690 24900 11086
rect 25148 11082 25176 11494
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 26252 11354 26280 11766
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 25042 11047 25098 11056
rect 25136 11076 25188 11082
rect 25056 10810 25084 11047
rect 25136 11018 25188 11024
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 24872 10662 25176 10690
rect 26344 10674 26372 12242
rect 26712 11762 26740 12582
rect 27540 11830 27568 14894
rect 27724 13841 27752 15846
rect 27816 15094 27844 17002
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28080 15428 28132 15434
rect 28080 15370 28132 15376
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 28092 14074 28120 15370
rect 28184 15162 28212 16050
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 27710 13832 27766 13841
rect 27710 13767 27766 13776
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27632 12850 27660 13670
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27528 11824 27580 11830
rect 26974 11792 27030 11801
rect 26700 11756 26752 11762
rect 27528 11766 27580 11772
rect 26974 11727 27030 11736
rect 26700 11698 26752 11704
rect 26988 11150 27016 11727
rect 27724 11626 27752 13767
rect 28080 13252 28132 13258
rect 28080 13194 28132 13200
rect 28092 12986 28120 13194
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 27712 11620 27764 11626
rect 27712 11562 27764 11568
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 25148 10062 25176 10662
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24492 9716 24544 9722
rect 24492 9658 24544 9664
rect 24504 9586 24532 9658
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24766 9480 24822 9489
rect 24400 9444 24452 9450
rect 24766 9415 24822 9424
rect 24400 9386 24452 9392
rect 24780 9178 24808 9415
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24688 8430 24716 8910
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23768 6798 23796 7278
rect 24030 6896 24086 6905
rect 24030 6831 24086 6840
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23388 6384 23440 6390
rect 23386 6352 23388 6361
rect 23440 6352 23442 6361
rect 23204 6316 23256 6322
rect 23386 6287 23442 6296
rect 23204 6258 23256 6264
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22756 5234 22784 5646
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22388 4185 22416 4694
rect 22374 4176 22430 4185
rect 22374 4111 22430 4120
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22296 3890 22324 3946
rect 22560 3936 22612 3942
rect 22296 3862 22416 3890
rect 22560 3878 22612 3884
rect 21914 3496 21970 3505
rect 21914 3431 21916 3440
rect 21968 3431 21970 3440
rect 21916 3402 21968 3408
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21744 2922 21772 3130
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21928 2689 21956 2994
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 21914 2680 21970 2689
rect 21914 2615 21970 2624
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 22020 2530 22048 2926
rect 22296 2854 22324 3334
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22020 2514 22140 2530
rect 22020 2508 22152 2514
rect 22020 2502 22100 2508
rect 22100 2450 22152 2456
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 21546 2136 21602 2145
rect 21546 2071 21602 2080
rect 21560 1970 21588 2071
rect 21548 1964 21600 1970
rect 21548 1906 21600 1912
rect 21652 1834 21680 2382
rect 22388 2310 22416 3862
rect 22572 3602 22600 3878
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22664 3534 22692 4082
rect 22756 4010 22784 5170
rect 23216 4622 23244 6258
rect 23388 6112 23440 6118
rect 23572 6112 23624 6118
rect 23440 6060 23520 6066
rect 23388 6054 23520 6060
rect 23572 6054 23624 6060
rect 23400 6038 23520 6054
rect 23492 5914 23520 6038
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23584 5794 23612 6054
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23400 5766 23612 5794
rect 23400 5710 23428 5766
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23388 4208 23440 4214
rect 23386 4176 23388 4185
rect 23440 4176 23442 4185
rect 23204 4140 23256 4146
rect 23492 4146 23520 4558
rect 23386 4111 23442 4120
rect 23480 4140 23532 4146
rect 23204 4082 23256 4088
rect 23480 4082 23532 4088
rect 22836 4072 22888 4078
rect 22888 4020 23060 4026
rect 22836 4014 23060 4020
rect 22744 4004 22796 4010
rect 22848 3998 23060 4014
rect 22744 3946 22796 3952
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22756 3346 22784 3946
rect 23032 3466 23060 3998
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 22572 3318 22784 3346
rect 22572 2514 22600 3318
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 22376 2304 22428 2310
rect 22376 2246 22428 2252
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 22572 2038 22600 2450
rect 22560 2032 22612 2038
rect 22560 1974 22612 1980
rect 21640 1828 21692 1834
rect 21640 1770 21692 1776
rect 22572 1358 22600 1974
rect 22664 1766 22692 2790
rect 22652 1760 22704 1766
rect 22652 1702 22704 1708
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 21456 1352 21508 1358
rect 21456 1294 21508 1300
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 23216 1290 23244 4082
rect 23952 4078 23980 5850
rect 24044 5370 24072 6831
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24228 6186 24256 6258
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24504 5914 24532 7754
rect 24688 7410 24716 8366
rect 24872 8090 24900 9930
rect 25148 9722 25176 9998
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25226 8936 25282 8945
rect 25226 8871 25282 8880
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24688 6798 24716 7346
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6254 24716 6734
rect 24964 6730 24992 8774
rect 25240 8566 25268 8871
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25148 6916 25176 7890
rect 25686 7304 25742 7313
rect 25686 7239 25742 7248
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25148 6888 25268 6916
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24688 5794 24716 6190
rect 24596 5766 24716 5794
rect 24596 5710 24624 5766
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24780 5658 24808 6598
rect 25148 6458 25176 6666
rect 25240 6458 25268 6888
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 24780 5642 24900 5658
rect 24216 5636 24268 5642
rect 24780 5636 24912 5642
rect 24780 5630 24860 5636
rect 24216 5578 24268 5584
rect 24860 5578 24912 5584
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24122 5128 24178 5137
rect 24122 5063 24178 5072
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23386 3904 23442 3913
rect 23386 3839 23442 3848
rect 23400 2922 23428 3839
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23400 1834 23428 2382
rect 23848 2032 23900 2038
rect 23848 1974 23900 1980
rect 23860 1902 23888 1974
rect 23848 1896 23900 1902
rect 23848 1838 23900 1844
rect 23388 1828 23440 1834
rect 23388 1770 23440 1776
rect 23480 1760 23532 1766
rect 23480 1702 23532 1708
rect 23492 1562 23520 1702
rect 23480 1556 23532 1562
rect 23480 1498 23532 1504
rect 23860 1426 23888 1838
rect 23848 1420 23900 1426
rect 23848 1362 23900 1368
rect 24044 1358 24072 3334
rect 24136 3126 24164 5063
rect 24228 4010 24256 5578
rect 24676 5568 24728 5574
rect 24676 5510 24728 5516
rect 24688 5234 24716 5510
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24412 2990 24440 3538
rect 24688 3210 24716 4218
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24780 3602 24808 4082
rect 25056 3738 25084 6190
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 25148 4690 25176 5102
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 24872 3346 24900 3402
rect 24872 3318 24992 3346
rect 24688 3182 24900 3210
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24412 2446 24440 2926
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24872 1358 24900 3182
rect 24964 2378 24992 3318
rect 24952 2372 25004 2378
rect 24952 2314 25004 2320
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 23204 1284 23256 1290
rect 23204 1226 23256 1232
rect 25056 1222 25084 3402
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25261 1660 25569 1669
rect 25261 1658 25267 1660
rect 25323 1658 25347 1660
rect 25403 1658 25427 1660
rect 25483 1658 25507 1660
rect 25563 1658 25569 1660
rect 25323 1606 25325 1658
rect 25505 1606 25507 1658
rect 25261 1604 25267 1606
rect 25323 1604 25347 1606
rect 25403 1604 25427 1606
rect 25483 1604 25507 1606
rect 25563 1604 25569 1606
rect 25261 1595 25569 1604
rect 25608 1222 25636 4150
rect 25700 2650 25728 7239
rect 26160 5642 26188 10406
rect 26712 10062 26740 11086
rect 26792 10532 26844 10538
rect 26792 10474 26844 10480
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26252 9654 26280 9930
rect 26514 9752 26570 9761
rect 26712 9722 26740 9998
rect 26514 9687 26570 9696
rect 26700 9716 26752 9722
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26528 9586 26556 9687
rect 26700 9658 26752 9664
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26712 9042 26740 9658
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26804 8974 26832 10474
rect 28000 9178 28028 12922
rect 28276 11898 28304 13874
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27250 9072 27306 9081
rect 27250 9007 27306 9016
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 27158 8800 27214 8809
rect 27158 8735 27214 8744
rect 26330 8392 26386 8401
rect 26330 8327 26332 8336
rect 26384 8327 26386 8336
rect 26332 8298 26384 8304
rect 27172 8090 27200 8735
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26606 7848 26662 7857
rect 26436 6798 26464 7822
rect 26606 7783 26662 7792
rect 26516 7268 26568 7274
rect 26516 7210 26568 7216
rect 26528 6798 26556 7210
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26436 6361 26464 6734
rect 26620 6458 26648 7783
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26422 6352 26478 6361
rect 26422 6287 26478 6296
rect 26436 5778 26464 6287
rect 27068 6112 27120 6118
rect 27068 6054 27120 6060
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26252 5234 26280 5510
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 25778 3632 25834 3641
rect 25778 3567 25834 3576
rect 25792 2922 25820 3567
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 26528 3194 26556 3334
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26238 2952 26294 2961
rect 25780 2916 25832 2922
rect 26238 2887 26240 2896
rect 25780 2858 25832 2864
rect 26292 2887 26294 2896
rect 26240 2858 26292 2864
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 25686 2544 25742 2553
rect 25686 2479 25742 2488
rect 25700 1834 25728 2479
rect 26514 2408 26570 2417
rect 26514 2343 26570 2352
rect 26332 2100 26384 2106
rect 26332 2042 26384 2048
rect 26344 2009 26372 2042
rect 26330 2000 26386 2009
rect 26528 1970 26556 2343
rect 26330 1935 26386 1944
rect 26516 1964 26568 1970
rect 26516 1906 26568 1912
rect 25688 1828 25740 1834
rect 25688 1770 25740 1776
rect 26608 1352 26660 1358
rect 26608 1294 26660 1300
rect 20812 1216 20864 1222
rect 20812 1158 20864 1164
rect 23388 1216 23440 1222
rect 23388 1158 23440 1164
rect 25044 1216 25096 1222
rect 25044 1158 25096 1164
rect 25596 1216 25648 1222
rect 25596 1158 25648 1164
rect 26424 1216 26476 1222
rect 26424 1158 26476 1164
rect 20824 746 20852 1158
rect 21788 1116 22096 1125
rect 21788 1114 21794 1116
rect 21850 1114 21874 1116
rect 21930 1114 21954 1116
rect 22010 1114 22034 1116
rect 22090 1114 22096 1116
rect 21850 1062 21852 1114
rect 22032 1062 22034 1114
rect 21788 1060 21794 1062
rect 21850 1060 21874 1062
rect 21930 1060 21954 1062
rect 22010 1060 22034 1062
rect 22090 1060 22096 1062
rect 21788 1051 22096 1060
rect 23400 746 23428 1158
rect 26436 1018 26464 1158
rect 26424 1012 26476 1018
rect 26424 954 26476 960
rect 26620 950 26648 1294
rect 26608 944 26660 950
rect 26608 886 26660 892
rect 26712 814 26740 3878
rect 26804 2446 26832 5306
rect 27080 3534 27108 6054
rect 27264 5370 27292 9007
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 28356 8016 28408 8022
rect 28356 7958 28408 7964
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27264 4690 27292 5306
rect 27710 5264 27766 5273
rect 27344 5228 27396 5234
rect 27710 5199 27766 5208
rect 27344 5170 27396 5176
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27356 4593 27384 5170
rect 27724 4826 27752 5199
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27618 4720 27674 4729
rect 27618 4655 27674 4664
rect 27632 4622 27660 4655
rect 27620 4616 27672 4622
rect 27342 4584 27398 4593
rect 27620 4558 27672 4564
rect 27342 4519 27398 4528
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27356 4049 27384 4082
rect 27342 4040 27398 4049
rect 27342 3975 27398 3984
rect 28368 3738 28396 7958
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 27068 3528 27120 3534
rect 27068 3470 27120 3476
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 27344 1352 27396 1358
rect 27344 1294 27396 1300
rect 27160 1216 27212 1222
rect 27160 1158 27212 1164
rect 27172 882 27200 1158
rect 27160 876 27212 882
rect 27160 818 27212 824
rect 26700 808 26752 814
rect 26700 750 26752 756
rect 20812 740 20864 746
rect 20812 682 20864 688
rect 23388 740 23440 746
rect 23388 682 23440 688
rect 27356 678 27384 1294
rect 28734 1116 29042 1125
rect 28734 1114 28740 1116
rect 28796 1114 28820 1116
rect 28876 1114 28900 1116
rect 28956 1114 28980 1116
rect 29036 1114 29042 1116
rect 28796 1062 28798 1114
rect 28978 1062 28980 1114
rect 28734 1060 28740 1062
rect 28796 1060 28820 1062
rect 28876 1060 28900 1062
rect 28956 1060 28980 1062
rect 29036 1060 29042 1062
rect 28734 1051 29042 1060
rect 27344 672 27396 678
rect 27344 614 27396 620
rect 15568 604 15620 610
rect 15568 546 15620 552
rect 18880 604 18932 610
rect 18880 546 18932 552
rect 19064 604 19116 610
rect 19064 546 19116 552
<< via2 >>
rect 2502 31340 2558 31376
rect 2502 31320 2504 31340
rect 2504 31320 2556 31340
rect 2556 31320 2558 31340
rect 2134 30268 2136 30288
rect 2136 30268 2188 30288
rect 2188 30268 2190 30288
rect 2134 30232 2190 30268
rect 478 28192 534 28248
rect 478 22072 534 22128
rect 478 20032 534 20088
rect 938 20848 994 20904
rect 570 17992 626 18048
rect 478 15952 534 16008
rect 478 13912 534 13968
rect 754 12688 810 12744
rect 478 9832 534 9888
rect 478 5752 534 5808
rect 2410 29588 2412 29608
rect 2412 29588 2464 29608
rect 2464 29588 2466 29608
rect 2410 29552 2466 29588
rect 1766 23740 1768 23760
rect 1768 23740 1820 23760
rect 1820 23740 1822 23760
rect 1766 23704 1822 23740
rect 3422 32272 3478 32328
rect 4429 32122 4485 32124
rect 4509 32122 4565 32124
rect 4589 32122 4645 32124
rect 4669 32122 4725 32124
rect 4429 32070 4475 32122
rect 4475 32070 4485 32122
rect 4509 32070 4539 32122
rect 4539 32070 4551 32122
rect 4551 32070 4565 32122
rect 4589 32070 4603 32122
rect 4603 32070 4615 32122
rect 4615 32070 4645 32122
rect 4669 32070 4679 32122
rect 4679 32070 4725 32122
rect 4429 32068 4485 32070
rect 4509 32068 4565 32070
rect 4589 32068 4645 32070
rect 4669 32068 4725 32070
rect 2778 30640 2834 30696
rect 3330 30796 3386 30832
rect 3330 30776 3332 30796
rect 3332 30776 3384 30796
rect 3384 30776 3386 30796
rect 2226 25064 2282 25120
rect 1858 22072 1914 22128
rect 1490 21800 1546 21856
rect 1398 16224 1454 16280
rect 2134 22208 2190 22264
rect 2962 23044 3018 23080
rect 2962 23024 2964 23044
rect 2964 23024 3016 23044
rect 3016 23024 3018 23044
rect 2686 22772 2742 22808
rect 2686 22752 2688 22772
rect 2688 22752 2740 22772
rect 2740 22752 2742 22772
rect 2594 22480 2650 22536
rect 2502 21548 2558 21584
rect 2502 21528 2504 21548
rect 2504 21528 2556 21548
rect 2556 21528 2558 21548
rect 2870 22072 2926 22128
rect 3422 25916 3424 25936
rect 3424 25916 3476 25936
rect 3476 25916 3478 25936
rect 3422 25880 3478 25916
rect 2410 20848 2466 20904
rect 2134 20304 2190 20360
rect 2226 20168 2282 20224
rect 2502 20440 2558 20496
rect 2410 19488 2466 19544
rect 2778 21936 2834 21992
rect 2870 19896 2926 19952
rect 2134 18420 2190 18456
rect 2134 18400 2136 18420
rect 2136 18400 2188 18420
rect 2188 18400 2190 18420
rect 2134 14456 2190 14512
rect 1766 14184 1822 14240
rect 1950 13912 2006 13968
rect 2318 12280 2374 12336
rect 3054 21936 3110 21992
rect 3054 21548 3110 21584
rect 3054 21528 3056 21548
rect 3056 21528 3108 21548
rect 3108 21528 3110 21548
rect 3238 22636 3294 22672
rect 3238 22616 3240 22636
rect 3240 22616 3292 22636
rect 3292 22616 3294 22636
rect 3238 22208 3294 22264
rect 3146 20440 3202 20496
rect 4066 30096 4122 30152
rect 5262 31900 5264 31920
rect 5264 31900 5316 31920
rect 5316 31900 5318 31920
rect 5262 31864 5318 31900
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 3790 26152 3846 26208
rect 4158 28600 4214 28656
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 4710 29144 4766 29200
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 4342 28464 4398 28520
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 4066 26852 4122 26888
rect 4066 26832 4068 26852
rect 4068 26832 4120 26852
rect 4120 26832 4122 26852
rect 3974 24112 4030 24168
rect 3422 19896 3478 19952
rect 2962 18536 3018 18592
rect 2686 15544 2742 15600
rect 1766 12008 1822 12064
rect 1398 9596 1400 9616
rect 1400 9596 1452 9616
rect 1452 9596 1454 9616
rect 1398 9560 1454 9596
rect 478 3712 534 3768
rect 1858 11076 1914 11112
rect 1858 11056 1860 11076
rect 1860 11056 1912 11076
rect 1912 11056 1914 11076
rect 1858 9696 1914 9752
rect 1766 9560 1822 9616
rect 1766 9172 1822 9208
rect 1766 9152 1768 9172
rect 1768 9152 1820 9172
rect 1820 9152 1822 9172
rect 1858 5772 1914 5808
rect 1858 5752 1860 5772
rect 1860 5752 1912 5772
rect 1912 5752 1914 5772
rect 2318 8200 2374 8256
rect 3330 17992 3386 18048
rect 3514 19352 3570 19408
rect 2870 12416 2926 12472
rect 3790 18708 3792 18728
rect 3792 18708 3844 18728
rect 3844 18708 3846 18728
rect 3790 18672 3846 18708
rect 3790 17584 3846 17640
rect 3698 16632 3754 16688
rect 2594 10376 2650 10432
rect 3146 10376 3202 10432
rect 3146 9560 3202 9616
rect 3238 9016 3294 9072
rect 3054 7928 3110 7984
rect 2962 6704 3018 6760
rect 1674 2488 1730 2544
rect 2594 1980 2596 2000
rect 2596 1980 2648 2000
rect 2648 1980 2650 2000
rect 2594 1944 2650 1980
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4802 26016 4858 26072
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 5262 27956 5264 27976
rect 5264 27956 5316 27976
rect 5316 27956 5318 27976
rect 5262 27920 5318 27956
rect 5262 26324 5264 26344
rect 5264 26324 5316 26344
rect 5316 26324 5318 26344
rect 4894 25200 4950 25256
rect 4802 24656 4858 24712
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4342 23568 4398 23624
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4618 22480 4674 22536
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4894 23296 4950 23352
rect 4894 22752 4950 22808
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 3974 19896 4030 19952
rect 4434 20884 4436 20904
rect 4436 20884 4488 20904
rect 4488 20884 4490 20904
rect 4434 20848 4490 20884
rect 4158 20168 4214 20224
rect 4434 20460 4490 20496
rect 4434 20440 4436 20460
rect 4436 20440 4488 20460
rect 4488 20440 4490 20460
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4434 19760 4490 19816
rect 5262 26288 5318 26324
rect 5354 24928 5410 24984
rect 5906 27784 5962 27840
rect 5538 24148 5540 24168
rect 5540 24148 5592 24168
rect 5592 24148 5594 24168
rect 5538 24112 5594 24148
rect 5354 22344 5410 22400
rect 5538 21836 5540 21856
rect 5540 21836 5592 21856
rect 5592 21836 5594 21856
rect 5538 21800 5594 21836
rect 5354 21392 5410 21448
rect 5446 21140 5502 21176
rect 5446 21120 5448 21140
rect 5448 21120 5500 21140
rect 5500 21120 5502 21140
rect 5170 20984 5226 21040
rect 5354 20984 5410 21040
rect 5078 20440 5134 20496
rect 4710 19216 4766 19272
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4158 16632 4214 16688
rect 4986 19488 5042 19544
rect 5262 19488 5318 19544
rect 4526 18128 4582 18184
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4342 17740 4398 17776
rect 4342 17720 4344 17740
rect 4344 17720 4396 17740
rect 4396 17720 4398 17740
rect 4986 17856 5042 17912
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 3790 15408 3846 15464
rect 3514 5480 3570 5536
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 5170 18672 5226 18728
rect 5446 20440 5502 20496
rect 5446 20340 5448 20360
rect 5448 20340 5500 20360
rect 5500 20340 5502 20360
rect 5446 20304 5502 20340
rect 5814 24812 5870 24848
rect 5814 24792 5816 24812
rect 5816 24792 5868 24812
rect 5868 24792 5870 24812
rect 5814 23432 5870 23488
rect 5722 23296 5778 23352
rect 5722 23160 5778 23216
rect 5722 22072 5778 22128
rect 6642 26424 6698 26480
rect 6550 25336 6606 25392
rect 6550 25200 6606 25256
rect 6458 24012 6460 24032
rect 6460 24012 6512 24032
rect 6512 24012 6514 24032
rect 6458 23976 6514 24012
rect 5630 19660 5632 19680
rect 5632 19660 5684 19680
rect 5684 19660 5686 19680
rect 5630 19624 5686 19660
rect 5538 19488 5594 19544
rect 5538 18536 5594 18592
rect 6366 22344 6422 22400
rect 6274 21936 6330 21992
rect 6826 28500 6828 28520
rect 6828 28500 6880 28520
rect 6880 28500 6882 28520
rect 6826 28464 6882 28500
rect 6918 26968 6974 27024
rect 6826 25200 6882 25256
rect 7010 24112 7066 24168
rect 6918 23840 6974 23896
rect 7010 23568 7066 23624
rect 6642 21004 6698 21040
rect 6642 20984 6644 21004
rect 6644 20984 6696 21004
rect 6696 20984 6698 21004
rect 6090 17856 6146 17912
rect 5814 17040 5870 17096
rect 4526 14184 4582 14240
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4342 12824 4398 12880
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 3974 10260 4030 10296
rect 3974 10240 3976 10260
rect 3976 10240 4028 10260
rect 4028 10240 4030 10260
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4158 11056 4214 11112
rect 4342 11092 4344 11112
rect 4344 11092 4396 11112
rect 4396 11092 4398 11112
rect 4342 11056 4398 11092
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 5170 13232 5226 13288
rect 5078 12280 5134 12336
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4710 7268 4766 7304
rect 4710 7248 4712 7268
rect 4712 7248 4764 7268
rect 4764 7248 4766 7268
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 4618 6452 4674 6488
rect 4618 6432 4620 6452
rect 4620 6432 4672 6452
rect 4672 6432 4674 6452
rect 5906 13776 5962 13832
rect 4158 6160 4214 6216
rect 4802 6024 4858 6080
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4986 5752 5042 5808
rect 4986 4820 5042 4856
rect 4986 4800 4988 4820
rect 4988 4800 5040 4820
rect 5040 4800 5042 4820
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 5078 3984 5134 4040
rect 5906 12436 5962 12472
rect 5906 12416 5908 12436
rect 5908 12416 5960 12436
rect 5960 12416 5962 12436
rect 5906 11464 5962 11520
rect 5538 8508 5540 8528
rect 5540 8508 5592 8528
rect 5592 8508 5594 8528
rect 5538 8472 5594 8508
rect 5538 8336 5594 8392
rect 5446 6160 5502 6216
rect 5906 10004 5908 10024
rect 5908 10004 5960 10024
rect 5960 10004 5962 10024
rect 5906 9968 5962 10004
rect 5998 9832 6054 9888
rect 5630 3848 5686 3904
rect 5814 5092 5870 5128
rect 5814 5072 5816 5092
rect 5816 5072 5868 5092
rect 5868 5072 5870 5092
rect 5722 3476 5724 3496
rect 5724 3476 5776 3496
rect 5776 3476 5778 3496
rect 5722 3440 5778 3476
rect 5354 3052 5410 3088
rect 5354 3032 5356 3052
rect 5356 3032 5408 3052
rect 5408 3032 5410 3052
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 4802 2352 4858 2408
rect 4429 1658 4485 1660
rect 4509 1658 4565 1660
rect 4589 1658 4645 1660
rect 4669 1658 4725 1660
rect 4429 1606 4475 1658
rect 4475 1606 4485 1658
rect 4509 1606 4539 1658
rect 4539 1606 4551 1658
rect 4551 1606 4565 1658
rect 4589 1606 4603 1658
rect 4603 1606 4615 1658
rect 4615 1606 4645 1658
rect 4669 1606 4679 1658
rect 4679 1606 4725 1658
rect 4429 1604 4485 1606
rect 4509 1604 4565 1606
rect 4589 1604 4645 1606
rect 4669 1604 4725 1606
rect 6458 18128 6514 18184
rect 7902 32666 7958 32668
rect 7982 32666 8038 32668
rect 8062 32666 8118 32668
rect 8142 32666 8198 32668
rect 7902 32614 7948 32666
rect 7948 32614 7958 32666
rect 7982 32614 8012 32666
rect 8012 32614 8024 32666
rect 8024 32614 8038 32666
rect 8062 32614 8076 32666
rect 8076 32614 8088 32666
rect 8088 32614 8118 32666
rect 8142 32614 8152 32666
rect 8152 32614 8198 32666
rect 7902 32612 7958 32614
rect 7982 32612 8038 32614
rect 8062 32612 8118 32614
rect 8142 32612 8198 32614
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 8482 31900 8484 31920
rect 8484 31900 8536 31920
rect 8536 31900 8538 31920
rect 8482 31864 8538 31900
rect 8298 31456 8354 31512
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 7654 30132 7656 30152
rect 7656 30132 7708 30152
rect 7708 30132 7710 30152
rect 7654 30096 7710 30132
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 8298 29008 8354 29064
rect 7286 25336 7342 25392
rect 7286 25064 7342 25120
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 7562 25472 7618 25528
rect 7010 22072 7066 22128
rect 6826 17992 6882 18048
rect 6458 16124 6460 16144
rect 6460 16124 6512 16144
rect 6512 16124 6514 16144
rect 6458 16088 6514 16124
rect 6458 13912 6514 13968
rect 6642 15272 6698 15328
rect 6734 13912 6790 13968
rect 6458 12416 6514 12472
rect 7102 21548 7158 21584
rect 7102 21528 7104 21548
rect 7104 21528 7156 21548
rect 7156 21528 7158 21548
rect 7010 20576 7066 20632
rect 7102 20168 7158 20224
rect 7194 19216 7250 19272
rect 7010 16088 7066 16144
rect 7378 21800 7434 21856
rect 7654 25200 7710 25256
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 9402 31184 9458 31240
rect 8114 25608 8170 25664
rect 8942 26288 8998 26344
rect 8758 26016 8814 26072
rect 9126 26444 9182 26480
rect 9126 26424 9128 26444
rect 9128 26424 9180 26444
rect 9180 26424 9182 26444
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7930 24676 7986 24712
rect 7930 24656 7932 24676
rect 7932 24656 7984 24676
rect 7984 24656 7986 24676
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 8574 23432 8630 23488
rect 8482 23160 8538 23216
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 8482 20712 8538 20768
rect 7654 19896 7710 19952
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7746 19352 7802 19408
rect 7562 17720 7618 17776
rect 8298 19216 8354 19272
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7746 18128 7802 18184
rect 8758 24248 8814 24304
rect 9126 23024 9182 23080
rect 8850 19760 8906 19816
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 8114 17040 8170 17096
rect 7746 16516 7802 16552
rect 7746 16496 7748 16516
rect 7748 16496 7800 16516
rect 7800 16496 7802 16516
rect 7562 16224 7618 16280
rect 7010 13640 7066 13696
rect 6918 13232 6974 13288
rect 6458 12008 6514 12064
rect 6182 7964 6184 7984
rect 6184 7964 6236 7984
rect 6236 7964 6238 7984
rect 6182 7928 6238 7964
rect 6550 9696 6606 9752
rect 6918 12416 6974 12472
rect 6826 12144 6882 12200
rect 6182 6296 6238 6352
rect 7194 13912 7250 13968
rect 7562 15544 7618 15600
rect 7470 15136 7526 15192
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7562 13776 7618 13832
rect 7286 12688 7342 12744
rect 7286 12416 7342 12472
rect 7194 12008 7250 12064
rect 7194 10668 7250 10704
rect 7194 10648 7196 10668
rect 7196 10648 7248 10668
rect 7248 10648 7250 10668
rect 7562 12724 7564 12744
rect 7564 12724 7616 12744
rect 7616 12724 7618 12744
rect 7562 12688 7618 12724
rect 7654 12552 7710 12608
rect 8206 14320 8262 14376
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7930 13932 7986 13968
rect 7930 13912 7932 13932
rect 7932 13912 7984 13932
rect 7984 13912 7986 13932
rect 8022 13368 8078 13424
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 8206 12316 8208 12336
rect 8208 12316 8260 12336
rect 8260 12316 8262 12336
rect 8206 12280 8262 12316
rect 8758 18808 8814 18864
rect 9310 23296 9366 23352
rect 9310 22616 9366 22672
rect 10506 31884 10562 31920
rect 10506 31864 10508 31884
rect 10508 31864 10560 31884
rect 10560 31864 10562 31884
rect 10138 30368 10194 30424
rect 9586 26580 9642 26616
rect 9586 26560 9588 26580
rect 9588 26560 9640 26580
rect 9640 26560 9642 26580
rect 9402 22072 9458 22128
rect 9770 25744 9826 25800
rect 9586 24132 9642 24168
rect 9586 24112 9588 24132
rect 9588 24112 9640 24132
rect 9640 24112 9642 24132
rect 9402 21412 9458 21448
rect 9402 21392 9404 21412
rect 9404 21392 9456 21412
rect 9456 21392 9458 21412
rect 10046 23840 10102 23896
rect 9034 18808 9090 18864
rect 9034 18264 9090 18320
rect 8850 15408 8906 15464
rect 8758 13776 8814 13832
rect 8666 13504 8722 13560
rect 9126 17992 9182 18048
rect 9034 13232 9090 13288
rect 8666 12552 8722 12608
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7838 10412 7840 10432
rect 7840 10412 7892 10432
rect 7892 10412 7894 10432
rect 7838 10376 7894 10412
rect 7654 9832 7710 9888
rect 7654 9152 7710 9208
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7930 9580 7986 9616
rect 7930 9560 7932 9580
rect 7932 9560 7984 9580
rect 7984 9560 7986 9580
rect 7378 7928 7434 7984
rect 6918 7420 6920 7440
rect 6920 7420 6972 7440
rect 6972 7420 6974 7440
rect 6918 7384 6974 7420
rect 6918 7248 6974 7304
rect 6734 5480 6790 5536
rect 6642 5228 6698 5264
rect 6642 5208 6644 5228
rect 6644 5208 6696 5228
rect 6696 5208 6698 5228
rect 7010 5888 7066 5944
rect 7378 4664 7434 4720
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 8850 12416 8906 12472
rect 8114 7284 8116 7304
rect 8116 7284 8168 7304
rect 8168 7284 8170 7304
rect 8114 7248 8170 7284
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 8206 2488 8262 2544
rect 9034 12588 9036 12608
rect 9036 12588 9088 12608
rect 9088 12588 9090 12608
rect 9034 12552 9090 12588
rect 9218 13912 9274 13968
rect 9402 20032 9458 20088
rect 9402 17584 9458 17640
rect 9310 13368 9366 13424
rect 9954 21684 10010 21720
rect 9954 21664 9956 21684
rect 9956 21664 10008 21684
rect 10008 21664 10010 21684
rect 9770 20324 9826 20360
rect 9770 20304 9772 20324
rect 9772 20304 9824 20324
rect 9824 20304 9826 20324
rect 10506 26152 10562 26208
rect 10506 25608 10562 25664
rect 11375 32122 11431 32124
rect 11455 32122 11511 32124
rect 11535 32122 11591 32124
rect 11615 32122 11671 32124
rect 11375 32070 11421 32122
rect 11421 32070 11431 32122
rect 11455 32070 11485 32122
rect 11485 32070 11497 32122
rect 11497 32070 11511 32122
rect 11535 32070 11549 32122
rect 11549 32070 11561 32122
rect 11561 32070 11591 32122
rect 11615 32070 11625 32122
rect 11625 32070 11671 32122
rect 11375 32068 11431 32070
rect 11455 32068 11511 32070
rect 11535 32068 11591 32070
rect 11615 32068 11671 32070
rect 11978 32136 12034 32192
rect 11794 31456 11850 31512
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 11794 30912 11850 30968
rect 10690 29996 10692 30016
rect 10692 29996 10744 30016
rect 10744 29996 10746 30016
rect 10690 29960 10746 29996
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 10690 28056 10746 28112
rect 10506 23976 10562 24032
rect 10506 23160 10562 23216
rect 9770 19080 9826 19136
rect 9770 18536 9826 18592
rect 9862 17756 9864 17776
rect 9864 17756 9916 17776
rect 9916 17756 9918 17776
rect 9862 17720 9918 17756
rect 9586 15272 9642 15328
rect 10322 17740 10378 17776
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11150 27512 11206 27568
rect 11058 27376 11114 27432
rect 11058 25608 11114 25664
rect 11058 25472 11114 25528
rect 10782 21684 10838 21720
rect 10782 21664 10784 21684
rect 10784 21664 10836 21684
rect 10836 21664 10838 21684
rect 10598 20848 10654 20904
rect 10782 19252 10784 19272
rect 10784 19252 10836 19272
rect 10836 19252 10838 19272
rect 10782 19216 10838 19252
rect 10322 17720 10324 17740
rect 10324 17720 10376 17740
rect 10376 17720 10378 17740
rect 10230 17176 10286 17232
rect 9862 16360 9918 16416
rect 10046 16396 10048 16416
rect 10048 16396 10100 16416
rect 10100 16396 10102 16416
rect 10046 16360 10102 16396
rect 10046 16088 10102 16144
rect 9494 13504 9550 13560
rect 9402 12416 9458 12472
rect 8942 11756 8998 11792
rect 8942 11736 8944 11756
rect 8944 11736 8996 11756
rect 8996 11736 8998 11756
rect 8942 11328 8998 11384
rect 8942 9696 8998 9752
rect 9126 11056 9182 11112
rect 9310 11600 9366 11656
rect 9218 10512 9274 10568
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 9402 11192 9458 11248
rect 9402 9596 9404 9616
rect 9404 9596 9456 9616
rect 9456 9596 9458 9616
rect 9402 9560 9458 9596
rect 10230 16516 10286 16552
rect 10230 16496 10232 16516
rect 10232 16496 10284 16516
rect 10284 16496 10286 16516
rect 10782 16360 10838 16416
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11518 24656 11574 24712
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11610 23976 11666 24032
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11886 29824 11942 29880
rect 12254 28872 12310 28928
rect 12254 27784 12310 27840
rect 11794 23316 11850 23352
rect 11794 23296 11796 23316
rect 11796 23296 11848 23316
rect 11848 23296 11850 23316
rect 11058 19352 11114 19408
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11426 20712 11482 20768
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 12714 29280 12770 29336
rect 13726 31084 13728 31104
rect 13728 31084 13780 31104
rect 13780 31084 13782 31104
rect 13726 31048 13782 31084
rect 13726 29688 13782 29744
rect 13358 28736 13414 28792
rect 12898 26968 12954 27024
rect 11610 19372 11666 19408
rect 11610 19352 11612 19372
rect 11612 19352 11664 19372
rect 11664 19352 11666 19372
rect 11058 19080 11114 19136
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11518 18828 11574 18864
rect 11518 18808 11520 18828
rect 11520 18808 11572 18828
rect 11572 18808 11574 18828
rect 11150 18572 11152 18592
rect 11152 18572 11204 18592
rect 11204 18572 11206 18592
rect 11150 18536 11206 18572
rect 11058 18400 11114 18456
rect 11610 18536 11666 18592
rect 11610 18164 11612 18184
rect 11612 18164 11664 18184
rect 11664 18164 11666 18184
rect 11610 18128 11666 18164
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 10874 14340 10930 14376
rect 10874 14320 10876 14340
rect 10876 14320 10928 14340
rect 10928 14320 10930 14340
rect 9954 13640 10010 13696
rect 9954 12416 10010 12472
rect 9770 12008 9826 12064
rect 9678 11892 9734 11928
rect 9678 11872 9680 11892
rect 9680 11872 9732 11892
rect 9732 11872 9734 11892
rect 11426 17196 11482 17232
rect 11426 17176 11428 17196
rect 11428 17176 11480 17196
rect 11480 17176 11482 17196
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11426 16516 11482 16552
rect 11426 16496 11428 16516
rect 11428 16496 11480 16516
rect 11480 16496 11482 16516
rect 11518 16360 11574 16416
rect 11242 16108 11298 16144
rect 11242 16088 11244 16108
rect 11244 16088 11296 16108
rect 11296 16088 11298 16108
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11150 15136 11206 15192
rect 12070 19760 12126 19816
rect 11978 18300 11980 18320
rect 11980 18300 12032 18320
rect 12032 18300 12034 18320
rect 11978 18264 12034 18300
rect 11978 18128 12034 18184
rect 11886 17992 11942 18048
rect 12438 20884 12440 20904
rect 12440 20884 12492 20904
rect 12492 20884 12494 20904
rect 12438 20848 12494 20884
rect 13174 24928 13230 24984
rect 13358 24384 13414 24440
rect 13266 23840 13322 23896
rect 12714 20848 12770 20904
rect 12438 18400 12494 18456
rect 11978 17040 12034 17096
rect 11886 15564 11942 15600
rect 11886 15544 11888 15564
rect 11888 15544 11940 15564
rect 11940 15544 11942 15564
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 10322 13096 10378 13152
rect 10230 12688 10286 12744
rect 10138 11872 10194 11928
rect 10230 11636 10232 11656
rect 10232 11636 10284 11656
rect 10284 11636 10286 11656
rect 10230 11600 10286 11636
rect 10138 11192 10194 11248
rect 9862 10784 9918 10840
rect 10046 10648 10102 10704
rect 9586 9716 9642 9752
rect 9586 9696 9588 9716
rect 9588 9696 9640 9716
rect 9640 9696 9642 9716
rect 9586 8608 9642 8664
rect 9586 8372 9588 8392
rect 9588 8372 9640 8392
rect 9640 8372 9642 8392
rect 9586 8336 9642 8372
rect 9402 6024 9458 6080
rect 9770 6704 9826 6760
rect 10046 10260 10102 10296
rect 10046 10240 10048 10260
rect 10048 10240 10100 10260
rect 10100 10240 10102 10260
rect 10414 11348 10470 11384
rect 10414 11328 10416 11348
rect 10416 11328 10468 11348
rect 10468 11328 10470 11348
rect 10782 12416 10838 12472
rect 11058 13504 11114 13560
rect 11334 14048 11390 14104
rect 12070 14592 12126 14648
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11794 13640 11850 13696
rect 11610 12688 11666 12744
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11702 11872 11758 11928
rect 11610 11600 11666 11656
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 10782 8372 10784 8392
rect 10784 8372 10836 8392
rect 10836 8372 10838 8392
rect 10782 8336 10838 8372
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11610 10104 11666 10160
rect 11242 9560 11298 9616
rect 14848 32666 14904 32668
rect 14928 32666 14984 32668
rect 15008 32666 15064 32668
rect 15088 32666 15144 32668
rect 14848 32614 14894 32666
rect 14894 32614 14904 32666
rect 14928 32614 14958 32666
rect 14958 32614 14970 32666
rect 14970 32614 14984 32666
rect 15008 32614 15022 32666
rect 15022 32614 15034 32666
rect 15034 32614 15064 32666
rect 15088 32614 15098 32666
rect 15098 32614 15144 32666
rect 14848 32612 14904 32614
rect 14928 32612 14984 32614
rect 15008 32612 15064 32614
rect 15088 32612 15144 32614
rect 14094 29280 14150 29336
rect 15290 31628 15292 31648
rect 15292 31628 15344 31648
rect 15344 31628 15346 31648
rect 15290 31592 15346 31628
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 14646 30368 14702 30424
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 14002 26580 14058 26616
rect 14002 26560 14004 26580
rect 14004 26560 14056 26580
rect 14056 26560 14058 26580
rect 13910 25472 13966 25528
rect 13082 20340 13084 20360
rect 13084 20340 13136 20360
rect 13136 20340 13138 20360
rect 13082 20304 13138 20340
rect 13082 20168 13138 20224
rect 12898 19352 12954 19408
rect 12806 18264 12862 18320
rect 13266 19216 13322 19272
rect 14186 26696 14242 26752
rect 15014 29960 15070 30016
rect 14646 29416 14702 29472
rect 14646 29008 14702 29064
rect 14370 27668 14426 27704
rect 14370 27648 14372 27668
rect 14372 27648 14424 27668
rect 14424 27648 14426 27668
rect 14278 23568 14334 23624
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 15474 31048 15530 31104
rect 15290 30540 15292 30560
rect 15292 30540 15344 30560
rect 15344 30540 15346 30560
rect 15290 30504 15346 30540
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 14738 27784 14794 27840
rect 15934 30368 15990 30424
rect 15382 29300 15438 29336
rect 15382 29280 15384 29300
rect 15384 29280 15436 29300
rect 15436 29280 15438 29300
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14646 26188 14648 26208
rect 14648 26188 14700 26208
rect 14700 26188 14702 26208
rect 14646 26152 14702 26188
rect 14554 25744 14610 25800
rect 14554 25200 14610 25256
rect 14554 25064 14610 25120
rect 14830 26560 14886 26616
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14738 25744 14794 25800
rect 15014 25492 15070 25528
rect 15014 25472 15016 25492
rect 15016 25472 15068 25492
rect 15068 25472 15070 25492
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 15014 24384 15070 24440
rect 15290 27240 15346 27296
rect 15474 27104 15530 27160
rect 15290 26560 15346 26616
rect 15290 26188 15292 26208
rect 15292 26188 15344 26208
rect 15344 26188 15346 26208
rect 15290 26152 15346 26188
rect 14462 23604 14464 23624
rect 14464 23604 14516 23624
rect 14516 23604 14518 23624
rect 14462 23568 14518 23604
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 13910 22616 13966 22672
rect 13726 22072 13782 22128
rect 13634 20440 13690 20496
rect 13266 17620 13268 17640
rect 13268 17620 13320 17640
rect 13320 17620 13322 17640
rect 13266 17584 13322 17620
rect 12254 14356 12256 14376
rect 12256 14356 12308 14376
rect 12308 14356 12310 14376
rect 12254 14320 12310 14356
rect 12162 14048 12218 14104
rect 12438 14864 12494 14920
rect 12438 13096 12494 13152
rect 12070 11464 12126 11520
rect 11610 9424 11666 9480
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11334 8744 11390 8800
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11978 10260 12034 10296
rect 11978 10240 11980 10260
rect 11980 10240 12032 10260
rect 12032 10240 12034 10260
rect 11978 9832 12034 9888
rect 13266 16904 13322 16960
rect 13082 15544 13138 15600
rect 14094 21392 14150 21448
rect 14830 23468 14832 23488
rect 14832 23468 14884 23488
rect 14884 23468 14886 23488
rect 14830 23432 14886 23468
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 15014 22208 15070 22264
rect 14186 19080 14242 19136
rect 13910 18672 13966 18728
rect 13818 17876 13874 17912
rect 13818 17856 13820 17876
rect 13820 17856 13872 17876
rect 13872 17856 13874 17876
rect 14002 17992 14058 18048
rect 14002 17856 14058 17912
rect 13910 17448 13966 17504
rect 13542 15952 13598 16008
rect 12714 13776 12770 13832
rect 12254 11892 12310 11928
rect 12254 11872 12256 11892
rect 12256 11872 12308 11892
rect 12308 11872 12310 11892
rect 12254 11600 12310 11656
rect 12254 10784 12310 10840
rect 12530 12280 12586 12336
rect 12162 10104 12218 10160
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11242 6740 11244 6760
rect 11244 6740 11296 6760
rect 11296 6740 11298 6760
rect 11242 6704 11298 6740
rect 8206 1284 8262 1320
rect 8206 1264 8208 1284
rect 8208 1264 8260 1284
rect 8260 1264 8262 1284
rect 7902 1114 7958 1116
rect 7982 1114 8038 1116
rect 8062 1114 8118 1116
rect 8142 1114 8198 1116
rect 7902 1062 7948 1114
rect 7948 1062 7958 1114
rect 7982 1062 8012 1114
rect 8012 1062 8024 1114
rect 8024 1062 8038 1114
rect 8062 1062 8076 1114
rect 8076 1062 8088 1114
rect 8088 1062 8118 1114
rect 8142 1062 8152 1114
rect 8152 1062 8198 1114
rect 7902 1060 7958 1062
rect 7982 1060 8038 1062
rect 8062 1060 8118 1062
rect 8142 1060 8198 1062
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 11978 7248 12034 7304
rect 11375 1658 11431 1660
rect 11455 1658 11511 1660
rect 11535 1658 11591 1660
rect 11615 1658 11671 1660
rect 11375 1606 11421 1658
rect 11421 1606 11431 1658
rect 11455 1606 11485 1658
rect 11485 1606 11497 1658
rect 11497 1606 11511 1658
rect 11535 1606 11549 1658
rect 11549 1606 11561 1658
rect 11561 1606 11591 1658
rect 11615 1606 11625 1658
rect 11625 1606 11671 1658
rect 11375 1604 11431 1606
rect 11455 1604 11511 1606
rect 11535 1604 11591 1606
rect 11615 1604 11671 1606
rect 12162 9288 12218 9344
rect 12346 7928 12402 7984
rect 12162 6840 12218 6896
rect 12898 12688 12954 12744
rect 13358 14456 13414 14512
rect 13542 13776 13598 13832
rect 13542 13232 13598 13288
rect 12530 7928 12586 7984
rect 12438 6704 12494 6760
rect 13082 10648 13138 10704
rect 12898 9424 12954 9480
rect 13174 10512 13230 10568
rect 13174 9968 13230 10024
rect 12898 8744 12954 8800
rect 12990 5480 13046 5536
rect 13910 15408 13966 15464
rect 14002 15136 14058 15192
rect 13726 13932 13782 13968
rect 13726 13912 13728 13932
rect 13728 13912 13780 13932
rect 13780 13912 13782 13932
rect 13726 11736 13782 11792
rect 13450 11056 13506 11112
rect 13450 8608 13506 8664
rect 13450 8336 13506 8392
rect 13910 12144 13966 12200
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14646 19488 14702 19544
rect 14278 14592 14334 14648
rect 15106 19760 15162 19816
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14922 19352 14978 19408
rect 15842 28464 15898 28520
rect 16118 29996 16120 30016
rect 16120 29996 16172 30016
rect 16172 29996 16174 30016
rect 16118 29960 16174 29996
rect 16302 31456 16358 31512
rect 16302 29960 16358 30016
rect 16210 29280 16266 29336
rect 16670 29824 16726 29880
rect 15842 24928 15898 24984
rect 16026 24656 16082 24712
rect 16302 25064 16358 25120
rect 15934 23568 15990 23624
rect 16026 22752 16082 22808
rect 16026 20204 16028 20224
rect 16028 20204 16080 20224
rect 16080 20204 16082 20224
rect 16026 20168 16082 20204
rect 15750 19896 15806 19952
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14646 18264 14702 18320
rect 15014 18148 15070 18184
rect 15014 18128 15016 18148
rect 15016 18128 15068 18148
rect 15068 18128 15070 18148
rect 15290 17992 15346 18048
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14186 13368 14242 13424
rect 14370 13912 14426 13968
rect 14646 14320 14702 14376
rect 14554 13368 14610 13424
rect 13174 6024 13230 6080
rect 13358 5888 13414 5944
rect 13818 6024 13874 6080
rect 13726 5480 13782 5536
rect 13450 2896 13506 2952
rect 14278 11192 14334 11248
rect 14370 9696 14426 9752
rect 15014 14456 15070 14512
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 15106 12844 15162 12880
rect 15106 12824 15108 12844
rect 15108 12824 15160 12844
rect 15160 12824 15162 12844
rect 15106 12316 15108 12336
rect 15108 12316 15160 12336
rect 15160 12316 15162 12336
rect 15106 12280 15162 12316
rect 15474 17856 15530 17912
rect 15382 16088 15438 16144
rect 15658 18944 15714 19000
rect 15658 18400 15714 18456
rect 15658 17992 15714 18048
rect 15658 17756 15660 17776
rect 15660 17756 15712 17776
rect 15712 17756 15714 17776
rect 15658 17720 15714 17756
rect 15842 19216 15898 19272
rect 15658 14728 15714 14784
rect 16302 23568 16358 23624
rect 16486 23976 16542 24032
rect 16578 23432 16634 23488
rect 17130 31864 17186 31920
rect 17590 32136 17646 32192
rect 17498 32000 17554 32056
rect 17406 31864 17462 31920
rect 18321 32122 18377 32124
rect 18401 32122 18457 32124
rect 18481 32122 18537 32124
rect 18561 32122 18617 32124
rect 18321 32070 18367 32122
rect 18367 32070 18377 32122
rect 18401 32070 18431 32122
rect 18431 32070 18443 32122
rect 18443 32070 18457 32122
rect 18481 32070 18495 32122
rect 18495 32070 18507 32122
rect 18507 32070 18537 32122
rect 18561 32070 18571 32122
rect 18571 32070 18617 32122
rect 18321 32068 18377 32070
rect 18401 32068 18457 32070
rect 18481 32068 18537 32070
rect 18561 32068 18617 32070
rect 18050 32000 18106 32056
rect 18418 31864 18474 31920
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 17038 27104 17094 27160
rect 16946 24928 17002 24984
rect 17130 23296 17186 23352
rect 16210 20052 16266 20088
rect 16210 20032 16212 20052
rect 16212 20032 16264 20052
rect 16264 20032 16266 20052
rect 16210 19760 16266 19816
rect 16210 19372 16266 19408
rect 16210 19352 16212 19372
rect 16212 19352 16264 19372
rect 16264 19352 16266 19372
rect 16210 18944 16266 19000
rect 16026 17992 16082 18048
rect 16118 17720 16174 17776
rect 16026 16904 16082 16960
rect 16394 18808 16450 18864
rect 16394 18128 16450 18184
rect 16394 17876 16450 17912
rect 16394 17856 16396 17876
rect 16396 17856 16448 17876
rect 16448 17856 16450 17876
rect 16302 17332 16358 17368
rect 16302 17312 16304 17332
rect 16304 17312 16356 17332
rect 16356 17312 16358 17332
rect 16670 19352 16726 19408
rect 17314 24248 17370 24304
rect 17314 23976 17370 24032
rect 18050 30368 18106 30424
rect 18878 31456 18934 31512
rect 18970 30776 19026 30832
rect 18970 30504 19026 30560
rect 17958 29960 18014 30016
rect 17958 28736 18014 28792
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 18694 28872 18750 28928
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18142 26696 18198 26752
rect 18326 28192 18382 28248
rect 18510 28192 18566 28248
rect 19062 28192 19118 28248
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 18694 27648 18750 27704
rect 18694 27240 18750 27296
rect 19062 27820 19064 27840
rect 19064 27820 19116 27840
rect 19116 27820 19118 27840
rect 19062 27784 19118 27820
rect 19062 27648 19118 27704
rect 18970 27104 19026 27160
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 17682 23568 17738 23624
rect 17314 22072 17370 22128
rect 16946 20712 17002 20768
rect 17774 22072 17830 22128
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18694 23296 18750 23352
rect 17314 20712 17370 20768
rect 17498 20304 17554 20360
rect 17038 18672 17094 18728
rect 16026 15000 16082 15056
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14830 11328 14886 11384
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 15382 11872 15438 11928
rect 15658 13096 15714 13152
rect 15566 12688 15622 12744
rect 15566 12180 15568 12200
rect 15568 12180 15620 12200
rect 15620 12180 15622 12200
rect 15566 12144 15622 12180
rect 15566 12008 15622 12064
rect 15382 11192 15438 11248
rect 15106 10240 15162 10296
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 15106 9596 15108 9616
rect 15108 9596 15160 9616
rect 15160 9596 15162 9616
rect 15106 9560 15162 9596
rect 15014 9424 15070 9480
rect 14462 8880 14518 8936
rect 14278 6024 14334 6080
rect 14278 5480 14334 5536
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14646 8336 14702 8392
rect 15106 8200 15162 8256
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14738 7248 14794 7304
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 15290 9460 15292 9480
rect 15292 9460 15344 9480
rect 15344 9460 15346 9480
rect 15290 9424 15346 9460
rect 15474 9172 15530 9208
rect 15474 9152 15476 9172
rect 15476 9152 15528 9172
rect 15528 9152 15530 9172
rect 16394 17040 16450 17096
rect 16394 16532 16396 16552
rect 16396 16532 16448 16552
rect 16448 16532 16450 16552
rect 16394 16496 16450 16532
rect 16302 15272 16358 15328
rect 16118 13912 16174 13968
rect 16026 12008 16082 12064
rect 16026 11872 16082 11928
rect 15934 11192 15990 11248
rect 16302 13640 16358 13696
rect 16118 10784 16174 10840
rect 15934 10648 15990 10704
rect 15198 6160 15254 6216
rect 15198 5652 15200 5672
rect 15200 5652 15252 5672
rect 15252 5652 15254 5672
rect 15198 5616 15254 5652
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 15474 6996 15530 7032
rect 15474 6976 15476 6996
rect 15476 6976 15528 6996
rect 15528 6976 15530 6996
rect 15474 6724 15530 6760
rect 15474 6704 15476 6724
rect 15476 6704 15528 6724
rect 15528 6704 15530 6724
rect 15474 6432 15530 6488
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 15750 9324 15752 9344
rect 15752 9324 15804 9344
rect 15804 9324 15806 9344
rect 15750 9288 15806 9324
rect 16118 9424 16174 9480
rect 16118 8472 16174 8528
rect 16670 14320 16726 14376
rect 17038 18264 17094 18320
rect 17130 17856 17186 17912
rect 17130 17176 17186 17232
rect 16946 17040 17002 17096
rect 17130 16632 17186 16688
rect 17314 17584 17370 17640
rect 17314 17040 17370 17096
rect 16946 14592 17002 14648
rect 17130 13912 17186 13968
rect 16854 13368 16910 13424
rect 17038 13368 17094 13424
rect 16578 11464 16634 11520
rect 16302 10104 16358 10160
rect 16302 8880 16358 8936
rect 15750 6432 15806 6488
rect 16486 9580 16542 9616
rect 16486 9560 16488 9580
rect 16488 9560 16540 9580
rect 16540 9560 16542 9580
rect 16486 9152 16542 9208
rect 16486 6876 16488 6896
rect 16488 6876 16540 6896
rect 16540 6876 16542 6896
rect 16486 6840 16542 6876
rect 15842 6160 15898 6216
rect 16026 6160 16082 6216
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 14848 1114 14904 1116
rect 14928 1114 14984 1116
rect 15008 1114 15064 1116
rect 15088 1114 15144 1116
rect 14848 1062 14894 1114
rect 14894 1062 14904 1114
rect 14928 1062 14958 1114
rect 14958 1062 14970 1114
rect 14970 1062 14984 1114
rect 15008 1062 15022 1114
rect 15022 1062 15034 1114
rect 15034 1062 15064 1114
rect 15088 1062 15098 1114
rect 15098 1062 15144 1114
rect 14848 1060 14904 1062
rect 14928 1060 14984 1062
rect 15008 1060 15064 1062
rect 15088 1060 15144 1062
rect 16026 6024 16082 6080
rect 16762 9968 16818 10024
rect 16578 5888 16634 5944
rect 17038 9424 17094 9480
rect 18602 22888 18658 22944
rect 19062 23976 19118 24032
rect 18970 23568 19026 23624
rect 21794 32666 21850 32668
rect 21874 32666 21930 32668
rect 21954 32666 22010 32668
rect 22034 32666 22090 32668
rect 21794 32614 21840 32666
rect 21840 32614 21850 32666
rect 21874 32614 21904 32666
rect 21904 32614 21916 32666
rect 21916 32614 21930 32666
rect 21954 32614 21968 32666
rect 21968 32614 21980 32666
rect 21980 32614 22010 32666
rect 22034 32614 22044 32666
rect 22044 32614 22090 32666
rect 21794 32612 21850 32614
rect 21874 32612 21930 32614
rect 21954 32612 22010 32614
rect 22034 32612 22090 32614
rect 20810 31728 20866 31784
rect 20718 31592 20774 31648
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18234 22072 18290 22128
rect 17958 19624 18014 19680
rect 17498 18672 17554 18728
rect 17498 17312 17554 17368
rect 17406 13640 17462 13696
rect 17314 11872 17370 11928
rect 17314 11348 17370 11384
rect 17314 11328 17316 11348
rect 17316 11328 17368 11348
rect 17368 11328 17370 11348
rect 17222 9988 17278 10024
rect 17222 9968 17224 9988
rect 17224 9968 17276 9988
rect 17276 9968 17278 9988
rect 17222 7112 17278 7168
rect 17774 15852 17776 15872
rect 17776 15852 17828 15872
rect 17828 15852 17830 15872
rect 17774 15816 17830 15852
rect 17866 15156 17922 15192
rect 17866 15136 17868 15156
rect 17868 15136 17920 15156
rect 17920 15136 17922 15156
rect 17682 14864 17738 14920
rect 18326 21836 18328 21856
rect 18328 21836 18380 21856
rect 18380 21836 18382 21856
rect 18326 21800 18382 21836
rect 18418 21392 18474 21448
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18234 19488 18290 19544
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18326 18420 18382 18456
rect 18326 18400 18328 18420
rect 18328 18400 18380 18420
rect 18380 18400 18382 18420
rect 19062 22380 19064 22400
rect 19064 22380 19116 22400
rect 19116 22380 19118 22400
rect 19062 22344 19118 22380
rect 18878 21664 18934 21720
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 19062 20984 19118 21040
rect 18326 17720 18382 17776
rect 17774 13676 17776 13696
rect 17776 13676 17828 13696
rect 17828 13676 17830 13696
rect 17774 13640 17830 13676
rect 17498 12436 17554 12472
rect 17498 12416 17500 12436
rect 17500 12416 17552 12436
rect 17552 12416 17554 12436
rect 17498 11756 17554 11792
rect 17498 11736 17500 11756
rect 17500 11736 17552 11756
rect 17552 11736 17554 11756
rect 17866 12824 17922 12880
rect 17866 11872 17922 11928
rect 18142 14456 18198 14512
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18602 16632 18658 16688
rect 18694 16360 18750 16416
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18510 13912 18566 13968
rect 18326 13776 18382 13832
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18786 13776 18842 13832
rect 19338 24520 19394 24576
rect 19430 22228 19486 22264
rect 19706 23432 19762 23488
rect 19706 22888 19762 22944
rect 19430 22208 19432 22228
rect 19432 22208 19484 22228
rect 19484 22208 19486 22228
rect 19246 20576 19302 20632
rect 19246 19624 19302 19680
rect 19430 19080 19486 19136
rect 19338 18944 19394 19000
rect 19614 18944 19670 19000
rect 18970 15272 19026 15328
rect 19246 16360 19302 16416
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18418 11872 18474 11928
rect 18878 12824 18934 12880
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18142 9424 18198 9480
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 17866 7248 17922 7304
rect 19062 13232 19118 13288
rect 19338 16088 19394 16144
rect 19614 17448 19670 17504
rect 18878 9424 18934 9480
rect 18694 8472 18750 8528
rect 18694 8336 18750 8392
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18694 5752 18750 5808
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 19246 11192 19302 11248
rect 20442 26560 20498 26616
rect 19982 22616 20038 22672
rect 19890 22072 19946 22128
rect 20258 22752 20314 22808
rect 20718 25608 20774 25664
rect 20718 25472 20774 25528
rect 20166 21936 20222 21992
rect 20534 22072 20590 22128
rect 20074 21800 20130 21856
rect 19798 18400 19854 18456
rect 19890 17992 19946 18048
rect 20442 21392 20498 21448
rect 20442 19216 20498 19272
rect 20166 19080 20222 19136
rect 19982 17040 20038 17096
rect 19890 16224 19946 16280
rect 19982 14456 20038 14512
rect 19982 14320 20038 14376
rect 20350 18400 20406 18456
rect 20626 20168 20682 20224
rect 21362 27512 21418 27568
rect 21546 27376 21602 27432
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 20902 21956 20958 21992
rect 20902 21936 20904 21956
rect 20904 21936 20956 21956
rect 20956 21936 20958 21956
rect 21454 26696 21510 26752
rect 21638 26560 21694 26616
rect 21638 26152 21694 26208
rect 22190 26152 22246 26208
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21178 23840 21234 23896
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 22834 27240 22890 27296
rect 22650 24520 22706 24576
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 20534 17720 20590 17776
rect 20350 14456 20406 14512
rect 19890 13640 19946 13696
rect 19982 12552 20038 12608
rect 19614 11076 19670 11112
rect 19614 11056 19616 11076
rect 19616 11056 19668 11076
rect 19668 11056 19670 11076
rect 19798 12280 19854 12336
rect 20718 14864 20774 14920
rect 20902 17040 20958 17096
rect 21546 20984 21602 21040
rect 21362 19352 21418 19408
rect 20994 16496 21050 16552
rect 20810 14320 20866 14376
rect 19890 11620 19946 11656
rect 19890 11600 19892 11620
rect 19892 11600 19944 11620
rect 19944 11600 19946 11620
rect 20258 11736 20314 11792
rect 19982 10784 20038 10840
rect 19522 8492 19578 8528
rect 19522 8472 19524 8492
rect 19524 8472 19576 8492
rect 19576 8472 19578 8492
rect 19062 6316 19118 6352
rect 19062 6296 19064 6316
rect 19064 6296 19116 6316
rect 19116 6296 19118 6316
rect 18786 3032 18842 3088
rect 17314 1536 17370 1592
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 17866 1536 17922 1592
rect 18321 1658 18377 1660
rect 18401 1658 18457 1660
rect 18481 1658 18537 1660
rect 18561 1658 18617 1660
rect 18321 1606 18367 1658
rect 18367 1606 18377 1658
rect 18401 1606 18431 1658
rect 18431 1606 18443 1658
rect 18443 1606 18457 1658
rect 18481 1606 18495 1658
rect 18495 1606 18507 1658
rect 18507 1606 18537 1658
rect 18561 1606 18571 1658
rect 18571 1606 18617 1658
rect 18321 1604 18377 1606
rect 18401 1604 18457 1606
rect 18481 1604 18537 1606
rect 18561 1604 18617 1606
rect 19890 7828 19892 7848
rect 19892 7828 19944 7848
rect 19944 7828 19946 7848
rect 19890 7792 19946 7828
rect 19982 7268 20038 7304
rect 19982 7248 19984 7268
rect 19984 7248 20036 7268
rect 20036 7248 20038 7268
rect 21086 16224 21142 16280
rect 20442 8608 20498 8664
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 22742 23296 22798 23352
rect 22558 22208 22614 22264
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21362 15816 21418 15872
rect 21362 14456 21418 14512
rect 21086 11192 21142 11248
rect 19798 3612 19800 3632
rect 19800 3612 19852 3632
rect 19852 3612 19854 3632
rect 19798 3576 19854 3612
rect 20442 3848 20498 3904
rect 19430 2624 19486 2680
rect 20442 3440 20498 3496
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21546 16360 21602 16416
rect 21546 15816 21602 15872
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 23754 29008 23810 29064
rect 23202 26308 23258 26344
rect 23202 26288 23204 26308
rect 23204 26288 23256 26308
rect 23256 26288 23258 26308
rect 23294 25472 23350 25528
rect 23386 24656 23442 24712
rect 23110 24248 23166 24304
rect 23018 23296 23074 23352
rect 24122 27820 24124 27840
rect 24124 27820 24176 27840
rect 24176 27820 24178 27840
rect 23846 24792 23902 24848
rect 23202 21528 23258 21584
rect 22926 20848 22982 20904
rect 23110 19760 23166 19816
rect 23662 23568 23718 23624
rect 22374 14456 22430 14512
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 22190 13912 22246 13968
rect 22098 13812 22100 13832
rect 22100 13812 22152 13832
rect 22152 13812 22154 13832
rect 22098 13776 22154 13812
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 22098 12144 22154 12200
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 22006 8880 22062 8936
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21914 8472 21970 8528
rect 22098 8472 22154 8528
rect 23110 15000 23166 15056
rect 22926 12144 22982 12200
rect 24122 27784 24178 27820
rect 24122 23296 24178 23352
rect 24858 30912 24914 30968
rect 25267 32122 25323 32124
rect 25347 32122 25403 32124
rect 25427 32122 25483 32124
rect 25507 32122 25563 32124
rect 25267 32070 25313 32122
rect 25313 32070 25323 32122
rect 25347 32070 25377 32122
rect 25377 32070 25389 32122
rect 25389 32070 25403 32122
rect 25427 32070 25441 32122
rect 25441 32070 25453 32122
rect 25453 32070 25483 32122
rect 25507 32070 25517 32122
rect 25517 32070 25563 32122
rect 25267 32068 25323 32070
rect 25347 32068 25403 32070
rect 25427 32068 25483 32070
rect 25507 32068 25563 32070
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 24858 30368 24914 30424
rect 24766 28600 24822 28656
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 26146 31184 26202 31240
rect 25870 30368 25926 30424
rect 25870 29180 25872 29200
rect 25872 29180 25924 29200
rect 25924 29180 25926 29200
rect 25870 29144 25926 29180
rect 25778 29008 25834 29064
rect 25134 28872 25190 28928
rect 24950 27648 25006 27704
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 25594 28464 25650 28520
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 25134 27276 25136 27296
rect 25136 27276 25188 27296
rect 25188 27276 25190 27296
rect 25134 27240 25190 27276
rect 25042 26696 25098 26752
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 26238 30268 26240 30288
rect 26240 30268 26292 30288
rect 26292 30268 26294 30288
rect 26238 30232 26294 30268
rect 25686 26424 25742 26480
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25686 25900 25742 25936
rect 25686 25880 25688 25900
rect 25688 25880 25740 25900
rect 25740 25880 25742 25900
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25042 24112 25098 24168
rect 24674 23704 24730 23760
rect 24306 23024 24362 23080
rect 24582 23160 24638 23216
rect 24674 22500 24730 22536
rect 24674 22480 24676 22500
rect 24676 22480 24728 22500
rect 24728 22480 24730 22500
rect 24306 20304 24362 20360
rect 23294 12588 23296 12608
rect 23296 12588 23348 12608
rect 23348 12588 23350 12608
rect 23294 12552 23350 12588
rect 22742 11600 22798 11656
rect 22834 9696 22890 9752
rect 22374 8744 22430 8800
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 20994 6180 21050 6216
rect 20994 6160 20996 6180
rect 20996 6160 21048 6180
rect 21048 6160 21050 6180
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 21178 2080 21234 2136
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25686 23160 25742 23216
rect 26054 26968 26110 27024
rect 27066 31320 27122 31376
rect 26422 30640 26478 30696
rect 26514 27920 26570 27976
rect 26146 26832 26202 26888
rect 25870 25764 25926 25800
rect 25870 25744 25872 25764
rect 25872 25744 25924 25764
rect 25924 25744 25926 25764
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 27802 30812 27804 30832
rect 27804 30812 27856 30832
rect 27856 30812 27858 30832
rect 27802 30776 27858 30812
rect 27618 30096 27674 30152
rect 27802 29688 27858 29744
rect 27158 29552 27214 29608
rect 28740 32666 28796 32668
rect 28820 32666 28876 32668
rect 28900 32666 28956 32668
rect 28980 32666 29036 32668
rect 28740 32614 28786 32666
rect 28786 32614 28796 32666
rect 28820 32614 28850 32666
rect 28850 32614 28862 32666
rect 28862 32614 28876 32666
rect 28900 32614 28914 32666
rect 28914 32614 28926 32666
rect 28926 32614 28956 32666
rect 28980 32614 28990 32666
rect 28990 32614 29036 32666
rect 28740 32612 28796 32614
rect 28820 32612 28876 32614
rect 28900 32612 28956 32614
rect 28980 32612 29036 32614
rect 27618 28076 27674 28112
rect 27618 28056 27620 28076
rect 27620 28056 27672 28076
rect 27672 28056 27674 28076
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 27986 25336 28042 25392
rect 25870 20984 25926 21040
rect 24674 19352 24730 19408
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 24582 16904 24638 16960
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 24306 14864 24362 14920
rect 26606 22072 26662 22128
rect 27434 21936 27490 21992
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 27802 17756 27804 17776
rect 27804 17756 27856 17776
rect 27856 17756 27858 17776
rect 27802 17720 27858 17756
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25502 13948 25504 13968
rect 25504 13948 25556 13968
rect 25556 13948 25558 13968
rect 25502 13912 25558 13948
rect 24398 12688 24454 12744
rect 22926 7928 22982 7984
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25318 12688 25374 12744
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25134 12144 25190 12200
rect 25042 11056 25098 11112
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 27710 13776 27766 13832
rect 26974 11736 27030 11792
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 24766 9424 24822 9480
rect 24030 6840 24086 6896
rect 23386 6332 23388 6352
rect 23388 6332 23440 6352
rect 23440 6332 23442 6352
rect 23386 6296 23442 6332
rect 22374 4120 22430 4176
rect 21914 3460 21970 3496
rect 21914 3440 21916 3460
rect 21916 3440 21968 3460
rect 21968 3440 21970 3460
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21914 2624 21970 2680
rect 21546 2080 21602 2136
rect 23386 4156 23388 4176
rect 23388 4156 23440 4176
rect 23440 4156 23442 4176
rect 23386 4120 23442 4156
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25226 8880 25282 8936
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25686 7248 25742 7304
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 24122 5072 24178 5128
rect 23386 3848 23442 3904
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 25267 1658 25323 1660
rect 25347 1658 25403 1660
rect 25427 1658 25483 1660
rect 25507 1658 25563 1660
rect 25267 1606 25313 1658
rect 25313 1606 25323 1658
rect 25347 1606 25377 1658
rect 25377 1606 25389 1658
rect 25389 1606 25403 1658
rect 25427 1606 25441 1658
rect 25441 1606 25453 1658
rect 25453 1606 25483 1658
rect 25507 1606 25517 1658
rect 25517 1606 25563 1658
rect 25267 1604 25323 1606
rect 25347 1604 25403 1606
rect 25427 1604 25483 1606
rect 25507 1604 25563 1606
rect 26514 9696 26570 9752
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 27250 9016 27306 9072
rect 27158 8744 27214 8800
rect 26330 8356 26386 8392
rect 26330 8336 26332 8356
rect 26332 8336 26384 8356
rect 26384 8336 26386 8356
rect 26606 7792 26662 7848
rect 26422 6296 26478 6352
rect 25778 3576 25834 3632
rect 26238 2916 26294 2952
rect 26238 2896 26240 2916
rect 26240 2896 26292 2916
rect 26292 2896 26294 2916
rect 25686 2488 25742 2544
rect 26514 2352 26570 2408
rect 26330 1944 26386 2000
rect 21794 1114 21850 1116
rect 21874 1114 21930 1116
rect 21954 1114 22010 1116
rect 22034 1114 22090 1116
rect 21794 1062 21840 1114
rect 21840 1062 21850 1114
rect 21874 1062 21904 1114
rect 21904 1062 21916 1114
rect 21916 1062 21930 1114
rect 21954 1062 21968 1114
rect 21968 1062 21980 1114
rect 21980 1062 22010 1114
rect 22034 1062 22044 1114
rect 22044 1062 22090 1114
rect 21794 1060 21850 1062
rect 21874 1060 21930 1062
rect 21954 1060 22010 1062
rect 22034 1060 22090 1062
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 27710 5208 27766 5264
rect 27618 4664 27674 4720
rect 27342 4528 27398 4584
rect 27342 3984 27398 4040
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 28740 1114 28796 1116
rect 28820 1114 28876 1116
rect 28900 1114 28956 1116
rect 28980 1114 29036 1116
rect 28740 1062 28786 1114
rect 28786 1062 28796 1114
rect 28820 1062 28850 1114
rect 28850 1062 28862 1114
rect 28862 1062 28876 1114
rect 28900 1062 28914 1114
rect 28914 1062 28926 1114
rect 28926 1062 28956 1114
rect 28980 1062 28990 1114
rect 28990 1062 29036 1114
rect 28740 1060 28796 1062
rect 28820 1060 28876 1062
rect 28900 1060 28956 1062
rect 28980 1060 29036 1062
<< metal3 >>
rect 7892 32672 8208 32673
rect 7892 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8208 32672
rect 7892 32607 8208 32608
rect 14838 32672 15154 32673
rect 14838 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15154 32672
rect 14838 32607 15154 32608
rect 21784 32672 22100 32673
rect 21784 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22100 32672
rect 21784 32607 22100 32608
rect 28730 32672 29046 32673
rect 28730 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29046 32672
rect 28730 32607 29046 32608
rect 0 32330 400 32360
rect 3417 32330 3483 32333
rect 0 32328 3483 32330
rect 0 32272 3422 32328
rect 3478 32272 3483 32328
rect 0 32270 3483 32272
rect 0 32240 400 32270
rect 3417 32267 3483 32270
rect 11973 32194 12039 32197
rect 17585 32194 17651 32197
rect 11973 32192 17651 32194
rect 11973 32136 11978 32192
rect 12034 32136 17590 32192
rect 17646 32136 17651 32192
rect 11973 32134 17651 32136
rect 11973 32131 12039 32134
rect 17585 32131 17651 32134
rect 4419 32128 4735 32129
rect 4419 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4735 32128
rect 4419 32063 4735 32064
rect 11365 32128 11681 32129
rect 11365 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11681 32128
rect 11365 32063 11681 32064
rect 18311 32128 18627 32129
rect 18311 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18627 32128
rect 18311 32063 18627 32064
rect 25257 32128 25573 32129
rect 25257 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25573 32128
rect 25257 32063 25573 32064
rect 17493 32058 17559 32061
rect 18045 32058 18111 32061
rect 17493 32056 18111 32058
rect 17493 32000 17498 32056
rect 17554 32000 18050 32056
rect 18106 32000 18111 32056
rect 17493 31998 18111 32000
rect 17493 31995 17559 31998
rect 18045 31995 18111 31998
rect 5257 31922 5323 31925
rect 8477 31922 8543 31925
rect 5257 31920 8543 31922
rect 5257 31864 5262 31920
rect 5318 31864 8482 31920
rect 8538 31864 8543 31920
rect 5257 31862 8543 31864
rect 5257 31859 5323 31862
rect 8477 31859 8543 31862
rect 10501 31922 10567 31925
rect 17125 31922 17191 31925
rect 10501 31920 17191 31922
rect 10501 31864 10506 31920
rect 10562 31864 17130 31920
rect 17186 31864 17191 31920
rect 10501 31862 17191 31864
rect 10501 31859 10567 31862
rect 17125 31859 17191 31862
rect 17401 31922 17467 31925
rect 18413 31922 18479 31925
rect 17401 31920 18479 31922
rect 17401 31864 17406 31920
rect 17462 31864 18418 31920
rect 18474 31864 18479 31920
rect 17401 31862 18479 31864
rect 17401 31859 17467 31862
rect 18413 31859 18479 31862
rect 14590 31724 14596 31788
rect 14660 31786 14666 31788
rect 20805 31786 20871 31789
rect 14660 31784 20871 31786
rect 14660 31728 20810 31784
rect 20866 31728 20871 31784
rect 14660 31726 20871 31728
rect 14660 31724 14666 31726
rect 20805 31723 20871 31726
rect 15285 31650 15351 31653
rect 15878 31650 15884 31652
rect 15285 31648 15884 31650
rect 15285 31592 15290 31648
rect 15346 31592 15884 31648
rect 15285 31590 15884 31592
rect 15285 31587 15351 31590
rect 15878 31588 15884 31590
rect 15948 31650 15954 31652
rect 20713 31650 20779 31653
rect 15948 31648 20779 31650
rect 15948 31592 20718 31648
rect 20774 31592 20779 31648
rect 15948 31590 20779 31592
rect 15948 31588 15954 31590
rect 20713 31587 20779 31590
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 8293 31514 8359 31517
rect 11789 31514 11855 31517
rect 8293 31512 11855 31514
rect 8293 31456 8298 31512
rect 8354 31456 11794 31512
rect 11850 31456 11855 31512
rect 8293 31454 11855 31456
rect 8293 31451 8359 31454
rect 11789 31451 11855 31454
rect 16297 31514 16363 31517
rect 18873 31514 18939 31517
rect 16297 31512 18939 31514
rect 16297 31456 16302 31512
rect 16358 31456 18878 31512
rect 18934 31456 18939 31512
rect 16297 31454 18939 31456
rect 16297 31451 16363 31454
rect 18873 31451 18939 31454
rect 2497 31378 2563 31381
rect 27061 31378 27127 31381
rect 2497 31376 27127 31378
rect 2497 31320 2502 31376
rect 2558 31320 27066 31376
rect 27122 31320 27127 31376
rect 2497 31318 27127 31320
rect 2497 31315 2563 31318
rect 27061 31315 27127 31318
rect 9397 31242 9463 31245
rect 26141 31242 26207 31245
rect 9397 31240 26207 31242
rect 9397 31184 9402 31240
rect 9458 31184 26146 31240
rect 26202 31184 26207 31240
rect 9397 31182 26207 31184
rect 9397 31179 9463 31182
rect 26141 31179 26207 31182
rect 13721 31106 13787 31109
rect 15469 31106 15535 31109
rect 13721 31104 15535 31106
rect 13721 31048 13726 31104
rect 13782 31048 15474 31104
rect 15530 31048 15535 31104
rect 13721 31046 15535 31048
rect 13721 31043 13787 31046
rect 15469 31043 15535 31046
rect 4419 31040 4735 31041
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 11789 30970 11855 30973
rect 24853 30970 24919 30973
rect 11789 30968 17418 30970
rect 11789 30912 11794 30968
rect 11850 30912 17418 30968
rect 11789 30910 17418 30912
rect 11789 30907 11855 30910
rect 3325 30834 3391 30837
rect 17166 30834 17172 30836
rect 3325 30832 17172 30834
rect 3325 30776 3330 30832
rect 3386 30776 17172 30832
rect 3325 30774 17172 30776
rect 3325 30771 3391 30774
rect 17166 30772 17172 30774
rect 17236 30772 17242 30836
rect 17358 30834 17418 30910
rect 18830 30968 24919 30970
rect 18830 30912 24858 30968
rect 24914 30912 24919 30968
rect 18830 30910 24919 30912
rect 18830 30834 18890 30910
rect 24853 30907 24919 30910
rect 17358 30774 18890 30834
rect 18965 30834 19031 30837
rect 27797 30834 27863 30837
rect 18965 30832 27863 30834
rect 18965 30776 18970 30832
rect 19026 30776 27802 30832
rect 27858 30776 27863 30832
rect 18965 30774 27863 30776
rect 18965 30771 19031 30774
rect 27797 30771 27863 30774
rect 2773 30698 2839 30701
rect 26417 30698 26483 30701
rect 2773 30696 26483 30698
rect 2773 30640 2778 30696
rect 2834 30640 26422 30696
rect 26478 30640 26483 30696
rect 2773 30638 26483 30640
rect 2773 30635 2839 30638
rect 26417 30635 26483 30638
rect 15285 30562 15351 30565
rect 18965 30562 19031 30565
rect 15285 30560 19031 30562
rect 15285 30504 15290 30560
rect 15346 30504 18970 30560
rect 19026 30504 19031 30560
rect 15285 30502 19031 30504
rect 15285 30499 15351 30502
rect 18965 30499 19031 30502
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 28730 30431 29046 30432
rect 10133 30426 10199 30429
rect 14641 30426 14707 30429
rect 10133 30424 14707 30426
rect 10133 30368 10138 30424
rect 10194 30368 14646 30424
rect 14702 30368 14707 30424
rect 10133 30366 14707 30368
rect 10133 30363 10199 30366
rect 14641 30363 14707 30366
rect 15929 30426 15995 30429
rect 18045 30426 18111 30429
rect 15929 30424 18111 30426
rect 15929 30368 15934 30424
rect 15990 30368 18050 30424
rect 18106 30368 18111 30424
rect 15929 30366 18111 30368
rect 15929 30363 15995 30366
rect 18045 30363 18111 30366
rect 24853 30426 24919 30429
rect 25865 30426 25931 30429
rect 24853 30424 25931 30426
rect 24853 30368 24858 30424
rect 24914 30368 25870 30424
rect 25926 30368 25931 30424
rect 24853 30366 25931 30368
rect 24853 30363 24919 30366
rect 25865 30363 25931 30366
rect 0 30290 400 30320
rect 2129 30290 2195 30293
rect 26233 30290 26299 30293
rect 0 30230 1962 30290
rect 0 30200 400 30230
rect 1902 30154 1962 30230
rect 2129 30288 26299 30290
rect 2129 30232 2134 30288
rect 2190 30232 26238 30288
rect 26294 30232 26299 30288
rect 2129 30230 26299 30232
rect 2129 30227 2195 30230
rect 26233 30227 26299 30230
rect 4061 30154 4127 30157
rect 1902 30152 4127 30154
rect 1902 30096 4066 30152
rect 4122 30096 4127 30152
rect 1902 30094 4127 30096
rect 4061 30091 4127 30094
rect 7649 30154 7715 30157
rect 27613 30154 27679 30157
rect 7649 30152 27679 30154
rect 7649 30096 7654 30152
rect 7710 30096 27618 30152
rect 27674 30096 27679 30152
rect 7649 30094 27679 30096
rect 7649 30091 7715 30094
rect 27613 30091 27679 30094
rect 10542 29956 10548 30020
rect 10612 30018 10618 30020
rect 10685 30018 10751 30021
rect 10612 30016 10751 30018
rect 10612 29960 10690 30016
rect 10746 29960 10751 30016
rect 10612 29958 10751 29960
rect 10612 29956 10618 29958
rect 10685 29955 10751 29958
rect 15009 30018 15075 30021
rect 16113 30018 16179 30021
rect 15009 30016 16179 30018
rect 15009 29960 15014 30016
rect 15070 29960 16118 30016
rect 16174 29960 16179 30016
rect 15009 29958 16179 29960
rect 15009 29955 15075 29958
rect 16113 29955 16179 29958
rect 16297 30018 16363 30021
rect 17953 30018 18019 30021
rect 16297 30016 18019 30018
rect 16297 29960 16302 30016
rect 16358 29960 17958 30016
rect 18014 29960 18019 30016
rect 16297 29958 18019 29960
rect 16297 29955 16363 29958
rect 17953 29955 18019 29958
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 11881 29882 11947 29885
rect 16665 29882 16731 29885
rect 11881 29880 16731 29882
rect 11881 29824 11886 29880
rect 11942 29824 16670 29880
rect 16726 29824 16731 29880
rect 11881 29822 16731 29824
rect 11881 29819 11947 29822
rect 16665 29819 16731 29822
rect 13721 29746 13787 29749
rect 27797 29746 27863 29749
rect 13721 29744 27863 29746
rect 13721 29688 13726 29744
rect 13782 29688 27802 29744
rect 27858 29688 27863 29744
rect 13721 29686 27863 29688
rect 13721 29683 13787 29686
rect 27797 29683 27863 29686
rect 2405 29610 2471 29613
rect 27153 29610 27219 29613
rect 2405 29608 27219 29610
rect 2405 29552 2410 29608
rect 2466 29552 27158 29608
rect 27214 29552 27219 29608
rect 2405 29550 27219 29552
rect 2405 29547 2471 29550
rect 27153 29547 27219 29550
rect 14641 29474 14707 29477
rect 12390 29472 14707 29474
rect 12390 29416 14646 29472
rect 14702 29416 14707 29472
rect 12390 29414 14707 29416
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 12390 29338 12450 29414
rect 14641 29411 14707 29414
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 8342 29278 12450 29338
rect 12709 29338 12775 29341
rect 14089 29338 14155 29341
rect 12709 29336 14155 29338
rect 12709 29280 12714 29336
rect 12770 29280 14094 29336
rect 14150 29280 14155 29336
rect 12709 29278 14155 29280
rect 4705 29202 4771 29205
rect 8342 29202 8402 29278
rect 12709 29275 12775 29278
rect 14089 29275 14155 29278
rect 15377 29338 15443 29341
rect 16205 29338 16271 29341
rect 15377 29336 16271 29338
rect 15377 29280 15382 29336
rect 15438 29280 16210 29336
rect 16266 29280 16271 29336
rect 15377 29278 16271 29280
rect 15377 29275 15443 29278
rect 16205 29275 16271 29278
rect 25865 29202 25931 29205
rect 4705 29200 8402 29202
rect 4705 29144 4710 29200
rect 4766 29144 8402 29200
rect 4705 29142 8402 29144
rect 12390 29200 25931 29202
rect 12390 29144 25870 29200
rect 25926 29144 25931 29200
rect 12390 29142 25931 29144
rect 4705 29139 4771 29142
rect 8293 29066 8359 29069
rect 12390 29066 12450 29142
rect 25865 29139 25931 29142
rect 8293 29064 12450 29066
rect 8293 29008 8298 29064
rect 8354 29008 12450 29064
rect 8293 29006 12450 29008
rect 14641 29066 14707 29069
rect 23749 29066 23815 29069
rect 25773 29066 25839 29069
rect 14641 29064 25839 29066
rect 14641 29008 14646 29064
rect 14702 29008 23754 29064
rect 23810 29008 25778 29064
rect 25834 29008 25839 29064
rect 14641 29006 25839 29008
rect 8293 29003 8359 29006
rect 14641 29003 14707 29006
rect 23749 29003 23815 29006
rect 25773 29003 25839 29006
rect 12249 28930 12315 28933
rect 18689 28930 18755 28933
rect 25129 28930 25195 28933
rect 12249 28928 18154 28930
rect 12249 28872 12254 28928
rect 12310 28872 18154 28928
rect 12249 28870 18154 28872
rect 12249 28867 12315 28870
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 13353 28794 13419 28797
rect 17953 28794 18019 28797
rect 13353 28792 18019 28794
rect 13353 28736 13358 28792
rect 13414 28736 17958 28792
rect 18014 28736 18019 28792
rect 13353 28734 18019 28736
rect 13353 28731 13419 28734
rect 17953 28731 18019 28734
rect 4153 28658 4219 28661
rect 17902 28658 17908 28660
rect 4153 28656 17908 28658
rect 4153 28600 4158 28656
rect 4214 28600 17908 28656
rect 4153 28598 17908 28600
rect 4153 28595 4219 28598
rect 17902 28596 17908 28598
rect 17972 28596 17978 28660
rect 18094 28658 18154 28870
rect 18689 28928 25195 28930
rect 18689 28872 18694 28928
rect 18750 28872 25134 28928
rect 25190 28872 25195 28928
rect 18689 28870 25195 28872
rect 18689 28867 18755 28870
rect 25129 28867 25195 28870
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 24761 28658 24827 28661
rect 18094 28656 24827 28658
rect 18094 28600 24766 28656
rect 24822 28600 24827 28656
rect 18094 28598 24827 28600
rect 24761 28595 24827 28598
rect 4337 28522 4403 28525
rect 5206 28522 5212 28524
rect 4337 28520 5212 28522
rect 4337 28464 4342 28520
rect 4398 28464 5212 28520
rect 4337 28462 5212 28464
rect 4337 28459 4403 28462
rect 5206 28460 5212 28462
rect 5276 28460 5282 28524
rect 6821 28522 6887 28525
rect 15837 28522 15903 28525
rect 25589 28522 25655 28525
rect 6821 28520 15903 28522
rect 6821 28464 6826 28520
rect 6882 28464 15842 28520
rect 15898 28464 15903 28520
rect 6821 28462 15903 28464
rect 6821 28459 6887 28462
rect 15837 28459 15903 28462
rect 16990 28520 25655 28522
rect 16990 28464 25594 28520
rect 25650 28464 25655 28520
rect 16990 28462 25655 28464
rect 7892 28320 8208 28321
rect 0 28250 400 28280
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 473 28250 539 28253
rect 0 28248 539 28250
rect 0 28192 478 28248
rect 534 28192 539 28248
rect 0 28190 539 28192
rect 0 28160 400 28190
rect 473 28187 539 28190
rect 10685 28114 10751 28117
rect 16990 28114 17050 28462
rect 25589 28459 25655 28462
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 17350 28188 17356 28252
rect 17420 28250 17426 28252
rect 18321 28250 18387 28253
rect 17420 28248 18387 28250
rect 17420 28192 18326 28248
rect 18382 28192 18387 28248
rect 17420 28190 18387 28192
rect 17420 28188 17426 28190
rect 18321 28187 18387 28190
rect 18505 28250 18571 28253
rect 19057 28250 19123 28253
rect 18505 28248 19123 28250
rect 18505 28192 18510 28248
rect 18566 28192 19062 28248
rect 19118 28192 19123 28248
rect 18505 28190 19123 28192
rect 18505 28187 18571 28190
rect 19057 28187 19123 28190
rect 10685 28112 17050 28114
rect 10685 28056 10690 28112
rect 10746 28056 17050 28112
rect 10685 28054 17050 28056
rect 10685 28051 10751 28054
rect 17166 28052 17172 28116
rect 17236 28114 17242 28116
rect 27613 28114 27679 28117
rect 17236 28112 27679 28114
rect 17236 28056 27618 28112
rect 27674 28056 27679 28112
rect 17236 28054 27679 28056
rect 17236 28052 17242 28054
rect 27613 28051 27679 28054
rect 5257 27978 5323 27981
rect 26509 27978 26575 27981
rect 5257 27976 26575 27978
rect 5257 27920 5262 27976
rect 5318 27920 26514 27976
rect 26570 27920 26575 27976
rect 5257 27918 26575 27920
rect 5257 27915 5323 27918
rect 26509 27915 26575 27918
rect 5574 27780 5580 27844
rect 5644 27842 5650 27844
rect 5901 27842 5967 27845
rect 5644 27840 5967 27842
rect 5644 27784 5906 27840
rect 5962 27784 5967 27840
rect 5644 27782 5967 27784
rect 5644 27780 5650 27782
rect 5901 27779 5967 27782
rect 12249 27842 12315 27845
rect 14733 27842 14799 27845
rect 19057 27842 19123 27845
rect 12249 27840 14799 27842
rect 12249 27784 12254 27840
rect 12310 27784 14738 27840
rect 14794 27784 14799 27840
rect 12249 27782 14799 27784
rect 12249 27779 12315 27782
rect 14733 27779 14799 27782
rect 18692 27840 19123 27842
rect 18692 27784 19062 27840
rect 19118 27784 19123 27840
rect 18692 27782 19123 27784
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 18692 27709 18752 27782
rect 19057 27779 19123 27782
rect 19374 27780 19380 27844
rect 19444 27842 19450 27844
rect 24117 27842 24183 27845
rect 19444 27840 24183 27842
rect 19444 27784 24122 27840
rect 24178 27784 24183 27840
rect 19444 27782 24183 27784
rect 19444 27780 19450 27782
rect 24117 27779 24183 27782
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 14365 27708 14431 27709
rect 14365 27704 14412 27708
rect 14476 27706 14482 27708
rect 14365 27648 14370 27704
rect 14365 27644 14412 27648
rect 14476 27646 14522 27706
rect 18689 27704 18755 27709
rect 18689 27648 18694 27704
rect 18750 27648 18755 27704
rect 14476 27644 14482 27646
rect 14365 27643 14431 27644
rect 18689 27643 18755 27648
rect 19057 27706 19123 27709
rect 24945 27706 25011 27709
rect 19057 27704 25011 27706
rect 19057 27648 19062 27704
rect 19118 27648 24950 27704
rect 25006 27648 25011 27704
rect 19057 27646 25011 27648
rect 19057 27643 19123 27646
rect 24945 27643 25011 27646
rect 11145 27570 11211 27573
rect 21357 27570 21423 27573
rect 11145 27568 21423 27570
rect 11145 27512 11150 27568
rect 11206 27512 21362 27568
rect 21418 27512 21423 27568
rect 11145 27510 21423 27512
rect 11145 27507 11211 27510
rect 21357 27507 21423 27510
rect 11053 27434 11119 27437
rect 21541 27434 21607 27437
rect 11053 27432 21607 27434
rect 11053 27376 11058 27432
rect 11114 27376 21546 27432
rect 21602 27376 21607 27432
rect 11053 27374 21607 27376
rect 11053 27371 11119 27374
rect 21541 27371 21607 27374
rect 15285 27298 15351 27301
rect 18689 27298 18755 27301
rect 15285 27296 18755 27298
rect 15285 27240 15290 27296
rect 15346 27240 18694 27296
rect 18750 27240 18755 27296
rect 15285 27238 18755 27240
rect 15285 27235 15351 27238
rect 18689 27235 18755 27238
rect 22829 27298 22895 27301
rect 25129 27298 25195 27301
rect 22829 27296 25195 27298
rect 22829 27240 22834 27296
rect 22890 27240 25134 27296
rect 25190 27240 25195 27296
rect 22829 27238 25195 27240
rect 22829 27235 22895 27238
rect 25129 27235 25195 27238
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 15469 27162 15535 27165
rect 17033 27162 17099 27165
rect 18965 27162 19031 27165
rect 15469 27160 19031 27162
rect 15469 27104 15474 27160
rect 15530 27104 17038 27160
rect 17094 27104 18970 27160
rect 19026 27104 19031 27160
rect 15469 27102 19031 27104
rect 15469 27099 15535 27102
rect 17033 27099 17099 27102
rect 18965 27099 19031 27102
rect 6913 27026 6979 27029
rect 12893 27026 12959 27029
rect 26049 27026 26115 27029
rect 6913 27024 26115 27026
rect 6913 26968 6918 27024
rect 6974 26968 12898 27024
rect 12954 26968 26054 27024
rect 26110 26968 26115 27024
rect 6913 26966 26115 26968
rect 6913 26963 6979 26966
rect 12893 26963 12959 26966
rect 26049 26963 26115 26966
rect 4061 26890 4127 26893
rect 26141 26890 26207 26893
rect 4061 26888 26207 26890
rect 4061 26832 4066 26888
rect 4122 26832 26146 26888
rect 26202 26832 26207 26888
rect 4061 26830 26207 26832
rect 4061 26827 4127 26830
rect 26141 26827 26207 26830
rect 13302 26692 13308 26756
rect 13372 26754 13378 26756
rect 14181 26754 14247 26757
rect 18137 26754 18203 26757
rect 13372 26752 18203 26754
rect 13372 26696 14186 26752
rect 14242 26696 18142 26752
rect 18198 26696 18203 26752
rect 13372 26694 18203 26696
rect 13372 26692 13378 26694
rect 14181 26691 14247 26694
rect 18137 26691 18203 26694
rect 21449 26754 21515 26757
rect 25037 26754 25103 26757
rect 21449 26752 25103 26754
rect 21449 26696 21454 26752
rect 21510 26696 25042 26752
rect 25098 26696 25103 26752
rect 21449 26694 25103 26696
rect 21449 26691 21515 26694
rect 25037 26691 25103 26694
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 5206 26556 5212 26620
rect 5276 26618 5282 26620
rect 9581 26618 9647 26621
rect 5276 26616 9647 26618
rect 5276 26560 9586 26616
rect 9642 26560 9647 26616
rect 5276 26558 9647 26560
rect 5276 26556 5282 26558
rect 9581 26555 9647 26558
rect 13997 26620 14063 26621
rect 13997 26616 14044 26620
rect 14108 26618 14114 26620
rect 14825 26618 14891 26621
rect 15285 26618 15351 26621
rect 13997 26560 14002 26616
rect 13997 26556 14044 26560
rect 14108 26558 14154 26618
rect 14825 26616 15351 26618
rect 14825 26560 14830 26616
rect 14886 26560 15290 26616
rect 15346 26560 15351 26616
rect 14825 26558 15351 26560
rect 14108 26556 14114 26558
rect 13997 26555 14063 26556
rect 14825 26555 14891 26558
rect 15285 26555 15351 26558
rect 20437 26618 20503 26621
rect 21633 26618 21699 26621
rect 20437 26616 21699 26618
rect 20437 26560 20442 26616
rect 20498 26560 21638 26616
rect 21694 26560 21699 26616
rect 20437 26558 21699 26560
rect 20437 26555 20503 26558
rect 21633 26555 21699 26558
rect 6637 26484 6703 26485
rect 6637 26480 6684 26484
rect 6748 26482 6754 26484
rect 9121 26482 9187 26485
rect 25681 26482 25747 26485
rect 6637 26424 6642 26480
rect 6637 26420 6684 26424
rect 6748 26422 6794 26482
rect 9121 26480 25747 26482
rect 9121 26424 9126 26480
rect 9182 26424 25686 26480
rect 25742 26424 25747 26480
rect 9121 26422 25747 26424
rect 6748 26420 6754 26422
rect 6637 26419 6703 26420
rect 9121 26419 9187 26422
rect 25681 26419 25747 26422
rect 5257 26348 5323 26349
rect 5206 26284 5212 26348
rect 5276 26346 5323 26348
rect 8937 26346 9003 26349
rect 9254 26346 9260 26348
rect 5276 26344 5368 26346
rect 5318 26288 5368 26344
rect 5276 26286 5368 26288
rect 8937 26344 9260 26346
rect 8937 26288 8942 26344
rect 8998 26288 9260 26344
rect 8937 26286 9260 26288
rect 5276 26284 5323 26286
rect 5257 26283 5323 26284
rect 8937 26283 9003 26286
rect 9254 26284 9260 26286
rect 9324 26284 9330 26348
rect 23197 26346 23263 26349
rect 9630 26344 23263 26346
rect 9630 26288 23202 26344
rect 23258 26288 23263 26344
rect 9630 26286 23263 26288
rect 0 26210 400 26240
rect 3785 26210 3851 26213
rect 0 26208 3851 26210
rect 0 26152 3790 26208
rect 3846 26152 3851 26208
rect 0 26150 3851 26152
rect 0 26120 400 26150
rect 3785 26147 3851 26150
rect 8334 26148 8340 26212
rect 8404 26210 8410 26212
rect 9630 26210 9690 26286
rect 23197 26283 23263 26286
rect 8404 26150 9690 26210
rect 8404 26148 8410 26150
rect 10358 26148 10364 26212
rect 10428 26210 10434 26212
rect 10501 26210 10567 26213
rect 14641 26210 14707 26213
rect 10428 26208 10567 26210
rect 10428 26152 10506 26208
rect 10562 26152 10567 26208
rect 10428 26150 10567 26152
rect 10428 26148 10434 26150
rect 10501 26147 10567 26150
rect 12390 26208 14707 26210
rect 12390 26152 14646 26208
rect 14702 26152 14707 26208
rect 12390 26150 14707 26152
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 4102 26012 4108 26076
rect 4172 26074 4178 26076
rect 4797 26074 4863 26077
rect 4172 26072 4863 26074
rect 4172 26016 4802 26072
rect 4858 26016 4863 26072
rect 4172 26014 4863 26016
rect 4172 26012 4178 26014
rect 4797 26011 4863 26014
rect 8753 26074 8819 26077
rect 12390 26074 12450 26150
rect 14641 26147 14707 26150
rect 15285 26210 15351 26213
rect 21633 26210 21699 26213
rect 15285 26208 21699 26210
rect 15285 26152 15290 26208
rect 15346 26152 21638 26208
rect 21694 26152 21699 26208
rect 15285 26150 21699 26152
rect 15285 26147 15351 26150
rect 21633 26147 21699 26150
rect 22185 26210 22251 26213
rect 22318 26210 22324 26212
rect 22185 26208 22324 26210
rect 22185 26152 22190 26208
rect 22246 26152 22324 26208
rect 22185 26150 22324 26152
rect 22185 26147 22251 26150
rect 22318 26148 22324 26150
rect 22388 26148 22394 26212
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 8753 26072 12450 26074
rect 8753 26016 8758 26072
rect 8814 26016 12450 26072
rect 8753 26014 12450 26016
rect 8753 26011 8819 26014
rect 17902 26012 17908 26076
rect 17972 26074 17978 26076
rect 17972 26014 19626 26074
rect 17972 26012 17978 26014
rect 3417 25938 3483 25941
rect 19374 25938 19380 25940
rect 3417 25936 19380 25938
rect 3417 25880 3422 25936
rect 3478 25880 19380 25936
rect 3417 25878 19380 25880
rect 3417 25875 3483 25878
rect 19374 25876 19380 25878
rect 19444 25876 19450 25940
rect 19566 25938 19626 26014
rect 25681 25938 25747 25941
rect 19566 25936 25747 25938
rect 19566 25880 25686 25936
rect 25742 25880 25747 25936
rect 19566 25878 25747 25880
rect 25681 25875 25747 25878
rect 9765 25804 9831 25805
rect 9765 25802 9812 25804
rect 9720 25800 9812 25802
rect 9876 25802 9882 25804
rect 14549 25802 14615 25805
rect 9876 25800 14615 25802
rect 9720 25744 9770 25800
rect 9876 25744 14554 25800
rect 14610 25744 14615 25800
rect 9720 25742 9812 25744
rect 9765 25740 9812 25742
rect 9876 25742 14615 25744
rect 9876 25740 9882 25742
rect 9765 25739 9831 25740
rect 14549 25739 14615 25742
rect 14733 25802 14799 25805
rect 25865 25802 25931 25805
rect 14733 25800 25931 25802
rect 14733 25744 14738 25800
rect 14794 25744 25870 25800
rect 25926 25744 25931 25800
rect 14733 25742 25931 25744
rect 14733 25739 14799 25742
rect 25865 25739 25931 25742
rect 7598 25604 7604 25668
rect 7668 25666 7674 25668
rect 8109 25666 8175 25669
rect 7668 25664 8175 25666
rect 7668 25608 8114 25664
rect 8170 25608 8175 25664
rect 7668 25606 8175 25608
rect 7668 25604 7674 25606
rect 8109 25603 8175 25606
rect 10501 25666 10567 25669
rect 11053 25666 11119 25669
rect 10501 25664 11119 25666
rect 10501 25608 10506 25664
rect 10562 25608 11058 25664
rect 11114 25608 11119 25664
rect 10501 25606 11119 25608
rect 10501 25603 10567 25606
rect 11053 25603 11119 25606
rect 18822 25604 18828 25668
rect 18892 25666 18898 25668
rect 20713 25666 20779 25669
rect 18892 25664 20779 25666
rect 18892 25608 20718 25664
rect 20774 25608 20779 25664
rect 18892 25606 20779 25608
rect 18892 25604 18898 25606
rect 20713 25603 20779 25606
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 7557 25530 7623 25533
rect 11053 25530 11119 25533
rect 7557 25528 11119 25530
rect 7557 25472 7562 25528
rect 7618 25472 11058 25528
rect 11114 25472 11119 25528
rect 7557 25470 11119 25472
rect 7557 25467 7623 25470
rect 11053 25467 11119 25470
rect 13905 25530 13971 25533
rect 14590 25530 14596 25532
rect 13905 25528 14596 25530
rect 13905 25472 13910 25528
rect 13966 25472 14596 25528
rect 13905 25470 14596 25472
rect 13905 25467 13971 25470
rect 14590 25468 14596 25470
rect 14660 25530 14666 25532
rect 15009 25530 15075 25533
rect 14660 25528 15075 25530
rect 14660 25472 15014 25528
rect 15070 25472 15075 25528
rect 14660 25470 15075 25472
rect 14660 25468 14666 25470
rect 15009 25467 15075 25470
rect 20713 25530 20779 25533
rect 23289 25530 23355 25533
rect 20713 25528 23355 25530
rect 20713 25472 20718 25528
rect 20774 25472 23294 25528
rect 23350 25472 23355 25528
rect 20713 25470 23355 25472
rect 20713 25467 20779 25470
rect 23289 25467 23355 25470
rect 3182 25332 3188 25396
rect 3252 25394 3258 25396
rect 6545 25394 6611 25397
rect 3252 25392 6611 25394
rect 3252 25336 6550 25392
rect 6606 25336 6611 25392
rect 3252 25334 6611 25336
rect 3252 25332 3258 25334
rect 6545 25331 6611 25334
rect 7281 25394 7347 25397
rect 27981 25394 28047 25397
rect 7281 25392 28047 25394
rect 7281 25336 7286 25392
rect 7342 25336 27986 25392
rect 28042 25336 28047 25392
rect 7281 25334 28047 25336
rect 7281 25331 7347 25334
rect 27981 25331 28047 25334
rect 4889 25258 4955 25261
rect 6545 25258 6611 25261
rect 4889 25256 6611 25258
rect 4889 25200 4894 25256
rect 4950 25200 6550 25256
rect 6606 25200 6611 25256
rect 4889 25198 6611 25200
rect 4889 25195 4955 25198
rect 6545 25195 6611 25198
rect 6821 25256 6887 25261
rect 6821 25200 6826 25256
rect 6882 25200 6887 25256
rect 6821 25195 6887 25200
rect 7649 25258 7715 25261
rect 14549 25258 14615 25261
rect 22318 25258 22324 25260
rect 7649 25256 9690 25258
rect 7649 25200 7654 25256
rect 7710 25200 9690 25256
rect 7649 25198 9690 25200
rect 7649 25195 7715 25198
rect 2221 25122 2287 25125
rect 6824 25122 6884 25195
rect 7281 25122 7347 25125
rect 2221 25120 7347 25122
rect 2221 25064 2226 25120
rect 2282 25064 7286 25120
rect 7342 25064 7347 25120
rect 2221 25062 7347 25064
rect 9630 25122 9690 25198
rect 14549 25256 22324 25258
rect 14549 25200 14554 25256
rect 14610 25200 22324 25256
rect 14549 25198 22324 25200
rect 14549 25195 14615 25198
rect 22318 25196 22324 25198
rect 22388 25196 22394 25260
rect 14549 25122 14615 25125
rect 9630 25120 14615 25122
rect 9630 25064 14554 25120
rect 14610 25064 14615 25120
rect 9630 25062 14615 25064
rect 2221 25059 2287 25062
rect 7281 25059 7347 25062
rect 14549 25059 14615 25062
rect 15326 25060 15332 25124
rect 15396 25122 15402 25124
rect 16297 25122 16363 25125
rect 15396 25120 16363 25122
rect 15396 25064 16302 25120
rect 16358 25064 16363 25120
rect 15396 25062 16363 25064
rect 15396 25060 15402 25062
rect 16297 25059 16363 25062
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 5349 24988 5415 24989
rect 13169 24988 13235 24989
rect 5349 24984 5396 24988
rect 5460 24986 5466 24988
rect 5349 24928 5354 24984
rect 5349 24924 5396 24928
rect 5460 24926 5506 24986
rect 5460 24924 5466 24926
rect 13118 24924 13124 24988
rect 13188 24986 13235 24988
rect 15837 24986 15903 24989
rect 16062 24986 16068 24988
rect 13188 24984 13280 24986
rect 13230 24928 13280 24984
rect 13188 24926 13280 24928
rect 15837 24984 16068 24986
rect 15837 24928 15842 24984
rect 15898 24928 16068 24984
rect 15837 24926 16068 24928
rect 13188 24924 13235 24926
rect 5349 24923 5415 24924
rect 13169 24923 13235 24924
rect 15837 24923 15903 24926
rect 16062 24924 16068 24926
rect 16132 24924 16138 24988
rect 16941 24986 17007 24989
rect 18822 24986 18828 24988
rect 16941 24984 18828 24986
rect 16941 24928 16946 24984
rect 17002 24928 18828 24984
rect 16941 24926 18828 24928
rect 16941 24923 17007 24926
rect 18822 24924 18828 24926
rect 18892 24924 18898 24988
rect 5809 24850 5875 24853
rect 23841 24850 23907 24853
rect 5809 24848 23907 24850
rect 5809 24792 5814 24848
rect 5870 24792 23846 24848
rect 23902 24792 23907 24848
rect 5809 24790 23907 24792
rect 5809 24787 5875 24790
rect 23841 24787 23907 24790
rect 4797 24714 4863 24717
rect 7925 24714 7991 24717
rect 4797 24712 7991 24714
rect 4797 24656 4802 24712
rect 4858 24656 7930 24712
rect 7986 24656 7991 24712
rect 4797 24654 7991 24656
rect 4797 24651 4863 24654
rect 7925 24651 7991 24654
rect 11513 24714 11579 24717
rect 11513 24712 12450 24714
rect 11513 24656 11518 24712
rect 11574 24656 12450 24712
rect 11513 24654 12450 24656
rect 11513 24651 11579 24654
rect 12390 24578 12450 24654
rect 15878 24652 15884 24716
rect 15948 24714 15954 24716
rect 16021 24714 16087 24717
rect 23381 24714 23447 24717
rect 15948 24712 16087 24714
rect 15948 24656 16026 24712
rect 16082 24656 16087 24712
rect 15948 24654 16087 24656
rect 15948 24652 15954 24654
rect 16021 24651 16087 24654
rect 17174 24712 23447 24714
rect 17174 24656 23386 24712
rect 23442 24656 23447 24712
rect 17174 24654 23447 24656
rect 17174 24578 17234 24654
rect 23381 24651 23447 24654
rect 12390 24518 17234 24578
rect 19333 24578 19399 24581
rect 22645 24578 22711 24581
rect 19333 24576 22711 24578
rect 19333 24520 19338 24576
rect 19394 24520 22650 24576
rect 22706 24520 22711 24576
rect 19333 24518 22711 24520
rect 19333 24515 19399 24518
rect 22645 24515 22711 24518
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 13353 24442 13419 24445
rect 15009 24442 15075 24445
rect 13353 24440 15075 24442
rect 13353 24384 13358 24440
rect 13414 24384 15014 24440
rect 15070 24384 15075 24440
rect 13353 24382 15075 24384
rect 13353 24379 13419 24382
rect 15009 24379 15075 24382
rect 8753 24306 8819 24309
rect 17309 24306 17375 24309
rect 23105 24306 23171 24309
rect 8753 24304 17234 24306
rect 8753 24248 8758 24304
rect 8814 24248 17234 24304
rect 8753 24246 17234 24248
rect 8753 24243 8819 24246
rect 0 24170 400 24200
rect 3969 24170 4035 24173
rect 0 24168 4035 24170
rect 0 24112 3974 24168
rect 4030 24112 4035 24168
rect 0 24110 4035 24112
rect 0 24080 400 24110
rect 3969 24107 4035 24110
rect 5533 24170 5599 24173
rect 7005 24170 7071 24173
rect 5533 24168 7071 24170
rect 5533 24112 5538 24168
rect 5594 24112 7010 24168
rect 7066 24112 7071 24168
rect 5533 24110 7071 24112
rect 5533 24107 5599 24110
rect 7005 24107 7071 24110
rect 9581 24170 9647 24173
rect 17174 24170 17234 24246
rect 17309 24304 23171 24306
rect 17309 24248 17314 24304
rect 17370 24248 23110 24304
rect 23166 24248 23171 24304
rect 17309 24246 23171 24248
rect 17309 24243 17375 24246
rect 23105 24243 23171 24246
rect 25037 24170 25103 24173
rect 9581 24168 13738 24170
rect 9581 24112 9586 24168
rect 9642 24112 13738 24168
rect 9581 24110 13738 24112
rect 9581 24107 9647 24110
rect 6310 23972 6316 24036
rect 6380 24034 6386 24036
rect 6453 24034 6519 24037
rect 6380 24032 6519 24034
rect 6380 23976 6458 24032
rect 6514 23976 6519 24032
rect 6380 23974 6519 23976
rect 6380 23972 6386 23974
rect 6453 23971 6519 23974
rect 10358 23972 10364 24036
rect 10428 24034 10434 24036
rect 10501 24034 10567 24037
rect 10428 24032 10567 24034
rect 10428 23976 10506 24032
rect 10562 23976 10567 24032
rect 10428 23974 10567 23976
rect 10428 23972 10434 23974
rect 10501 23971 10567 23974
rect 11605 24034 11671 24037
rect 13118 24034 13124 24036
rect 11605 24032 13124 24034
rect 11605 23976 11610 24032
rect 11666 23976 13124 24032
rect 11605 23974 13124 23976
rect 11605 23971 11671 23974
rect 13118 23972 13124 23974
rect 13188 23972 13194 24036
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 6913 23898 6979 23901
rect 7046 23898 7052 23900
rect 6913 23896 7052 23898
rect 6913 23840 6918 23896
rect 6974 23840 7052 23896
rect 6913 23838 7052 23840
rect 6913 23835 6979 23838
rect 7046 23836 7052 23838
rect 7116 23836 7122 23900
rect 10041 23898 10107 23901
rect 12014 23898 12020 23900
rect 10041 23896 12020 23898
rect 10041 23840 10046 23896
rect 10102 23840 12020 23896
rect 10041 23838 12020 23840
rect 10041 23835 10107 23838
rect 12014 23836 12020 23838
rect 12084 23898 12090 23900
rect 13261 23898 13327 23901
rect 12084 23896 13327 23898
rect 12084 23840 13266 23896
rect 13322 23840 13327 23896
rect 12084 23838 13327 23840
rect 13678 23898 13738 24110
rect 14230 24110 16314 24170
rect 17174 24168 25103 24170
rect 17174 24112 25042 24168
rect 25098 24112 25103 24168
rect 17174 24110 25103 24112
rect 14230 23898 14290 24110
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 13678 23838 14290 23898
rect 16254 23898 16314 24110
rect 25037 24107 25103 24110
rect 16481 24034 16547 24037
rect 17309 24034 17375 24037
rect 19057 24036 19123 24037
rect 16481 24032 17375 24034
rect 16481 23976 16486 24032
rect 16542 23976 17314 24032
rect 17370 23976 17375 24032
rect 16481 23974 17375 23976
rect 16481 23971 16547 23974
rect 17309 23971 17375 23974
rect 19006 23972 19012 24036
rect 19076 24034 19123 24036
rect 19076 24032 19168 24034
rect 19118 23976 19168 24032
rect 19076 23974 19168 23976
rect 19076 23972 19123 23974
rect 19057 23971 19123 23972
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 21173 23898 21239 23901
rect 16254 23896 21239 23898
rect 16254 23840 21178 23896
rect 21234 23840 21239 23896
rect 16254 23838 21239 23840
rect 12084 23836 12090 23838
rect 13261 23835 13327 23838
rect 21173 23835 21239 23838
rect 1761 23762 1827 23765
rect 24669 23762 24735 23765
rect 1761 23760 24735 23762
rect 1761 23704 1766 23760
rect 1822 23704 24674 23760
rect 24730 23704 24735 23760
rect 1761 23702 24735 23704
rect 1761 23699 1827 23702
rect 24669 23699 24735 23702
rect 4337 23628 4403 23629
rect 4286 23626 4292 23628
rect 4246 23566 4292 23626
rect 4356 23624 4403 23628
rect 4398 23568 4403 23624
rect 4286 23564 4292 23566
rect 4356 23564 4403 23568
rect 4337 23563 4403 23564
rect 7005 23626 7071 23629
rect 8334 23626 8340 23628
rect 7005 23624 8340 23626
rect 7005 23568 7010 23624
rect 7066 23568 8340 23624
rect 7005 23566 8340 23568
rect 7005 23563 7071 23566
rect 8334 23564 8340 23566
rect 8404 23564 8410 23628
rect 9438 23564 9444 23628
rect 9508 23626 9514 23628
rect 14273 23626 14339 23629
rect 9508 23624 14339 23626
rect 9508 23568 14278 23624
rect 14334 23568 14339 23624
rect 9508 23566 14339 23568
rect 9508 23564 9514 23566
rect 14273 23563 14339 23566
rect 14457 23626 14523 23629
rect 15929 23626 15995 23629
rect 14457 23624 15995 23626
rect 14457 23568 14462 23624
rect 14518 23568 15934 23624
rect 15990 23568 15995 23624
rect 14457 23566 15995 23568
rect 14457 23563 14523 23566
rect 15929 23563 15995 23566
rect 16297 23626 16363 23629
rect 17677 23626 17743 23629
rect 16297 23624 17743 23626
rect 16297 23568 16302 23624
rect 16358 23568 17682 23624
rect 17738 23568 17743 23624
rect 16297 23566 17743 23568
rect 16297 23563 16363 23566
rect 17677 23563 17743 23566
rect 18965 23626 19031 23629
rect 23657 23626 23723 23629
rect 18965 23624 23723 23626
rect 18965 23568 18970 23624
rect 19026 23568 23662 23624
rect 23718 23568 23723 23624
rect 18965 23566 23723 23568
rect 18965 23563 19031 23566
rect 23657 23563 23723 23566
rect 5809 23490 5875 23493
rect 8569 23490 8635 23493
rect 5809 23488 8635 23490
rect 5809 23432 5814 23488
rect 5870 23432 8574 23488
rect 8630 23432 8635 23488
rect 5809 23430 8635 23432
rect 5809 23427 5875 23430
rect 8569 23427 8635 23430
rect 14825 23490 14891 23493
rect 16573 23490 16639 23493
rect 14825 23488 16639 23490
rect 14825 23432 14830 23488
rect 14886 23432 16578 23488
rect 16634 23432 16639 23488
rect 14825 23430 16639 23432
rect 14825 23427 14891 23430
rect 16573 23427 16639 23430
rect 19701 23490 19767 23493
rect 19701 23488 25146 23490
rect 19701 23432 19706 23488
rect 19762 23432 25146 23488
rect 19701 23430 25146 23432
rect 19701 23427 19767 23430
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 4889 23354 4955 23357
rect 5717 23354 5783 23357
rect 4889 23352 5783 23354
rect 4889 23296 4894 23352
rect 4950 23296 5722 23352
rect 5778 23296 5783 23352
rect 4889 23294 5783 23296
rect 4889 23291 4955 23294
rect 5717 23291 5783 23294
rect 9305 23354 9371 23357
rect 11789 23354 11855 23357
rect 17125 23354 17191 23357
rect 9305 23352 10794 23354
rect 9305 23296 9310 23352
rect 9366 23296 10794 23352
rect 9305 23294 10794 23296
rect 9305 23291 9371 23294
rect 5717 23218 5783 23221
rect 8477 23218 8543 23221
rect 10501 23220 10567 23221
rect 10501 23218 10548 23220
rect 5717 23216 8543 23218
rect 5717 23160 5722 23216
rect 5778 23160 8482 23216
rect 8538 23160 8543 23216
rect 5717 23158 8543 23160
rect 10456 23216 10548 23218
rect 10456 23160 10506 23216
rect 10456 23158 10548 23160
rect 5717 23155 5783 23158
rect 8477 23155 8543 23158
rect 10501 23156 10548 23158
rect 10612 23156 10618 23220
rect 10734 23218 10794 23294
rect 11789 23352 17191 23354
rect 11789 23296 11794 23352
rect 11850 23296 17130 23352
rect 17186 23296 17191 23352
rect 11789 23294 17191 23296
rect 11789 23291 11855 23294
rect 17125 23291 17191 23294
rect 18689 23354 18755 23357
rect 22737 23354 22803 23357
rect 18689 23352 22803 23354
rect 18689 23296 18694 23352
rect 18750 23296 22742 23352
rect 22798 23296 22803 23352
rect 18689 23294 22803 23296
rect 18689 23291 18755 23294
rect 22737 23291 22803 23294
rect 23013 23354 23079 23357
rect 24117 23354 24183 23357
rect 23013 23352 24183 23354
rect 23013 23296 23018 23352
rect 23074 23296 24122 23352
rect 24178 23296 24183 23352
rect 23013 23294 24183 23296
rect 23013 23291 23079 23294
rect 24117 23291 24183 23294
rect 24577 23218 24643 23221
rect 10734 23216 24643 23218
rect 10734 23160 24582 23216
rect 24638 23160 24643 23216
rect 10734 23158 24643 23160
rect 25086 23218 25146 23430
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 25681 23218 25747 23221
rect 25086 23216 25747 23218
rect 25086 23160 25686 23216
rect 25742 23160 25747 23216
rect 25086 23158 25747 23160
rect 10501 23155 10567 23156
rect 24577 23155 24643 23158
rect 25681 23155 25747 23158
rect 2957 23082 3023 23085
rect 6678 23082 6684 23084
rect 2957 23080 6684 23082
rect 2957 23024 2962 23080
rect 3018 23024 6684 23080
rect 2957 23022 6684 23024
rect 2957 23019 3023 23022
rect 6678 23020 6684 23022
rect 6748 23020 6754 23084
rect 9121 23082 9187 23085
rect 24301 23082 24367 23085
rect 9121 23080 24367 23082
rect 9121 23024 9126 23080
rect 9182 23024 24306 23080
rect 24362 23024 24367 23080
rect 9121 23022 24367 23024
rect 9121 23019 9187 23022
rect 24301 23019 24367 23022
rect 16430 22884 16436 22948
rect 16500 22946 16506 22948
rect 18597 22946 18663 22949
rect 16500 22944 18663 22946
rect 16500 22888 18602 22944
rect 18658 22888 18663 22944
rect 16500 22886 18663 22888
rect 16500 22884 16506 22886
rect 18597 22883 18663 22886
rect 19374 22884 19380 22948
rect 19444 22946 19450 22948
rect 19701 22946 19767 22949
rect 19444 22944 19767 22946
rect 19444 22888 19706 22944
rect 19762 22888 19767 22944
rect 19444 22886 19767 22888
rect 19444 22884 19450 22886
rect 19701 22883 19767 22886
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 2681 22810 2747 22813
rect 4889 22810 4955 22813
rect 2681 22808 4955 22810
rect 2681 22752 2686 22808
rect 2742 22752 4894 22808
rect 4950 22752 4955 22808
rect 2681 22750 4955 22752
rect 2681 22747 2747 22750
rect 4889 22747 4955 22750
rect 16021 22810 16087 22813
rect 20253 22810 20319 22813
rect 16021 22808 20319 22810
rect 16021 22752 16026 22808
rect 16082 22752 20258 22808
rect 20314 22752 20319 22808
rect 16021 22750 20319 22752
rect 16021 22747 16087 22750
rect 20253 22747 20319 22750
rect 3233 22674 3299 22677
rect 5574 22674 5580 22676
rect 3233 22672 5580 22674
rect 3233 22616 3238 22672
rect 3294 22616 5580 22672
rect 3233 22614 5580 22616
rect 3233 22611 3299 22614
rect 5574 22612 5580 22614
rect 5644 22674 5650 22676
rect 9305 22674 9371 22677
rect 5644 22672 9371 22674
rect 5644 22616 9310 22672
rect 9366 22616 9371 22672
rect 5644 22614 9371 22616
rect 5644 22612 5650 22614
rect 9305 22611 9371 22614
rect 13905 22674 13971 22677
rect 17350 22674 17356 22676
rect 13905 22672 17356 22674
rect 13905 22616 13910 22672
rect 13966 22616 17356 22672
rect 13905 22614 17356 22616
rect 13905 22611 13971 22614
rect 17350 22612 17356 22614
rect 17420 22612 17426 22676
rect 18086 22612 18092 22676
rect 18156 22674 18162 22676
rect 19977 22674 20043 22677
rect 18156 22672 20043 22674
rect 18156 22616 19982 22672
rect 20038 22616 20043 22672
rect 18156 22614 20043 22616
rect 18156 22612 18162 22614
rect 19977 22611 20043 22614
rect 2589 22538 2655 22541
rect 4613 22538 4679 22541
rect 2589 22536 4679 22538
rect 2589 22480 2594 22536
rect 2650 22480 4618 22536
rect 4674 22480 4679 22536
rect 2589 22478 4679 22480
rect 2589 22475 2655 22478
rect 4613 22475 4679 22478
rect 7598 22476 7604 22540
rect 7668 22538 7674 22540
rect 24669 22538 24735 22541
rect 7668 22536 24735 22538
rect 7668 22480 24674 22536
rect 24730 22480 24735 22536
rect 7668 22478 24735 22480
rect 7668 22476 7674 22478
rect 24669 22475 24735 22478
rect 5349 22402 5415 22405
rect 6361 22402 6427 22405
rect 5349 22400 6427 22402
rect 5349 22344 5354 22400
rect 5410 22344 6366 22400
rect 6422 22344 6427 22400
rect 5349 22342 6427 22344
rect 5349 22339 5415 22342
rect 6361 22339 6427 22342
rect 19057 22402 19123 22405
rect 19190 22402 19196 22404
rect 19057 22400 19196 22402
rect 19057 22344 19062 22400
rect 19118 22344 19196 22400
rect 19057 22342 19196 22344
rect 19057 22339 19123 22342
rect 19190 22340 19196 22342
rect 19260 22340 19266 22404
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 2129 22266 2195 22269
rect 3233 22266 3299 22269
rect 2129 22264 3299 22266
rect 2129 22208 2134 22264
rect 2190 22208 3238 22264
rect 3294 22208 3299 22264
rect 2129 22206 3299 22208
rect 2129 22203 2195 22206
rect 3233 22203 3299 22206
rect 14590 22204 14596 22268
rect 14660 22266 14666 22268
rect 15009 22266 15075 22269
rect 14660 22264 15075 22266
rect 14660 22208 15014 22264
rect 15070 22208 15075 22264
rect 14660 22206 15075 22208
rect 14660 22204 14666 22206
rect 15009 22203 15075 22206
rect 19425 22266 19491 22269
rect 22553 22266 22619 22269
rect 19425 22264 22619 22266
rect 19425 22208 19430 22264
rect 19486 22208 22558 22264
rect 22614 22208 22619 22264
rect 19425 22206 22619 22208
rect 19425 22203 19491 22206
rect 22553 22203 22619 22206
rect 0 22130 400 22160
rect 473 22130 539 22133
rect 0 22128 539 22130
rect 0 22072 478 22128
rect 534 22072 539 22128
rect 0 22070 539 22072
rect 0 22040 400 22070
rect 473 22067 539 22070
rect 1853 22130 1919 22133
rect 2865 22130 2931 22133
rect 5717 22130 5783 22133
rect 1853 22128 5783 22130
rect 1853 22072 1858 22128
rect 1914 22072 2870 22128
rect 2926 22072 5722 22128
rect 5778 22072 5783 22128
rect 1853 22070 5783 22072
rect 1853 22067 1919 22070
rect 2865 22067 2931 22070
rect 5717 22067 5783 22070
rect 7005 22130 7071 22133
rect 9397 22130 9463 22133
rect 7005 22128 9463 22130
rect 7005 22072 7010 22128
rect 7066 22072 9402 22128
rect 9458 22072 9463 22128
rect 7005 22070 9463 22072
rect 7005 22067 7071 22070
rect 9397 22067 9463 22070
rect 13721 22130 13787 22133
rect 17309 22130 17375 22133
rect 13721 22128 17375 22130
rect 13721 22072 13726 22128
rect 13782 22072 17314 22128
rect 17370 22072 17375 22128
rect 13721 22070 17375 22072
rect 13721 22067 13787 22070
rect 17309 22067 17375 22070
rect 17769 22130 17835 22133
rect 18229 22130 18295 22133
rect 17769 22128 18295 22130
rect 17769 22072 17774 22128
rect 17830 22072 18234 22128
rect 18290 22072 18295 22128
rect 17769 22070 18295 22072
rect 17769 22067 17835 22070
rect 18229 22067 18295 22070
rect 19885 22130 19951 22133
rect 20529 22130 20595 22133
rect 26601 22130 26667 22133
rect 19885 22128 26667 22130
rect 19885 22072 19890 22128
rect 19946 22072 20534 22128
rect 20590 22072 26606 22128
rect 26662 22072 26667 22128
rect 19885 22070 26667 22072
rect 19885 22067 19951 22070
rect 20529 22067 20595 22070
rect 26601 22067 26667 22070
rect 2773 21994 2839 21997
rect 3049 21994 3115 21997
rect 6269 21994 6335 21997
rect 2773 21992 6335 21994
rect 2773 21936 2778 21992
rect 2834 21936 3054 21992
rect 3110 21936 6274 21992
rect 6330 21936 6335 21992
rect 2773 21934 6335 21936
rect 2773 21931 2839 21934
rect 3049 21931 3115 21934
rect 6269 21931 6335 21934
rect 16062 21932 16068 21996
rect 16132 21994 16138 21996
rect 20161 21994 20227 21997
rect 16132 21992 20227 21994
rect 16132 21936 20166 21992
rect 20222 21936 20227 21992
rect 16132 21934 20227 21936
rect 16132 21932 16138 21934
rect 20161 21931 20227 21934
rect 20897 21994 20963 21997
rect 27429 21994 27495 21997
rect 20897 21992 27495 21994
rect 20897 21936 20902 21992
rect 20958 21936 27434 21992
rect 27490 21936 27495 21992
rect 20897 21934 27495 21936
rect 20897 21931 20963 21934
rect 27429 21931 27495 21934
rect 1485 21858 1551 21861
rect 5533 21858 5599 21861
rect 6310 21858 6316 21860
rect 1485 21856 6316 21858
rect 1485 21800 1490 21856
rect 1546 21800 5538 21856
rect 5594 21800 6316 21856
rect 1485 21798 6316 21800
rect 1485 21795 1551 21798
rect 5533 21795 5599 21798
rect 6310 21796 6316 21798
rect 6380 21858 6386 21860
rect 7373 21858 7439 21861
rect 6380 21856 7439 21858
rect 6380 21800 7378 21856
rect 7434 21800 7439 21856
rect 6380 21798 7439 21800
rect 6380 21796 6386 21798
rect 7373 21795 7439 21798
rect 18321 21858 18387 21861
rect 20069 21858 20135 21861
rect 18321 21856 20135 21858
rect 18321 21800 18326 21856
rect 18382 21800 20074 21856
rect 20130 21800 20135 21856
rect 18321 21798 20135 21800
rect 18321 21795 18387 21798
rect 20069 21795 20135 21798
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 9949 21722 10015 21725
rect 10777 21722 10843 21725
rect 9949 21720 10843 21722
rect 9949 21664 9954 21720
rect 10010 21664 10782 21720
rect 10838 21664 10843 21720
rect 9949 21662 10843 21664
rect 9949 21659 10015 21662
rect 10777 21659 10843 21662
rect 18873 21722 18939 21725
rect 19006 21722 19012 21724
rect 18873 21720 19012 21722
rect 18873 21664 18878 21720
rect 18934 21664 19012 21720
rect 18873 21662 19012 21664
rect 18873 21659 18939 21662
rect 19006 21660 19012 21662
rect 19076 21660 19082 21724
rect 2497 21586 2563 21589
rect 3049 21586 3115 21589
rect 3182 21586 3188 21588
rect 2497 21584 2790 21586
rect 2497 21528 2502 21584
rect 2558 21528 2790 21584
rect 2497 21526 2790 21528
rect 2497 21523 2563 21526
rect 2730 21450 2790 21526
rect 3049 21584 3188 21586
rect 3049 21528 3054 21584
rect 3110 21528 3188 21584
rect 3049 21526 3188 21528
rect 3049 21523 3115 21526
rect 3182 21524 3188 21526
rect 3252 21524 3258 21588
rect 7097 21586 7163 21589
rect 23197 21586 23263 21589
rect 3374 21584 23263 21586
rect 3374 21528 7102 21584
rect 7158 21528 23202 21584
rect 23258 21528 23263 21584
rect 3374 21526 23263 21528
rect 3374 21450 3434 21526
rect 7097 21523 7163 21526
rect 23197 21523 23263 21526
rect 2730 21390 3434 21450
rect 5349 21448 5415 21453
rect 5349 21392 5354 21448
rect 5410 21392 5415 21448
rect 5349 21387 5415 21392
rect 9397 21450 9463 21453
rect 14089 21450 14155 21453
rect 15326 21450 15332 21452
rect 9397 21448 15332 21450
rect 9397 21392 9402 21448
rect 9458 21392 14094 21448
rect 14150 21392 15332 21448
rect 9397 21390 15332 21392
rect 9397 21387 9463 21390
rect 14089 21387 14155 21390
rect 15326 21388 15332 21390
rect 15396 21388 15402 21452
rect 18413 21450 18479 21453
rect 18822 21450 18828 21452
rect 18413 21448 18828 21450
rect 18413 21392 18418 21448
rect 18474 21392 18828 21448
rect 18413 21390 18828 21392
rect 18413 21387 18479 21390
rect 18822 21388 18828 21390
rect 18892 21388 18898 21452
rect 20294 21388 20300 21452
rect 20364 21450 20370 21452
rect 20437 21450 20503 21453
rect 20364 21448 20503 21450
rect 20364 21392 20442 21448
rect 20498 21392 20503 21448
rect 20364 21390 20503 21392
rect 20364 21388 20370 21390
rect 20437 21387 20503 21390
rect 5352 21314 5412 21387
rect 5352 21254 5642 21314
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 5206 21116 5212 21180
rect 5276 21178 5282 21180
rect 5441 21178 5507 21181
rect 5276 21176 5507 21178
rect 5276 21120 5446 21176
rect 5502 21120 5507 21176
rect 5276 21118 5507 21120
rect 5276 21116 5282 21118
rect 5441 21115 5507 21118
rect 5165 21044 5231 21045
rect 5165 21042 5212 21044
rect 5120 21040 5212 21042
rect 5120 20984 5170 21040
rect 5120 20982 5212 20984
rect 5165 20980 5212 20982
rect 5276 20980 5282 21044
rect 5349 21042 5415 21045
rect 5582 21042 5642 21254
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 6637 21044 6703 21045
rect 6637 21042 6684 21044
rect 5349 21040 5642 21042
rect 5349 20984 5354 21040
rect 5410 20984 5642 21040
rect 5349 20982 5642 20984
rect 6592 21040 6684 21042
rect 6592 20984 6642 21040
rect 6592 20982 6684 20984
rect 5165 20979 5231 20980
rect 5349 20979 5415 20982
rect 6637 20980 6684 20982
rect 6748 20980 6754 21044
rect 19057 21042 19123 21045
rect 19190 21042 19196 21044
rect 19057 21040 19196 21042
rect 19057 20984 19062 21040
rect 19118 20984 19196 21040
rect 19057 20982 19196 20984
rect 6637 20979 6703 20980
rect 19057 20979 19123 20982
rect 19190 20980 19196 20982
rect 19260 20980 19266 21044
rect 21541 21042 21607 21045
rect 25865 21042 25931 21045
rect 21541 21040 25931 21042
rect 21541 20984 21546 21040
rect 21602 20984 25870 21040
rect 25926 20984 25931 21040
rect 21541 20982 25931 20984
rect 21541 20979 21607 20982
rect 25865 20979 25931 20982
rect 933 20906 999 20909
rect 2405 20906 2471 20909
rect 4429 20906 4495 20909
rect 933 20904 4495 20906
rect 933 20848 938 20904
rect 994 20848 2410 20904
rect 2466 20848 4434 20904
rect 4490 20848 4495 20904
rect 933 20846 4495 20848
rect 933 20843 999 20846
rect 2405 20843 2471 20846
rect 4429 20843 4495 20846
rect 10593 20906 10659 20909
rect 12433 20906 12499 20909
rect 10593 20904 12499 20906
rect 10593 20848 10598 20904
rect 10654 20848 12438 20904
rect 12494 20848 12499 20904
rect 10593 20846 12499 20848
rect 10593 20843 10659 20846
rect 12433 20843 12499 20846
rect 12709 20906 12775 20909
rect 22921 20906 22987 20909
rect 12709 20904 22987 20906
rect 12709 20848 12714 20904
rect 12770 20848 22926 20904
rect 22982 20848 22987 20904
rect 12709 20846 22987 20848
rect 12709 20843 12775 20846
rect 22921 20843 22987 20846
rect 8477 20772 8543 20773
rect 8477 20768 8524 20772
rect 8588 20770 8594 20772
rect 11421 20770 11487 20773
rect 12014 20770 12020 20772
rect 8477 20712 8482 20768
rect 8477 20708 8524 20712
rect 8588 20710 8634 20770
rect 11421 20768 12020 20770
rect 11421 20712 11426 20768
rect 11482 20712 12020 20768
rect 11421 20710 12020 20712
rect 8588 20708 8594 20710
rect 8477 20707 8543 20708
rect 11421 20707 11487 20710
rect 12014 20708 12020 20710
rect 12084 20708 12090 20772
rect 16941 20770 17007 20773
rect 17309 20770 17375 20773
rect 16941 20768 17375 20770
rect 16941 20712 16946 20768
rect 17002 20712 17314 20768
rect 17370 20712 17375 20768
rect 16941 20710 17375 20712
rect 16941 20707 17007 20710
rect 17309 20707 17375 20710
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 7005 20634 7071 20637
rect 3144 20632 7071 20634
rect 3144 20576 7010 20632
rect 7066 20576 7071 20632
rect 3144 20574 7071 20576
rect 3144 20501 3204 20574
rect 7005 20571 7071 20574
rect 19241 20634 19307 20637
rect 19374 20634 19380 20636
rect 19241 20632 19380 20634
rect 19241 20576 19246 20632
rect 19302 20576 19380 20632
rect 19241 20574 19380 20576
rect 19241 20571 19307 20574
rect 19374 20572 19380 20574
rect 19444 20572 19450 20636
rect 2497 20498 2563 20501
rect 3141 20498 3207 20501
rect 2497 20496 3207 20498
rect 2497 20440 2502 20496
rect 2558 20440 3146 20496
rect 3202 20440 3207 20496
rect 2497 20438 3207 20440
rect 2497 20435 2563 20438
rect 3141 20435 3207 20438
rect 4429 20498 4495 20501
rect 5073 20498 5139 20501
rect 5441 20498 5507 20501
rect 4429 20496 5507 20498
rect 4429 20440 4434 20496
rect 4490 20440 5078 20496
rect 5134 20440 5446 20496
rect 5502 20440 5507 20496
rect 4429 20438 5507 20440
rect 4429 20435 4495 20438
rect 5073 20435 5139 20438
rect 5441 20435 5507 20438
rect 9254 20436 9260 20500
rect 9324 20498 9330 20500
rect 13629 20498 13695 20501
rect 9324 20496 13695 20498
rect 9324 20440 13634 20496
rect 13690 20440 13695 20496
rect 9324 20438 13695 20440
rect 9324 20436 9330 20438
rect 13629 20435 13695 20438
rect 1158 20300 1164 20364
rect 1228 20362 1234 20364
rect 2129 20362 2195 20365
rect 5441 20362 5507 20365
rect 1228 20360 5507 20362
rect 1228 20304 2134 20360
rect 2190 20304 5446 20360
rect 5502 20304 5507 20360
rect 1228 20302 5507 20304
rect 1228 20300 1234 20302
rect 2129 20299 2195 20302
rect 5441 20299 5507 20302
rect 9765 20362 9831 20365
rect 13077 20362 13143 20365
rect 9765 20360 13143 20362
rect 9765 20304 9770 20360
rect 9826 20304 13082 20360
rect 13138 20304 13143 20360
rect 9765 20302 13143 20304
rect 9765 20299 9831 20302
rect 13077 20299 13143 20302
rect 17493 20362 17559 20365
rect 24301 20362 24367 20365
rect 17493 20360 24367 20362
rect 17493 20304 17498 20360
rect 17554 20304 24306 20360
rect 24362 20304 24367 20360
rect 17493 20302 24367 20304
rect 17493 20299 17559 20302
rect 24301 20299 24367 20302
rect 2221 20226 2287 20229
rect 4153 20228 4219 20229
rect 7097 20228 7163 20229
rect 4102 20226 4108 20228
rect 2221 20224 4108 20226
rect 4172 20226 4219 20228
rect 4172 20224 4264 20226
rect 2221 20168 2226 20224
rect 2282 20168 4108 20224
rect 4214 20168 4264 20224
rect 2221 20166 4108 20168
rect 2221 20163 2287 20166
rect 4102 20164 4108 20166
rect 4172 20166 4264 20168
rect 4172 20164 4219 20166
rect 7046 20164 7052 20228
rect 7116 20226 7163 20228
rect 13077 20226 13143 20229
rect 16021 20226 16087 20229
rect 7116 20224 7208 20226
rect 7158 20168 7208 20224
rect 7116 20166 7208 20168
rect 13077 20224 16087 20226
rect 13077 20168 13082 20224
rect 13138 20168 16026 20224
rect 16082 20168 16087 20224
rect 13077 20166 16087 20168
rect 7116 20164 7163 20166
rect 4153 20163 4219 20164
rect 7097 20163 7163 20164
rect 13077 20163 13143 20166
rect 16021 20163 16087 20166
rect 20478 20164 20484 20228
rect 20548 20226 20554 20228
rect 20621 20226 20687 20229
rect 20548 20224 20687 20226
rect 20548 20168 20626 20224
rect 20682 20168 20687 20224
rect 20548 20166 20687 20168
rect 20548 20164 20554 20166
rect 20621 20163 20687 20166
rect 4419 20160 4735 20161
rect 0 20090 400 20120
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 473 20090 539 20093
rect 9397 20090 9463 20093
rect 0 20088 539 20090
rect 0 20032 478 20088
rect 534 20032 539 20088
rect 0 20030 539 20032
rect 0 20000 400 20030
rect 473 20027 539 20030
rect 4846 20088 9463 20090
rect 4846 20032 9402 20088
rect 9458 20032 9463 20088
rect 4846 20030 9463 20032
rect 2865 19954 2931 19957
rect 3417 19954 3483 19957
rect 2865 19952 3483 19954
rect 2865 19896 2870 19952
rect 2926 19896 3422 19952
rect 3478 19896 3483 19952
rect 2865 19894 3483 19896
rect 2865 19891 2931 19894
rect 3417 19891 3483 19894
rect 3969 19954 4035 19957
rect 4846 19954 4906 20030
rect 9397 20027 9463 20030
rect 13670 20028 13676 20092
rect 13740 20090 13746 20092
rect 16205 20090 16271 20093
rect 13740 20088 16271 20090
rect 13740 20032 16210 20088
rect 16266 20032 16271 20088
rect 13740 20030 16271 20032
rect 13740 20028 13746 20030
rect 16205 20027 16271 20030
rect 3969 19952 4906 19954
rect 3969 19896 3974 19952
rect 4030 19896 4906 19952
rect 3969 19894 4906 19896
rect 3969 19891 4035 19894
rect 5390 19892 5396 19956
rect 5460 19954 5466 19956
rect 7649 19954 7715 19957
rect 5460 19952 7715 19954
rect 5460 19896 7654 19952
rect 7710 19896 7715 19952
rect 5460 19894 7715 19896
rect 5460 19892 5466 19894
rect 7649 19891 7715 19894
rect 14222 19892 14228 19956
rect 14292 19954 14298 19956
rect 14590 19954 14596 19956
rect 14292 19894 14596 19954
rect 14292 19892 14298 19894
rect 14590 19892 14596 19894
rect 14660 19892 14666 19956
rect 15510 19892 15516 19956
rect 15580 19954 15586 19956
rect 15745 19954 15811 19957
rect 15580 19952 15811 19954
rect 15580 19896 15750 19952
rect 15806 19896 15811 19952
rect 15580 19894 15811 19896
rect 15580 19892 15586 19894
rect 15745 19891 15811 19894
rect 4429 19818 4495 19821
rect 8845 19818 8911 19821
rect 4429 19816 8911 19818
rect 4429 19760 4434 19816
rect 4490 19760 8850 19816
rect 8906 19760 8911 19816
rect 4429 19758 8911 19760
rect 4429 19755 4495 19758
rect 8845 19755 8911 19758
rect 12065 19818 12131 19821
rect 12065 19816 12266 19818
rect 12065 19760 12070 19816
rect 12126 19760 12266 19816
rect 12065 19758 12266 19760
rect 12065 19755 12131 19758
rect 790 19620 796 19684
rect 860 19682 866 19684
rect 5625 19682 5691 19685
rect 860 19680 5691 19682
rect 860 19624 5630 19680
rect 5686 19624 5691 19680
rect 860 19622 5691 19624
rect 860 19620 866 19622
rect 5625 19619 5691 19622
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 2405 19546 2471 19549
rect 4981 19546 5047 19549
rect 2405 19544 5047 19546
rect 2405 19488 2410 19544
rect 2466 19488 4986 19544
rect 5042 19488 5047 19544
rect 2405 19486 5047 19488
rect 2405 19483 2471 19486
rect 4981 19483 5047 19486
rect 5257 19546 5323 19549
rect 5390 19546 5396 19548
rect 5257 19544 5396 19546
rect 5257 19488 5262 19544
rect 5318 19488 5396 19544
rect 5257 19486 5396 19488
rect 5257 19483 5323 19486
rect 5390 19484 5396 19486
rect 5460 19484 5466 19548
rect 5533 19546 5599 19549
rect 12206 19548 12266 19758
rect 14590 19756 14596 19820
rect 14660 19818 14666 19820
rect 15101 19818 15167 19821
rect 14660 19816 15167 19818
rect 14660 19760 15106 19816
rect 15162 19760 15167 19816
rect 14660 19758 15167 19760
rect 14660 19756 14666 19758
rect 15101 19755 15167 19758
rect 16205 19818 16271 19821
rect 23105 19818 23171 19821
rect 16205 19816 23171 19818
rect 16205 19760 16210 19816
rect 16266 19760 23110 19816
rect 23166 19760 23171 19816
rect 16205 19758 23171 19760
rect 16205 19755 16271 19758
rect 23105 19755 23171 19758
rect 17953 19684 18019 19685
rect 17902 19620 17908 19684
rect 17972 19682 18019 19684
rect 19241 19682 19307 19685
rect 17972 19680 19307 19682
rect 18014 19624 19246 19680
rect 19302 19624 19307 19680
rect 17972 19622 19307 19624
rect 17972 19620 18019 19622
rect 17953 19619 18019 19620
rect 19241 19619 19307 19622
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 6494 19546 6500 19548
rect 5533 19544 6500 19546
rect 5533 19488 5538 19544
rect 5594 19488 6500 19544
rect 5533 19486 6500 19488
rect 5533 19483 5599 19486
rect 6494 19484 6500 19486
rect 6564 19484 6570 19548
rect 12198 19484 12204 19548
rect 12268 19546 12274 19548
rect 14641 19546 14707 19549
rect 18229 19546 18295 19549
rect 12268 19544 14707 19546
rect 12268 19488 14646 19544
rect 14702 19488 14707 19544
rect 12268 19486 14707 19488
rect 12268 19484 12274 19486
rect 14641 19483 14707 19486
rect 16208 19544 18295 19546
rect 16208 19488 18234 19544
rect 18290 19488 18295 19544
rect 16208 19486 18295 19488
rect 16208 19413 16268 19486
rect 18229 19483 18295 19486
rect 3509 19410 3575 19413
rect 7741 19410 7807 19413
rect 3509 19408 7807 19410
rect 3509 19352 3514 19408
rect 3570 19352 7746 19408
rect 7802 19352 7807 19408
rect 3509 19350 7807 19352
rect 3509 19347 3575 19350
rect 7741 19347 7807 19350
rect 11053 19410 11119 19413
rect 11605 19410 11671 19413
rect 11053 19408 11671 19410
rect 11053 19352 11058 19408
rect 11114 19352 11610 19408
rect 11666 19352 11671 19408
rect 11053 19350 11671 19352
rect 11053 19347 11119 19350
rect 11605 19347 11671 19350
rect 12893 19410 12959 19413
rect 13486 19410 13492 19412
rect 12893 19408 13492 19410
rect 12893 19352 12898 19408
rect 12954 19352 13492 19408
rect 12893 19350 13492 19352
rect 12893 19347 12959 19350
rect 13486 19348 13492 19350
rect 13556 19348 13562 19412
rect 14406 19348 14412 19412
rect 14476 19410 14482 19412
rect 14917 19410 14983 19413
rect 14476 19408 14983 19410
rect 14476 19352 14922 19408
rect 14978 19352 14983 19408
rect 14476 19350 14983 19352
rect 14476 19348 14482 19350
rect 14917 19347 14983 19350
rect 16205 19408 16271 19413
rect 16665 19412 16731 19413
rect 16614 19410 16620 19412
rect 16205 19352 16210 19408
rect 16266 19352 16271 19408
rect 16205 19347 16271 19352
rect 16574 19350 16620 19410
rect 16684 19408 16731 19412
rect 16726 19352 16731 19408
rect 16614 19348 16620 19350
rect 16684 19348 16731 19352
rect 16665 19347 16731 19348
rect 21357 19410 21423 19413
rect 24669 19410 24735 19413
rect 21357 19408 24735 19410
rect 21357 19352 21362 19408
rect 21418 19352 24674 19408
rect 24730 19352 24735 19408
rect 21357 19350 24735 19352
rect 21357 19347 21423 19350
rect 24669 19347 24735 19350
rect 4705 19274 4771 19277
rect 7189 19274 7255 19277
rect 4705 19272 7255 19274
rect 4705 19216 4710 19272
rect 4766 19216 7194 19272
rect 7250 19216 7255 19272
rect 4705 19214 7255 19216
rect 4705 19211 4771 19214
rect 7189 19211 7255 19214
rect 8293 19274 8359 19277
rect 10777 19274 10843 19277
rect 8293 19272 10843 19274
rect 8293 19216 8298 19272
rect 8354 19216 10782 19272
rect 10838 19216 10843 19272
rect 8293 19214 10843 19216
rect 8293 19211 8359 19214
rect 10777 19211 10843 19214
rect 13261 19276 13327 19277
rect 13261 19272 13308 19276
rect 13372 19274 13378 19276
rect 15837 19274 15903 19277
rect 20437 19274 20503 19277
rect 13261 19216 13266 19272
rect 13261 19212 13308 19216
rect 13372 19214 13418 19274
rect 15837 19272 20503 19274
rect 15837 19216 15842 19272
rect 15898 19216 20442 19272
rect 20498 19216 20503 19272
rect 15837 19214 20503 19216
rect 13372 19212 13378 19214
rect 13261 19211 13327 19212
rect 15837 19211 15903 19214
rect 20437 19211 20503 19214
rect 9765 19138 9831 19141
rect 11053 19138 11119 19141
rect 9765 19136 11119 19138
rect 9765 19080 9770 19136
rect 9826 19080 11058 19136
rect 11114 19080 11119 19136
rect 9765 19078 11119 19080
rect 9765 19075 9831 19078
rect 11053 19075 11119 19078
rect 14181 19138 14247 19141
rect 19425 19140 19491 19141
rect 20161 19140 20227 19141
rect 17902 19138 17908 19140
rect 14181 19136 17908 19138
rect 14181 19080 14186 19136
rect 14242 19080 17908 19136
rect 14181 19078 17908 19080
rect 14181 19075 14247 19078
rect 17902 19076 17908 19078
rect 17972 19076 17978 19140
rect 19374 19076 19380 19140
rect 19444 19138 19491 19140
rect 19444 19136 19536 19138
rect 19486 19080 19536 19136
rect 19444 19078 19536 19080
rect 19444 19076 19491 19078
rect 20110 19076 20116 19140
rect 20180 19138 20227 19140
rect 20180 19136 20272 19138
rect 20222 19080 20272 19136
rect 20180 19078 20272 19080
rect 20180 19076 20227 19078
rect 19425 19075 19491 19076
rect 20161 19075 20227 19076
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 15653 19002 15719 19005
rect 15653 19000 15762 19002
rect 15653 18944 15658 19000
rect 15714 18944 15762 19000
rect 15653 18939 15762 18944
rect 16062 18940 16068 19004
rect 16132 19002 16138 19004
rect 16205 19002 16271 19005
rect 16132 19000 16271 19002
rect 16132 18944 16210 19000
rect 16266 18944 16271 19000
rect 16132 18942 16271 18944
rect 16132 18940 16138 18942
rect 16205 18939 16271 18942
rect 19333 19002 19399 19005
rect 19609 19002 19675 19005
rect 19333 19000 19675 19002
rect 19333 18944 19338 19000
rect 19394 18944 19614 19000
rect 19670 18944 19675 19000
rect 19333 18942 19675 18944
rect 19333 18939 19399 18942
rect 19609 18939 19675 18942
rect 8753 18866 8819 18869
rect 9029 18866 9095 18869
rect 11513 18866 11579 18869
rect 8753 18864 11579 18866
rect 8753 18808 8758 18864
rect 8814 18808 9034 18864
rect 9090 18808 11518 18864
rect 11574 18808 11579 18864
rect 8753 18806 11579 18808
rect 15702 18866 15762 18939
rect 16389 18866 16455 18869
rect 22318 18866 22324 18868
rect 15702 18864 22324 18866
rect 15702 18808 16394 18864
rect 16450 18808 22324 18864
rect 15702 18806 22324 18808
rect 8753 18803 8819 18806
rect 9029 18803 9095 18806
rect 11513 18803 11579 18806
rect 16389 18803 16455 18806
rect 22318 18804 22324 18806
rect 22388 18804 22394 18868
rect 3785 18730 3851 18733
rect 5165 18730 5231 18733
rect 3785 18728 5231 18730
rect 3785 18672 3790 18728
rect 3846 18672 5170 18728
rect 5226 18672 5231 18728
rect 3785 18670 5231 18672
rect 3785 18667 3851 18670
rect 5165 18667 5231 18670
rect 13905 18730 13971 18733
rect 15878 18730 15884 18732
rect 13905 18728 15884 18730
rect 13905 18672 13910 18728
rect 13966 18672 15884 18728
rect 13905 18670 15884 18672
rect 13905 18667 13971 18670
rect 15878 18668 15884 18670
rect 15948 18730 15954 18732
rect 17033 18730 17099 18733
rect 15948 18728 17099 18730
rect 15948 18672 17038 18728
rect 17094 18672 17099 18728
rect 15948 18670 17099 18672
rect 15948 18668 15954 18670
rect 17033 18667 17099 18670
rect 17493 18730 17559 18733
rect 20294 18730 20300 18732
rect 17493 18728 20300 18730
rect 17493 18672 17498 18728
rect 17554 18672 20300 18728
rect 17493 18670 20300 18672
rect 17493 18667 17559 18670
rect 20294 18668 20300 18670
rect 20364 18668 20370 18732
rect 2957 18594 3023 18597
rect 5533 18594 5599 18597
rect 2957 18592 5599 18594
rect 2957 18536 2962 18592
rect 3018 18536 5538 18592
rect 5594 18536 5599 18592
rect 2957 18534 5599 18536
rect 2957 18531 3023 18534
rect 5533 18531 5599 18534
rect 9765 18594 9831 18597
rect 11145 18594 11211 18597
rect 11605 18594 11671 18597
rect 9765 18592 11671 18594
rect 9765 18536 9770 18592
rect 9826 18536 11150 18592
rect 11206 18536 11610 18592
rect 11666 18536 11671 18592
rect 9765 18534 11671 18536
rect 9765 18531 9831 18534
rect 11145 18531 11211 18534
rect 11605 18531 11671 18534
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 2129 18458 2195 18461
rect 11053 18458 11119 18461
rect 12433 18458 12499 18461
rect 2129 18456 2790 18458
rect 2129 18400 2134 18456
rect 2190 18400 2790 18456
rect 2129 18398 2790 18400
rect 2129 18395 2195 18398
rect 2730 18322 2790 18398
rect 11053 18456 12499 18458
rect 11053 18400 11058 18456
rect 11114 18400 12438 18456
rect 12494 18400 12499 18456
rect 11053 18398 12499 18400
rect 11053 18395 11119 18398
rect 12433 18395 12499 18398
rect 15653 18458 15719 18461
rect 18321 18458 18387 18461
rect 15653 18456 18387 18458
rect 15653 18400 15658 18456
rect 15714 18400 18326 18456
rect 18382 18400 18387 18456
rect 15653 18398 18387 18400
rect 15653 18395 15719 18398
rect 18321 18395 18387 18398
rect 19793 18458 19859 18461
rect 20345 18458 20411 18461
rect 19793 18456 20411 18458
rect 19793 18400 19798 18456
rect 19854 18400 20350 18456
rect 20406 18400 20411 18456
rect 19793 18398 20411 18400
rect 19793 18395 19859 18398
rect 20345 18395 20411 18398
rect 4286 18322 4292 18324
rect 2730 18262 4292 18322
rect 4286 18260 4292 18262
rect 4356 18322 4362 18324
rect 9029 18322 9095 18325
rect 4356 18320 9095 18322
rect 4356 18264 9034 18320
rect 9090 18264 9095 18320
rect 4356 18262 9095 18264
rect 4356 18260 4362 18262
rect 9029 18259 9095 18262
rect 11973 18322 12039 18325
rect 12801 18322 12867 18325
rect 11973 18320 12867 18322
rect 11973 18264 11978 18320
rect 12034 18264 12806 18320
rect 12862 18264 12867 18320
rect 11973 18262 12867 18264
rect 11973 18259 12039 18262
rect 12801 18259 12867 18262
rect 14641 18322 14707 18325
rect 17033 18322 17099 18325
rect 14641 18320 17099 18322
rect 14641 18264 14646 18320
rect 14702 18264 17038 18320
rect 17094 18264 17099 18320
rect 14641 18262 17099 18264
rect 14641 18259 14707 18262
rect 17033 18259 17099 18262
rect 4521 18186 4587 18189
rect 6453 18186 6519 18189
rect 4521 18184 6519 18186
rect 4521 18128 4526 18184
rect 4582 18128 6458 18184
rect 6514 18128 6519 18184
rect 4521 18126 6519 18128
rect 4521 18123 4587 18126
rect 6453 18123 6519 18126
rect 7598 18124 7604 18188
rect 7668 18186 7674 18188
rect 7741 18186 7807 18189
rect 7668 18184 7807 18186
rect 7668 18128 7746 18184
rect 7802 18128 7807 18184
rect 7668 18126 7807 18128
rect 7668 18124 7674 18126
rect 7741 18123 7807 18126
rect 11605 18186 11671 18189
rect 11973 18186 12039 18189
rect 11605 18184 12039 18186
rect 11605 18128 11610 18184
rect 11666 18128 11978 18184
rect 12034 18128 12039 18184
rect 11605 18126 12039 18128
rect 11605 18123 11671 18126
rect 11973 18123 12039 18126
rect 15009 18186 15075 18189
rect 16389 18186 16455 18189
rect 15009 18184 16455 18186
rect 15009 18128 15014 18184
rect 15070 18128 16394 18184
rect 16450 18128 16455 18184
rect 15009 18126 16455 18128
rect 15009 18123 15075 18126
rect 16389 18123 16455 18126
rect 0 18050 400 18080
rect 565 18050 631 18053
rect 0 18048 631 18050
rect 0 17992 570 18048
rect 626 17992 631 18048
rect 0 17990 631 17992
rect 0 17960 400 17990
rect 565 17987 631 17990
rect 1894 17988 1900 18052
rect 1964 18050 1970 18052
rect 3325 18050 3391 18053
rect 1964 18048 3391 18050
rect 1964 17992 3330 18048
rect 3386 17992 3391 18048
rect 1964 17990 3391 17992
rect 1964 17988 1970 17990
rect 3325 17987 3391 17990
rect 6821 18050 6887 18053
rect 9121 18050 9187 18053
rect 11881 18052 11947 18053
rect 11830 18050 11836 18052
rect 6821 18048 9187 18050
rect 6821 17992 6826 18048
rect 6882 17992 9126 18048
rect 9182 17992 9187 18048
rect 6821 17990 9187 17992
rect 11790 17990 11836 18050
rect 11900 18048 11947 18052
rect 11942 17992 11947 18048
rect 6821 17987 6887 17990
rect 9121 17987 9187 17990
rect 11830 17988 11836 17990
rect 11900 17988 11947 17992
rect 11881 17987 11947 17988
rect 13997 18050 14063 18053
rect 14406 18050 14412 18052
rect 13997 18048 14412 18050
rect 13997 17992 14002 18048
rect 14058 17992 14412 18048
rect 13997 17990 14412 17992
rect 13997 17987 14063 17990
rect 14406 17988 14412 17990
rect 14476 17988 14482 18052
rect 15285 18050 15351 18053
rect 15653 18050 15719 18053
rect 15285 18048 15719 18050
rect 15285 17992 15290 18048
rect 15346 17992 15658 18048
rect 15714 17992 15719 18048
rect 15285 17990 15719 17992
rect 15285 17987 15351 17990
rect 15653 17987 15719 17990
rect 16021 18050 16087 18053
rect 16021 18048 16682 18050
rect 16021 17992 16026 18048
rect 16082 17992 16682 18048
rect 16021 17990 16682 17992
rect 16021 17987 16087 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 4981 17916 5047 17917
rect 4981 17914 5028 17916
rect 4936 17912 5028 17914
rect 4936 17856 4986 17912
rect 4936 17854 5028 17856
rect 4981 17852 5028 17854
rect 5092 17852 5098 17916
rect 5206 17852 5212 17916
rect 5276 17914 5282 17916
rect 6085 17914 6151 17917
rect 5276 17912 6151 17914
rect 5276 17856 6090 17912
rect 6146 17856 6151 17912
rect 5276 17854 6151 17856
rect 5276 17852 5282 17854
rect 4981 17851 5047 17852
rect 6085 17851 6151 17854
rect 13118 17852 13124 17916
rect 13188 17914 13194 17916
rect 13813 17914 13879 17917
rect 13188 17912 13879 17914
rect 13188 17856 13818 17912
rect 13874 17856 13879 17912
rect 13188 17854 13879 17856
rect 13188 17852 13194 17854
rect 13813 17851 13879 17854
rect 13997 17916 14063 17917
rect 13997 17912 14044 17916
rect 14108 17914 14114 17916
rect 15469 17914 15535 17917
rect 16389 17916 16455 17917
rect 16246 17914 16252 17916
rect 13997 17856 14002 17912
rect 13997 17852 14044 17856
rect 14108 17854 14154 17914
rect 15469 17912 16252 17914
rect 15469 17856 15474 17912
rect 15530 17856 16252 17912
rect 15469 17854 16252 17856
rect 14108 17852 14114 17854
rect 13997 17851 14063 17852
rect 15469 17851 15535 17854
rect 16246 17852 16252 17854
rect 16316 17852 16322 17916
rect 16389 17912 16436 17916
rect 16500 17914 16506 17916
rect 16622 17914 16682 17990
rect 19742 17988 19748 18052
rect 19812 18050 19818 18052
rect 19885 18050 19951 18053
rect 19812 18048 19951 18050
rect 19812 17992 19890 18048
rect 19946 17992 19951 18048
rect 19812 17990 19951 17992
rect 19812 17988 19818 17990
rect 19885 17987 19951 17990
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 17125 17914 17191 17917
rect 16389 17856 16394 17912
rect 16389 17852 16436 17856
rect 16500 17854 16546 17914
rect 16622 17912 17191 17914
rect 16622 17856 17130 17912
rect 17186 17856 17191 17912
rect 16622 17854 17191 17856
rect 16500 17852 16506 17854
rect 16389 17851 16455 17852
rect 17125 17851 17191 17854
rect 4337 17778 4403 17781
rect 7557 17778 7623 17781
rect 4337 17776 7623 17778
rect 4337 17720 4342 17776
rect 4398 17720 7562 17776
rect 7618 17720 7623 17776
rect 4337 17718 7623 17720
rect 4337 17715 4403 17718
rect 7557 17715 7623 17718
rect 9857 17778 9923 17781
rect 9990 17778 9996 17780
rect 9857 17776 9996 17778
rect 9857 17720 9862 17776
rect 9918 17720 9996 17776
rect 9857 17718 9996 17720
rect 9857 17715 9923 17718
rect 9990 17716 9996 17718
rect 10060 17716 10066 17780
rect 10317 17778 10383 17781
rect 15472 17778 15532 17851
rect 10317 17776 15532 17778
rect 10317 17720 10322 17776
rect 10378 17720 15532 17776
rect 10317 17718 15532 17720
rect 15653 17778 15719 17781
rect 16113 17778 16179 17781
rect 18086 17778 18092 17780
rect 15653 17776 18092 17778
rect 15653 17720 15658 17776
rect 15714 17720 16118 17776
rect 16174 17720 18092 17776
rect 15653 17718 18092 17720
rect 10317 17715 10383 17718
rect 15653 17715 15719 17718
rect 16113 17715 16179 17718
rect 18086 17716 18092 17718
rect 18156 17716 18162 17780
rect 18321 17778 18387 17781
rect 20529 17778 20595 17781
rect 27797 17778 27863 17781
rect 18321 17776 20595 17778
rect 18321 17720 18326 17776
rect 18382 17720 20534 17776
rect 20590 17720 20595 17776
rect 18321 17718 20595 17720
rect 18321 17715 18387 17718
rect 20529 17715 20595 17718
rect 20670 17776 27863 17778
rect 20670 17720 27802 17776
rect 27858 17720 27863 17776
rect 20670 17718 27863 17720
rect 3785 17642 3851 17645
rect 9397 17642 9463 17645
rect 3785 17640 9463 17642
rect 3785 17584 3790 17640
rect 3846 17584 9402 17640
rect 9458 17584 9463 17640
rect 3785 17582 9463 17584
rect 3785 17579 3851 17582
rect 9397 17579 9463 17582
rect 13261 17642 13327 17645
rect 17309 17642 17375 17645
rect 13261 17640 17375 17642
rect 13261 17584 13266 17640
rect 13322 17584 17314 17640
rect 17370 17584 17375 17640
rect 13261 17582 17375 17584
rect 13261 17579 13327 17582
rect 17309 17579 17375 17582
rect 12198 17444 12204 17508
rect 12268 17506 12274 17508
rect 13905 17506 13971 17509
rect 19609 17508 19675 17509
rect 12268 17504 13971 17506
rect 12268 17448 13910 17504
rect 13966 17448 13971 17504
rect 12268 17446 13971 17448
rect 12268 17444 12274 17446
rect 13905 17443 13971 17446
rect 19558 17444 19564 17508
rect 19628 17506 19675 17508
rect 20670 17506 20730 17718
rect 27797 17715 27863 17718
rect 19628 17504 20730 17506
rect 19670 17448 20730 17504
rect 19628 17446 20730 17448
rect 19628 17444 19675 17446
rect 19609 17443 19675 17444
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 16297 17370 16363 17373
rect 17493 17370 17559 17373
rect 16297 17368 17559 17370
rect 16297 17312 16302 17368
rect 16358 17312 17498 17368
rect 17554 17312 17559 17368
rect 16297 17310 17559 17312
rect 16297 17307 16363 17310
rect 17493 17307 17559 17310
rect 2262 17172 2268 17236
rect 2332 17234 2338 17236
rect 10225 17234 10291 17237
rect 2332 17232 10291 17234
rect 2332 17176 10230 17232
rect 10286 17176 10291 17232
rect 2332 17174 10291 17176
rect 2332 17172 2338 17174
rect 10225 17171 10291 17174
rect 11421 17234 11487 17237
rect 13118 17234 13124 17236
rect 11421 17232 13124 17234
rect 11421 17176 11426 17232
rect 11482 17176 13124 17232
rect 11421 17174 13124 17176
rect 11421 17171 11487 17174
rect 13118 17172 13124 17174
rect 13188 17234 13194 17236
rect 17125 17234 17191 17237
rect 13188 17232 17191 17234
rect 13188 17176 17130 17232
rect 17186 17176 17191 17232
rect 13188 17174 17191 17176
rect 13188 17172 13194 17174
rect 17125 17171 17191 17174
rect 5809 17098 5875 17101
rect 8109 17098 8175 17101
rect 5809 17096 8175 17098
rect 5809 17040 5814 17096
rect 5870 17040 8114 17096
rect 8170 17040 8175 17096
rect 5809 17038 8175 17040
rect 5809 17035 5875 17038
rect 8109 17035 8175 17038
rect 11973 17098 12039 17101
rect 16389 17098 16455 17101
rect 11973 17096 16455 17098
rect 11973 17040 11978 17096
rect 12034 17040 16394 17096
rect 16450 17040 16455 17096
rect 11973 17038 16455 17040
rect 11973 17035 12039 17038
rect 16389 17035 16455 17038
rect 16941 17098 17007 17101
rect 17309 17098 17375 17101
rect 19977 17098 20043 17101
rect 20897 17098 20963 17101
rect 16941 17096 20963 17098
rect 16941 17040 16946 17096
rect 17002 17040 17314 17096
rect 17370 17040 19982 17096
rect 20038 17040 20902 17096
rect 20958 17040 20963 17096
rect 16941 17038 20963 17040
rect 16941 17035 17007 17038
rect 17309 17035 17375 17038
rect 19977 17035 20043 17038
rect 20897 17035 20963 17038
rect 13261 16962 13327 16965
rect 16021 16962 16087 16965
rect 13261 16960 16087 16962
rect 13261 16904 13266 16960
rect 13322 16904 16026 16960
rect 16082 16904 16087 16960
rect 13261 16902 16087 16904
rect 13261 16899 13327 16902
rect 16021 16899 16087 16902
rect 19374 16900 19380 16964
rect 19444 16962 19450 16964
rect 24577 16962 24643 16965
rect 19444 16960 24643 16962
rect 19444 16904 24582 16960
rect 24638 16904 24643 16960
rect 19444 16902 24643 16904
rect 19444 16900 19450 16902
rect 24577 16899 24643 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 3693 16692 3759 16693
rect 3693 16688 3740 16692
rect 3804 16690 3810 16692
rect 4153 16690 4219 16693
rect 4286 16690 4292 16692
rect 3693 16632 3698 16688
rect 3693 16628 3740 16632
rect 3804 16630 3850 16690
rect 4153 16688 4292 16690
rect 4153 16632 4158 16688
rect 4214 16632 4292 16688
rect 4153 16630 4292 16632
rect 3804 16628 3810 16630
rect 3693 16627 3759 16628
rect 4153 16627 4219 16630
rect 4286 16628 4292 16630
rect 4356 16628 4362 16692
rect 17125 16690 17191 16693
rect 18597 16690 18663 16693
rect 17125 16688 18663 16690
rect 17125 16632 17130 16688
rect 17186 16632 18602 16688
rect 18658 16632 18663 16688
rect 17125 16630 18663 16632
rect 17125 16627 17191 16630
rect 18597 16627 18663 16630
rect 6678 16492 6684 16556
rect 6748 16554 6754 16556
rect 7741 16554 7807 16557
rect 6748 16552 7807 16554
rect 6748 16496 7746 16552
rect 7802 16496 7807 16552
rect 6748 16494 7807 16496
rect 6748 16492 6754 16494
rect 7741 16491 7807 16494
rect 10225 16554 10291 16557
rect 11421 16554 11487 16557
rect 10225 16552 11487 16554
rect 10225 16496 10230 16552
rect 10286 16496 11426 16552
rect 11482 16496 11487 16552
rect 10225 16494 11487 16496
rect 10225 16491 10291 16494
rect 11421 16491 11487 16494
rect 16389 16554 16455 16557
rect 20989 16554 21055 16557
rect 16389 16552 21055 16554
rect 16389 16496 16394 16552
rect 16450 16496 20994 16552
rect 21050 16496 21055 16552
rect 16389 16494 21055 16496
rect 16389 16491 16455 16494
rect 20989 16491 21055 16494
rect 9857 16418 9923 16421
rect 10041 16418 10107 16421
rect 10777 16418 10843 16421
rect 11513 16418 11579 16421
rect 9857 16416 11579 16418
rect 9857 16360 9862 16416
rect 9918 16360 10046 16416
rect 10102 16360 10782 16416
rect 10838 16360 11518 16416
rect 11574 16360 11579 16416
rect 9857 16358 11579 16360
rect 9857 16355 9923 16358
rect 10041 16355 10107 16358
rect 10777 16355 10843 16358
rect 11513 16355 11579 16358
rect 18689 16418 18755 16421
rect 18822 16418 18828 16420
rect 18689 16416 18828 16418
rect 18689 16360 18694 16416
rect 18750 16360 18828 16416
rect 18689 16358 18828 16360
rect 18689 16355 18755 16358
rect 18822 16356 18828 16358
rect 18892 16356 18898 16420
rect 19241 16418 19307 16421
rect 21541 16418 21607 16421
rect 19241 16416 21607 16418
rect 19241 16360 19246 16416
rect 19302 16360 21546 16416
rect 21602 16360 21607 16416
rect 19241 16358 21607 16360
rect 19241 16355 19307 16358
rect 21541 16355 21607 16358
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 1393 16282 1459 16285
rect 7414 16282 7420 16284
rect 1393 16280 7420 16282
rect 1393 16224 1398 16280
rect 1454 16224 7420 16280
rect 1393 16222 7420 16224
rect 1393 16219 1459 16222
rect 7414 16220 7420 16222
rect 7484 16282 7490 16284
rect 7557 16282 7623 16285
rect 7484 16280 7623 16282
rect 7484 16224 7562 16280
rect 7618 16224 7623 16280
rect 7484 16222 7623 16224
rect 7484 16220 7490 16222
rect 7557 16219 7623 16222
rect 19885 16282 19951 16285
rect 21081 16282 21147 16285
rect 19885 16280 21147 16282
rect 19885 16224 19890 16280
rect 19946 16224 21086 16280
rect 21142 16224 21147 16280
rect 19885 16222 21147 16224
rect 19885 16219 19951 16222
rect 21081 16219 21147 16222
rect 6453 16148 6519 16149
rect 6453 16146 6500 16148
rect 6408 16144 6500 16146
rect 6408 16088 6458 16144
rect 6408 16086 6500 16088
rect 6453 16084 6500 16086
rect 6564 16084 6570 16148
rect 7005 16146 7071 16149
rect 9806 16146 9812 16148
rect 7005 16144 9812 16146
rect 7005 16088 7010 16144
rect 7066 16088 9812 16144
rect 7005 16086 9812 16088
rect 6453 16083 6519 16084
rect 7005 16083 7071 16086
rect 9806 16084 9812 16086
rect 9876 16084 9882 16148
rect 10041 16146 10107 16149
rect 11237 16146 11303 16149
rect 10041 16144 11303 16146
rect 10041 16088 10046 16144
rect 10102 16088 11242 16144
rect 11298 16088 11303 16144
rect 10041 16086 11303 16088
rect 10041 16083 10107 16086
rect 11237 16083 11303 16086
rect 11830 16084 11836 16148
rect 11900 16146 11906 16148
rect 15377 16146 15443 16149
rect 11900 16144 15443 16146
rect 11900 16088 15382 16144
rect 15438 16088 15443 16144
rect 11900 16086 15443 16088
rect 11900 16084 11906 16086
rect 15377 16083 15443 16086
rect 19333 16148 19399 16149
rect 19333 16144 19380 16148
rect 19444 16146 19450 16148
rect 19333 16088 19338 16144
rect 19333 16084 19380 16088
rect 19444 16086 19490 16146
rect 19444 16084 19450 16086
rect 19333 16083 19399 16084
rect 0 16010 400 16040
rect 473 16010 539 16013
rect 13537 16012 13603 16013
rect 0 16008 539 16010
rect 0 15952 478 16008
rect 534 15952 539 16008
rect 0 15950 539 15952
rect 0 15920 400 15950
rect 473 15947 539 15950
rect 13486 15948 13492 16012
rect 13556 16010 13603 16012
rect 13556 16008 13648 16010
rect 13598 15952 13648 16008
rect 13556 15950 13648 15952
rect 13556 15948 13603 15950
rect 13537 15947 13603 15948
rect 15326 15812 15332 15876
rect 15396 15874 15402 15876
rect 17769 15874 17835 15877
rect 15396 15872 17835 15874
rect 15396 15816 17774 15872
rect 17830 15816 17835 15872
rect 15396 15814 17835 15816
rect 15396 15812 15402 15814
rect 17769 15811 17835 15814
rect 21357 15874 21423 15877
rect 21541 15874 21607 15877
rect 21357 15872 21607 15874
rect 21357 15816 21362 15872
rect 21418 15816 21546 15872
rect 21602 15816 21607 15872
rect 21357 15814 21607 15816
rect 21357 15811 21423 15814
rect 21541 15811 21607 15814
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 2681 15602 2747 15605
rect 7557 15602 7623 15605
rect 2681 15600 7623 15602
rect 2681 15544 2686 15600
rect 2742 15544 7562 15600
rect 7618 15544 7623 15600
rect 2681 15542 7623 15544
rect 2681 15539 2747 15542
rect 7557 15539 7623 15542
rect 11881 15602 11947 15605
rect 13077 15602 13143 15605
rect 11881 15600 13143 15602
rect 11881 15544 11886 15600
rect 11942 15544 13082 15600
rect 13138 15544 13143 15600
rect 11881 15542 13143 15544
rect 11881 15539 11947 15542
rect 13077 15539 13143 15542
rect 3785 15466 3851 15469
rect 7046 15466 7052 15468
rect 3785 15464 7052 15466
rect 3785 15408 3790 15464
rect 3846 15408 7052 15464
rect 3785 15406 7052 15408
rect 3785 15403 3851 15406
rect 7046 15404 7052 15406
rect 7116 15466 7122 15468
rect 8845 15466 8911 15469
rect 7116 15464 8911 15466
rect 7116 15408 8850 15464
rect 8906 15408 8911 15464
rect 7116 15406 8911 15408
rect 7116 15404 7122 15406
rect 8845 15403 8911 15406
rect 13905 15466 13971 15469
rect 16614 15466 16620 15468
rect 13905 15464 16620 15466
rect 13905 15408 13910 15464
rect 13966 15408 16620 15464
rect 13905 15406 16620 15408
rect 13905 15403 13971 15406
rect 16614 15404 16620 15406
rect 16684 15404 16690 15468
rect 2630 15268 2636 15332
rect 2700 15330 2706 15332
rect 6637 15330 6703 15333
rect 2700 15328 6703 15330
rect 2700 15272 6642 15328
rect 6698 15272 6703 15328
rect 2700 15270 6703 15272
rect 2700 15268 2706 15270
rect 6637 15267 6703 15270
rect 9581 15330 9647 15333
rect 13670 15330 13676 15332
rect 9581 15328 13676 15330
rect 9581 15272 9586 15328
rect 9642 15272 13676 15328
rect 9581 15270 13676 15272
rect 9581 15267 9647 15270
rect 13670 15268 13676 15270
rect 13740 15268 13746 15332
rect 16297 15330 16363 15333
rect 18965 15330 19031 15333
rect 16297 15328 19031 15330
rect 16297 15272 16302 15328
rect 16358 15272 18970 15328
rect 19026 15272 19031 15328
rect 16297 15270 19031 15272
rect 16297 15267 16363 15270
rect 18965 15267 19031 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 7230 15132 7236 15196
rect 7300 15194 7306 15196
rect 7465 15194 7531 15197
rect 7300 15192 7531 15194
rect 7300 15136 7470 15192
rect 7526 15136 7531 15192
rect 7300 15134 7531 15136
rect 7300 15132 7306 15134
rect 7465 15131 7531 15134
rect 11145 15194 11211 15197
rect 13997 15194 14063 15197
rect 11145 15192 14063 15194
rect 11145 15136 11150 15192
rect 11206 15136 14002 15192
rect 14058 15136 14063 15192
rect 11145 15134 14063 15136
rect 11145 15131 11211 15134
rect 13997 15131 14063 15134
rect 17861 15194 17927 15197
rect 20478 15194 20484 15196
rect 17861 15192 20484 15194
rect 17861 15136 17866 15192
rect 17922 15136 20484 15192
rect 17861 15134 20484 15136
rect 17861 15131 17927 15134
rect 20478 15132 20484 15134
rect 20548 15132 20554 15196
rect 16021 15058 16087 15061
rect 23105 15058 23171 15061
rect 16021 15056 23171 15058
rect 16021 15000 16026 15056
rect 16082 15000 23110 15056
rect 23166 15000 23171 15056
rect 16021 14998 23171 15000
rect 16021 14995 16087 14998
rect 23105 14995 23171 14998
rect 12433 14922 12499 14925
rect 16062 14922 16068 14924
rect 12433 14920 16068 14922
rect 12433 14864 12438 14920
rect 12494 14864 16068 14920
rect 12433 14862 16068 14864
rect 12433 14859 12499 14862
rect 16062 14860 16068 14862
rect 16132 14922 16138 14924
rect 17677 14922 17743 14925
rect 16132 14920 17743 14922
rect 16132 14864 17682 14920
rect 17738 14864 17743 14920
rect 16132 14862 17743 14864
rect 16132 14860 16138 14862
rect 17677 14859 17743 14862
rect 20713 14922 20779 14925
rect 24301 14922 24367 14925
rect 20713 14920 24367 14922
rect 20713 14864 20718 14920
rect 20774 14864 24306 14920
rect 24362 14864 24367 14920
rect 20713 14862 24367 14864
rect 20713 14859 20779 14862
rect 24301 14859 24367 14862
rect 14406 14724 14412 14788
rect 14476 14786 14482 14788
rect 15653 14786 15719 14789
rect 14476 14784 15719 14786
rect 14476 14728 15658 14784
rect 15714 14728 15719 14784
rect 14476 14726 15719 14728
rect 14476 14724 14482 14726
rect 15653 14723 15719 14726
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 12065 14650 12131 14653
rect 14273 14650 14339 14653
rect 16941 14650 17007 14653
rect 12065 14648 17007 14650
rect 12065 14592 12070 14648
rect 12126 14592 14278 14648
rect 14334 14592 16946 14648
rect 17002 14592 17007 14648
rect 12065 14590 17007 14592
rect 12065 14587 12131 14590
rect 14273 14587 14339 14590
rect 16941 14587 17007 14590
rect 2129 14514 2195 14517
rect 13353 14514 13419 14517
rect 2129 14512 13419 14514
rect 2129 14456 2134 14512
rect 2190 14456 13358 14512
rect 13414 14456 13419 14512
rect 2129 14454 13419 14456
rect 2129 14451 2195 14454
rect 13353 14451 13419 14454
rect 15009 14514 15075 14517
rect 18137 14514 18203 14517
rect 19977 14516 20043 14517
rect 19926 14514 19932 14516
rect 15009 14512 18203 14514
rect 15009 14456 15014 14512
rect 15070 14456 18142 14512
rect 18198 14456 18203 14512
rect 15009 14454 18203 14456
rect 19886 14454 19932 14514
rect 19996 14512 20043 14516
rect 20038 14456 20043 14512
rect 15009 14451 15075 14454
rect 18137 14451 18203 14454
rect 19926 14452 19932 14454
rect 19996 14452 20043 14456
rect 19977 14451 20043 14452
rect 20345 14514 20411 14517
rect 21357 14514 21423 14517
rect 22369 14514 22435 14517
rect 20345 14512 22435 14514
rect 20345 14456 20350 14512
rect 20406 14456 21362 14512
rect 21418 14456 22374 14512
rect 22430 14456 22435 14512
rect 20345 14454 22435 14456
rect 20345 14451 20411 14454
rect 21357 14451 21423 14454
rect 22369 14451 22435 14454
rect 974 14316 980 14380
rect 1044 14378 1050 14380
rect 8201 14378 8267 14381
rect 1044 14376 8267 14378
rect 1044 14320 8206 14376
rect 8262 14320 8267 14376
rect 1044 14318 8267 14320
rect 1044 14316 1050 14318
rect 8201 14315 8267 14318
rect 10869 14378 10935 14381
rect 12249 14378 12315 14381
rect 10869 14376 12315 14378
rect 10869 14320 10874 14376
rect 10930 14320 12254 14376
rect 12310 14320 12315 14376
rect 10869 14318 12315 14320
rect 10869 14315 10935 14318
rect 12249 14315 12315 14318
rect 14641 14378 14707 14381
rect 16665 14378 16731 14381
rect 14641 14376 16731 14378
rect 14641 14320 14646 14376
rect 14702 14320 16670 14376
rect 16726 14320 16731 14376
rect 14641 14318 16731 14320
rect 14641 14315 14707 14318
rect 16665 14315 16731 14318
rect 19977 14378 20043 14381
rect 20805 14378 20871 14381
rect 19977 14376 20871 14378
rect 19977 14320 19982 14376
rect 20038 14320 20810 14376
rect 20866 14320 20871 14376
rect 19977 14318 20871 14320
rect 19977 14315 20043 14318
rect 20805 14315 20871 14318
rect 1761 14242 1827 14245
rect 4521 14242 4587 14245
rect 1761 14240 4587 14242
rect 1761 14184 1766 14240
rect 1822 14184 4526 14240
rect 4582 14184 4587 14240
rect 1761 14182 4587 14184
rect 1761 14179 1827 14182
rect 4521 14179 4587 14182
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 11329 14106 11395 14109
rect 12157 14106 12223 14109
rect 11329 14104 14612 14106
rect 11329 14048 11334 14104
rect 11390 14048 12162 14104
rect 12218 14048 14612 14104
rect 11329 14046 14612 14048
rect 11329 14043 11395 14046
rect 12157 14043 12223 14046
rect 0 13970 400 14000
rect 473 13970 539 13973
rect 0 13968 539 13970
rect 0 13912 478 13968
rect 534 13912 539 13968
rect 0 13910 539 13912
rect 0 13880 400 13910
rect 473 13907 539 13910
rect 1945 13970 2011 13973
rect 6453 13970 6519 13973
rect 1945 13968 6519 13970
rect 1945 13912 1950 13968
rect 2006 13912 6458 13968
rect 6514 13912 6519 13968
rect 1945 13910 6519 13912
rect 1945 13907 2011 13910
rect 6453 13907 6519 13910
rect 6729 13970 6795 13973
rect 7189 13970 7255 13973
rect 6729 13968 7255 13970
rect 6729 13912 6734 13968
rect 6790 13912 7194 13968
rect 7250 13912 7255 13968
rect 6729 13910 7255 13912
rect 6729 13907 6795 13910
rect 7189 13907 7255 13910
rect 7925 13970 7991 13973
rect 9213 13970 9279 13973
rect 7925 13968 9279 13970
rect 7925 13912 7930 13968
rect 7986 13912 9218 13968
rect 9274 13912 9279 13968
rect 7925 13910 9279 13912
rect 7925 13907 7991 13910
rect 9213 13907 9279 13910
rect 11094 13908 11100 13972
rect 11164 13970 11170 13972
rect 13721 13970 13787 13973
rect 11164 13968 13787 13970
rect 11164 13912 13726 13968
rect 13782 13912 13787 13968
rect 11164 13910 13787 13912
rect 11164 13908 11170 13910
rect 13721 13907 13787 13910
rect 14222 13908 14228 13972
rect 14292 13970 14298 13972
rect 14365 13970 14431 13973
rect 14292 13968 14431 13970
rect 14292 13912 14370 13968
rect 14426 13912 14431 13968
rect 14292 13910 14431 13912
rect 14552 13970 14612 14046
rect 16113 13970 16179 13973
rect 14552 13968 16179 13970
rect 14552 13912 16118 13968
rect 16174 13912 16179 13968
rect 14552 13910 16179 13912
rect 14292 13908 14298 13910
rect 14365 13907 14431 13910
rect 16113 13907 16179 13910
rect 17125 13970 17191 13973
rect 18505 13970 18571 13973
rect 17125 13968 18571 13970
rect 17125 13912 17130 13968
rect 17186 13912 18510 13968
rect 18566 13912 18571 13968
rect 17125 13910 18571 13912
rect 17125 13907 17191 13910
rect 18505 13907 18571 13910
rect 22185 13970 22251 13973
rect 25497 13970 25563 13973
rect 22185 13968 25563 13970
rect 22185 13912 22190 13968
rect 22246 13912 25502 13968
rect 25558 13912 25563 13968
rect 22185 13910 25563 13912
rect 22185 13907 22251 13910
rect 25497 13907 25563 13910
rect 5901 13834 5967 13837
rect 7557 13834 7623 13837
rect 8753 13834 8819 13837
rect 5901 13832 8819 13834
rect 5901 13776 5906 13832
rect 5962 13776 7562 13832
rect 7618 13776 8758 13832
rect 8814 13776 8819 13832
rect 5901 13774 8819 13776
rect 5901 13771 5967 13774
rect 7557 13771 7623 13774
rect 8753 13771 8819 13774
rect 9438 13772 9444 13836
rect 9508 13834 9514 13836
rect 12709 13834 12775 13837
rect 13537 13836 13603 13837
rect 13486 13834 13492 13836
rect 9508 13832 12775 13834
rect 9508 13776 12714 13832
rect 12770 13776 12775 13832
rect 9508 13774 12775 13776
rect 13446 13774 13492 13834
rect 13556 13832 13603 13836
rect 13598 13776 13603 13832
rect 9508 13772 9514 13774
rect 12709 13771 12775 13774
rect 13486 13772 13492 13774
rect 13556 13772 13603 13776
rect 13537 13771 13603 13772
rect 18321 13834 18387 13837
rect 18781 13834 18847 13837
rect 18321 13832 18847 13834
rect 18321 13776 18326 13832
rect 18382 13776 18786 13832
rect 18842 13776 18847 13832
rect 18321 13774 18847 13776
rect 18321 13771 18387 13774
rect 18781 13771 18847 13774
rect 22093 13834 22159 13837
rect 27705 13834 27771 13837
rect 22093 13832 27771 13834
rect 22093 13776 22098 13832
rect 22154 13776 27710 13832
rect 27766 13776 27771 13832
rect 22093 13774 27771 13776
rect 22093 13771 22159 13774
rect 27705 13771 27771 13774
rect 7005 13698 7071 13701
rect 9949 13698 10015 13701
rect 7005 13696 10015 13698
rect 7005 13640 7010 13696
rect 7066 13640 9954 13696
rect 10010 13640 10015 13696
rect 7005 13638 10015 13640
rect 7005 13635 7071 13638
rect 9949 13635 10015 13638
rect 11789 13698 11855 13701
rect 12014 13698 12020 13700
rect 11789 13696 12020 13698
rect 11789 13640 11794 13696
rect 11850 13640 12020 13696
rect 11789 13638 12020 13640
rect 11789 13635 11855 13638
rect 12014 13636 12020 13638
rect 12084 13698 12090 13700
rect 16297 13698 16363 13701
rect 12084 13696 16363 13698
rect 12084 13640 16302 13696
rect 16358 13640 16363 13696
rect 12084 13638 16363 13640
rect 12084 13636 12090 13638
rect 16297 13635 16363 13638
rect 17401 13698 17467 13701
rect 17769 13698 17835 13701
rect 17401 13696 17835 13698
rect 17401 13640 17406 13696
rect 17462 13640 17774 13696
rect 17830 13640 17835 13696
rect 17401 13638 17835 13640
rect 17401 13635 17467 13638
rect 17769 13635 17835 13638
rect 19885 13698 19951 13701
rect 20110 13698 20116 13700
rect 19885 13696 20116 13698
rect 19885 13640 19890 13696
rect 19946 13640 20116 13696
rect 19885 13638 20116 13640
rect 19885 13635 19951 13638
rect 20110 13636 20116 13638
rect 20180 13636 20186 13700
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 8661 13562 8727 13565
rect 9254 13562 9260 13564
rect 8661 13560 9260 13562
rect 8661 13504 8666 13560
rect 8722 13504 9260 13560
rect 8661 13502 9260 13504
rect 8661 13499 8727 13502
rect 9254 13500 9260 13502
rect 9324 13500 9330 13564
rect 9489 13562 9555 13565
rect 11053 13562 11119 13565
rect 15510 13562 15516 13564
rect 9489 13560 11119 13562
rect 9489 13504 9494 13560
rect 9550 13504 11058 13560
rect 11114 13504 11119 13560
rect 9489 13502 11119 13504
rect 9489 13499 9555 13502
rect 11053 13499 11119 13502
rect 12390 13502 15516 13562
rect 8017 13426 8083 13429
rect 5168 13424 8083 13426
rect 5168 13368 8022 13424
rect 8078 13368 8083 13424
rect 5168 13366 8083 13368
rect 5168 13293 5228 13366
rect 8017 13363 8083 13366
rect 9305 13426 9371 13429
rect 12390 13426 12450 13502
rect 15510 13500 15516 13502
rect 15580 13500 15586 13564
rect 9305 13424 12450 13426
rect 9305 13368 9310 13424
rect 9366 13368 12450 13424
rect 9305 13366 12450 13368
rect 14181 13426 14247 13429
rect 14406 13426 14412 13428
rect 14181 13424 14412 13426
rect 14181 13368 14186 13424
rect 14242 13368 14412 13424
rect 14181 13366 14412 13368
rect 9305 13363 9371 13366
rect 14181 13363 14247 13366
rect 14406 13364 14412 13366
rect 14476 13364 14482 13428
rect 14549 13426 14615 13429
rect 16849 13426 16915 13429
rect 14549 13424 16915 13426
rect 14549 13368 14554 13424
rect 14610 13368 16854 13424
rect 16910 13368 16915 13424
rect 14549 13366 16915 13368
rect 14549 13363 14615 13366
rect 16849 13363 16915 13366
rect 17033 13426 17099 13429
rect 19558 13426 19564 13428
rect 17033 13424 19564 13426
rect 17033 13368 17038 13424
rect 17094 13368 19564 13424
rect 17033 13366 19564 13368
rect 17033 13363 17099 13366
rect 19558 13364 19564 13366
rect 19628 13364 19634 13428
rect 5165 13288 5231 13293
rect 5165 13232 5170 13288
rect 5226 13232 5231 13288
rect 5165 13227 5231 13232
rect 6913 13290 6979 13293
rect 9029 13290 9095 13293
rect 6913 13288 9095 13290
rect 6913 13232 6918 13288
rect 6974 13232 9034 13288
rect 9090 13232 9095 13288
rect 6913 13230 9095 13232
rect 6913 13227 6979 13230
rect 9029 13227 9095 13230
rect 13537 13290 13603 13293
rect 19057 13290 19123 13293
rect 13537 13288 19123 13290
rect 13537 13232 13542 13288
rect 13598 13232 19062 13288
rect 19118 13232 19123 13288
rect 13537 13230 19123 13232
rect 13537 13227 13603 13230
rect 19057 13227 19123 13230
rect 10317 13154 10383 13157
rect 12433 13154 12499 13157
rect 10317 13152 12499 13154
rect 10317 13096 10322 13152
rect 10378 13096 12438 13152
rect 12494 13096 12499 13152
rect 10317 13094 12499 13096
rect 10317 13091 10383 13094
rect 12433 13091 12499 13094
rect 15653 13154 15719 13157
rect 17350 13154 17356 13156
rect 15653 13152 17356 13154
rect 15653 13096 15658 13152
rect 15714 13096 17356 13152
rect 15653 13094 17356 13096
rect 15653 13091 15719 13094
rect 17350 13092 17356 13094
rect 17420 13092 17426 13156
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 4337 12884 4403 12885
rect 4286 12820 4292 12884
rect 4356 12882 4403 12884
rect 4356 12880 4448 12882
rect 4398 12824 4448 12880
rect 4356 12822 4448 12824
rect 4356 12820 4403 12822
rect 5206 12820 5212 12884
rect 5276 12882 5282 12884
rect 5276 12822 7482 12882
rect 5276 12820 5282 12822
rect 4337 12819 4403 12820
rect 749 12746 815 12749
rect 7281 12746 7347 12749
rect 749 12744 7347 12746
rect 749 12688 754 12744
rect 810 12688 7286 12744
rect 7342 12688 7347 12744
rect 749 12686 7347 12688
rect 7422 12746 7482 12822
rect 14590 12820 14596 12884
rect 14660 12882 14666 12884
rect 15101 12882 15167 12885
rect 14660 12880 15167 12882
rect 14660 12824 15106 12880
rect 15162 12824 15167 12880
rect 14660 12822 15167 12824
rect 14660 12820 14666 12822
rect 15101 12819 15167 12822
rect 17861 12882 17927 12885
rect 18873 12882 18939 12885
rect 17861 12880 18939 12882
rect 17861 12824 17866 12880
rect 17922 12824 18878 12880
rect 18934 12824 18939 12880
rect 17861 12822 18939 12824
rect 17861 12819 17927 12822
rect 18873 12819 18939 12822
rect 7557 12748 7623 12749
rect 10225 12748 10291 12749
rect 7557 12746 7604 12748
rect 7422 12744 7604 12746
rect 7422 12688 7562 12744
rect 7422 12686 7604 12688
rect 749 12683 815 12686
rect 7281 12683 7347 12686
rect 7557 12684 7604 12686
rect 7668 12684 7674 12748
rect 10174 12746 10180 12748
rect 10134 12686 10180 12746
rect 10244 12744 10291 12748
rect 10286 12688 10291 12744
rect 10174 12684 10180 12686
rect 10244 12684 10291 12688
rect 7557 12683 7623 12684
rect 10225 12683 10291 12684
rect 11605 12746 11671 12749
rect 12893 12746 12959 12749
rect 11605 12744 12959 12746
rect 11605 12688 11610 12744
rect 11666 12688 12898 12744
rect 12954 12688 12959 12744
rect 11605 12686 12959 12688
rect 11605 12683 11671 12686
rect 12893 12683 12959 12686
rect 15561 12746 15627 12749
rect 17902 12746 17908 12748
rect 15561 12744 17908 12746
rect 15561 12688 15566 12744
rect 15622 12688 17908 12744
rect 15561 12686 17908 12688
rect 15561 12683 15627 12686
rect 17902 12684 17908 12686
rect 17972 12684 17978 12748
rect 24393 12746 24459 12749
rect 25313 12746 25379 12749
rect 24393 12744 25379 12746
rect 24393 12688 24398 12744
rect 24454 12688 25318 12744
rect 25374 12688 25379 12744
rect 24393 12686 25379 12688
rect 24393 12683 24459 12686
rect 25313 12683 25379 12686
rect 7649 12610 7715 12613
rect 6732 12608 7715 12610
rect 6732 12552 7654 12608
rect 7710 12552 7715 12608
rect 6732 12550 7715 12552
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 54 12412 60 12476
rect 124 12474 130 12476
rect 2865 12474 2931 12477
rect 124 12472 2931 12474
rect 124 12416 2870 12472
rect 2926 12416 2931 12472
rect 124 12414 2931 12416
rect 124 12412 130 12414
rect 2865 12411 2931 12414
rect 5390 12412 5396 12476
rect 5460 12474 5466 12476
rect 5901 12474 5967 12477
rect 5460 12472 5967 12474
rect 5460 12416 5906 12472
rect 5962 12416 5967 12472
rect 5460 12414 5967 12416
rect 5460 12412 5466 12414
rect 5901 12411 5967 12414
rect 6453 12474 6519 12477
rect 6732 12474 6792 12550
rect 7649 12547 7715 12550
rect 8661 12610 8727 12613
rect 9029 12610 9095 12613
rect 8661 12608 9095 12610
rect 8661 12552 8666 12608
rect 8722 12552 9034 12608
rect 9090 12552 9095 12608
rect 8661 12550 9095 12552
rect 8661 12547 8727 12550
rect 9029 12547 9095 12550
rect 19977 12610 20043 12613
rect 23289 12610 23355 12613
rect 19977 12608 23355 12610
rect 19977 12552 19982 12608
rect 20038 12552 23294 12608
rect 23350 12552 23355 12608
rect 19977 12550 23355 12552
rect 19977 12547 20043 12550
rect 23289 12547 23355 12550
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 6453 12472 6792 12474
rect 6453 12416 6458 12472
rect 6514 12416 6792 12472
rect 6453 12414 6792 12416
rect 6913 12474 6979 12477
rect 7281 12474 7347 12477
rect 6913 12472 7347 12474
rect 6913 12416 6918 12472
rect 6974 12416 7286 12472
rect 7342 12416 7347 12472
rect 6913 12414 7347 12416
rect 6453 12411 6519 12414
rect 6913 12411 6979 12414
rect 7281 12411 7347 12414
rect 8845 12474 8911 12477
rect 9397 12474 9463 12477
rect 8845 12472 9463 12474
rect 8845 12416 8850 12472
rect 8906 12416 9402 12472
rect 9458 12416 9463 12472
rect 8845 12414 9463 12416
rect 8845 12411 8911 12414
rect 9397 12411 9463 12414
rect 9949 12474 10015 12477
rect 10777 12474 10843 12477
rect 17493 12476 17559 12477
rect 17493 12474 17540 12476
rect 9949 12472 10843 12474
rect 9949 12416 9954 12472
rect 10010 12416 10782 12472
rect 10838 12416 10843 12472
rect 9949 12414 10843 12416
rect 17448 12472 17540 12474
rect 17448 12416 17498 12472
rect 17448 12414 17540 12416
rect 9949 12411 10015 12414
rect 10777 12411 10843 12414
rect 17493 12412 17540 12414
rect 17604 12412 17610 12476
rect 17493 12411 17559 12412
rect 2313 12338 2379 12341
rect 5073 12338 5139 12341
rect 2313 12336 5139 12338
rect 2313 12280 2318 12336
rect 2374 12280 5078 12336
rect 5134 12280 5139 12336
rect 2313 12278 5139 12280
rect 2313 12275 2379 12278
rect 5073 12275 5139 12278
rect 8201 12338 8267 12341
rect 12525 12338 12591 12341
rect 8201 12336 12591 12338
rect 8201 12280 8206 12336
rect 8262 12280 12530 12336
rect 12586 12280 12591 12336
rect 8201 12278 12591 12280
rect 8201 12275 8267 12278
rect 12525 12275 12591 12278
rect 15101 12338 15167 12341
rect 19793 12340 19859 12341
rect 15326 12338 15332 12340
rect 15101 12336 15332 12338
rect 15101 12280 15106 12336
rect 15162 12280 15332 12336
rect 15101 12278 15332 12280
rect 15101 12275 15167 12278
rect 15326 12276 15332 12278
rect 15396 12276 15402 12340
rect 19742 12276 19748 12340
rect 19812 12338 19859 12340
rect 19812 12336 19904 12338
rect 19854 12280 19904 12336
rect 19812 12278 19904 12280
rect 19812 12276 19859 12278
rect 19793 12275 19859 12276
rect 3918 12140 3924 12204
rect 3988 12202 3994 12204
rect 6821 12202 6887 12205
rect 3988 12200 6887 12202
rect 3988 12144 6826 12200
rect 6882 12144 6887 12200
rect 3988 12142 6887 12144
rect 3988 12140 3994 12142
rect 6821 12139 6887 12142
rect 13905 12202 13971 12205
rect 15561 12202 15627 12205
rect 13905 12200 15627 12202
rect 13905 12144 13910 12200
rect 13966 12144 15566 12200
rect 15622 12144 15627 12200
rect 13905 12142 15627 12144
rect 13905 12139 13971 12142
rect 15561 12139 15627 12142
rect 22093 12202 22159 12205
rect 22921 12202 22987 12205
rect 25129 12202 25195 12205
rect 22093 12200 25195 12202
rect 22093 12144 22098 12200
rect 22154 12144 22926 12200
rect 22982 12144 25134 12200
rect 25190 12144 25195 12200
rect 22093 12142 25195 12144
rect 22093 12139 22159 12142
rect 22921 12139 22987 12142
rect 25129 12139 25195 12142
rect 1761 12066 1827 12069
rect 2262 12066 2268 12068
rect 1761 12064 2268 12066
rect 1761 12008 1766 12064
rect 1822 12008 2268 12064
rect 1761 12006 2268 12008
rect 1761 12003 1827 12006
rect 2262 12004 2268 12006
rect 2332 12004 2338 12068
rect 6453 12066 6519 12069
rect 7189 12066 7255 12069
rect 6453 12064 7255 12066
rect 6453 12008 6458 12064
rect 6514 12008 7194 12064
rect 7250 12008 7255 12064
rect 6453 12006 7255 12008
rect 6453 12003 6519 12006
rect 7189 12003 7255 12006
rect 9765 12066 9831 12069
rect 10358 12066 10364 12068
rect 9765 12064 10364 12066
rect 9765 12008 9770 12064
rect 9826 12008 10364 12064
rect 9765 12006 10364 12008
rect 9765 12003 9831 12006
rect 10358 12004 10364 12006
rect 10428 12004 10434 12068
rect 15561 12066 15627 12069
rect 16021 12066 16087 12069
rect 15561 12064 16087 12066
rect 15561 12008 15566 12064
rect 15622 12008 16026 12064
rect 16082 12008 16087 12064
rect 15561 12006 16087 12008
rect 15561 12003 15627 12006
rect 16021 12003 16087 12006
rect 7892 12000 8208 12001
rect 0 11930 400 11960
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 5574 11930 5580 11932
rect 0 11870 5580 11930
rect 0 11840 400 11870
rect 5574 11868 5580 11870
rect 5644 11868 5650 11932
rect 9673 11930 9739 11933
rect 10133 11930 10199 11933
rect 9673 11928 10199 11930
rect 9673 11872 9678 11928
rect 9734 11872 10138 11928
rect 10194 11872 10199 11928
rect 9673 11870 10199 11872
rect 9673 11867 9739 11870
rect 10133 11867 10199 11870
rect 11697 11930 11763 11933
rect 12249 11930 12315 11933
rect 11697 11928 12315 11930
rect 11697 11872 11702 11928
rect 11758 11872 12254 11928
rect 12310 11872 12315 11928
rect 11697 11870 12315 11872
rect 11697 11867 11763 11870
rect 12249 11867 12315 11870
rect 15377 11930 15443 11933
rect 16021 11930 16087 11933
rect 17309 11930 17375 11933
rect 17861 11930 17927 11933
rect 18413 11930 18479 11933
rect 15377 11928 18479 11930
rect 15377 11872 15382 11928
rect 15438 11872 16026 11928
rect 16082 11872 17314 11928
rect 17370 11872 17866 11928
rect 17922 11872 18418 11928
rect 18474 11872 18479 11928
rect 15377 11870 18479 11872
rect 15377 11867 15443 11870
rect 16021 11867 16087 11870
rect 17309 11867 17375 11870
rect 17861 11867 17927 11870
rect 18413 11867 18479 11870
rect 8937 11794 9003 11797
rect 13721 11794 13787 11797
rect 8937 11792 13787 11794
rect 8937 11736 8942 11792
rect 8998 11736 13726 11792
rect 13782 11736 13787 11792
rect 8937 11734 13787 11736
rect 8937 11731 9003 11734
rect 13721 11731 13787 11734
rect 16062 11732 16068 11796
rect 16132 11794 16138 11796
rect 17493 11794 17559 11797
rect 16132 11792 17559 11794
rect 16132 11736 17498 11792
rect 17554 11736 17559 11792
rect 16132 11734 17559 11736
rect 16132 11732 16138 11734
rect 17493 11731 17559 11734
rect 20253 11794 20319 11797
rect 26969 11794 27035 11797
rect 20253 11792 27035 11794
rect 20253 11736 20258 11792
rect 20314 11736 26974 11792
rect 27030 11736 27035 11792
rect 20253 11734 27035 11736
rect 20253 11731 20319 11734
rect 26969 11731 27035 11734
rect 9305 11658 9371 11661
rect 10225 11658 10291 11661
rect 9305 11656 10291 11658
rect 9305 11600 9310 11656
rect 9366 11600 10230 11656
rect 10286 11600 10291 11656
rect 9305 11598 10291 11600
rect 9305 11595 9371 11598
rect 10225 11595 10291 11598
rect 11605 11658 11671 11661
rect 12249 11658 12315 11661
rect 11605 11656 12315 11658
rect 11605 11600 11610 11656
rect 11666 11600 12254 11656
rect 12310 11600 12315 11656
rect 11605 11598 12315 11600
rect 11605 11595 11671 11598
rect 12249 11595 12315 11598
rect 19885 11658 19951 11661
rect 22737 11658 22803 11661
rect 19885 11656 22803 11658
rect 19885 11600 19890 11656
rect 19946 11600 22742 11656
rect 22798 11600 22803 11656
rect 19885 11598 22803 11600
rect 19885 11595 19951 11598
rect 22737 11595 22803 11598
rect 5758 11460 5764 11524
rect 5828 11522 5834 11524
rect 5901 11522 5967 11525
rect 5828 11520 5967 11522
rect 5828 11464 5906 11520
rect 5962 11464 5967 11520
rect 5828 11462 5967 11464
rect 5828 11460 5834 11462
rect 5901 11459 5967 11462
rect 12065 11522 12131 11525
rect 16573 11522 16639 11525
rect 12065 11520 16639 11522
rect 12065 11464 12070 11520
rect 12126 11464 16578 11520
rect 16634 11464 16639 11520
rect 12065 11462 16639 11464
rect 12065 11459 12131 11462
rect 16573 11459 16639 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 8937 11386 9003 11389
rect 10409 11386 10475 11389
rect 8937 11384 10475 11386
rect 8937 11328 8942 11384
rect 8998 11328 10414 11384
rect 10470 11328 10475 11384
rect 8937 11326 10475 11328
rect 8937 11323 9003 11326
rect 10409 11323 10475 11326
rect 14825 11386 14891 11389
rect 17309 11386 17375 11389
rect 14825 11384 17375 11386
rect 14825 11328 14830 11384
rect 14886 11328 17314 11384
rect 17370 11328 17375 11384
rect 14825 11326 17375 11328
rect 14825 11323 14891 11326
rect 17309 11323 17375 11326
rect 9254 11188 9260 11252
rect 9324 11250 9330 11252
rect 9397 11250 9463 11253
rect 10133 11250 10199 11253
rect 14273 11250 14339 11253
rect 15377 11252 15443 11253
rect 15929 11252 15995 11253
rect 15326 11250 15332 11252
rect 9324 11248 14339 11250
rect 9324 11192 9402 11248
rect 9458 11192 10138 11248
rect 10194 11192 14278 11248
rect 14334 11192 14339 11248
rect 9324 11190 14339 11192
rect 15286 11190 15332 11250
rect 15396 11248 15443 11252
rect 15438 11192 15443 11248
rect 9324 11188 9330 11190
rect 9397 11187 9463 11190
rect 10133 11187 10199 11190
rect 14273 11187 14339 11190
rect 15326 11188 15332 11190
rect 15396 11188 15443 11192
rect 15878 11188 15884 11252
rect 15948 11250 15995 11252
rect 19241 11250 19307 11253
rect 21081 11250 21147 11253
rect 15948 11248 16040 11250
rect 15990 11192 16040 11248
rect 15948 11190 16040 11192
rect 19241 11248 21147 11250
rect 19241 11192 19246 11248
rect 19302 11192 21086 11248
rect 21142 11192 21147 11248
rect 19241 11190 21147 11192
rect 15948 11188 15995 11190
rect 15377 11187 15443 11188
rect 15929 11187 15995 11188
rect 19241 11187 19307 11190
rect 21081 11187 21147 11190
rect 1853 11114 1919 11117
rect 4153 11116 4219 11117
rect 2262 11114 2268 11116
rect 1853 11112 2268 11114
rect 1853 11056 1858 11112
rect 1914 11056 2268 11112
rect 1853 11054 2268 11056
rect 1853 11051 1919 11054
rect 2262 11052 2268 11054
rect 2332 11052 2338 11116
rect 4102 11114 4108 11116
rect 4062 11054 4108 11114
rect 4172 11112 4219 11116
rect 4214 11056 4219 11112
rect 4102 11052 4108 11054
rect 4172 11052 4219 11056
rect 4153 11051 4219 11052
rect 4337 11114 4403 11117
rect 4838 11114 4844 11116
rect 4337 11112 4844 11114
rect 4337 11056 4342 11112
rect 4398 11056 4844 11112
rect 4337 11054 4844 11056
rect 4337 11051 4403 11054
rect 4838 11052 4844 11054
rect 4908 11052 4914 11116
rect 9121 11114 9187 11117
rect 13445 11114 13511 11117
rect 9121 11112 13511 11114
rect 9121 11056 9126 11112
rect 9182 11056 13450 11112
rect 13506 11056 13511 11112
rect 9121 11054 13511 11056
rect 9121 11051 9187 11054
rect 13445 11051 13511 11054
rect 19609 11114 19675 11117
rect 25037 11114 25103 11117
rect 19609 11112 25103 11114
rect 19609 11056 19614 11112
rect 19670 11056 25042 11112
rect 25098 11056 25103 11112
rect 19609 11054 25103 11056
rect 19609 11051 19675 11054
rect 25037 11051 25103 11054
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 9857 10842 9923 10845
rect 12249 10842 12315 10845
rect 16113 10844 16179 10845
rect 19977 10844 20043 10845
rect 9857 10840 12315 10842
rect 9857 10784 9862 10840
rect 9918 10784 12254 10840
rect 12310 10784 12315 10840
rect 9857 10782 12315 10784
rect 9857 10779 9923 10782
rect 12249 10779 12315 10782
rect 16062 10780 16068 10844
rect 16132 10842 16179 10844
rect 16132 10840 16224 10842
rect 16174 10784 16224 10840
rect 16132 10782 16224 10784
rect 16132 10780 16179 10782
rect 19926 10780 19932 10844
rect 19996 10842 20043 10844
rect 19996 10840 20088 10842
rect 20038 10784 20088 10840
rect 19996 10782 20088 10784
rect 19996 10780 20043 10782
rect 16113 10779 16179 10780
rect 19977 10779 20043 10780
rect 7046 10644 7052 10708
rect 7116 10706 7122 10708
rect 7189 10706 7255 10709
rect 7116 10704 7255 10706
rect 7116 10648 7194 10704
rect 7250 10648 7255 10704
rect 7116 10646 7255 10648
rect 7116 10644 7122 10646
rect 7189 10643 7255 10646
rect 10041 10706 10107 10709
rect 10174 10706 10180 10708
rect 10041 10704 10180 10706
rect 10041 10648 10046 10704
rect 10102 10648 10180 10704
rect 10041 10646 10180 10648
rect 10041 10643 10107 10646
rect 10174 10644 10180 10646
rect 10244 10644 10250 10708
rect 13077 10706 13143 10709
rect 15929 10706 15995 10709
rect 13077 10704 15995 10706
rect 13077 10648 13082 10704
rect 13138 10648 15934 10704
rect 15990 10648 15995 10704
rect 13077 10646 15995 10648
rect 13077 10643 13143 10646
rect 15929 10643 15995 10646
rect 9213 10570 9279 10573
rect 13169 10570 13235 10573
rect 9213 10568 13235 10570
rect 9213 10512 9218 10568
rect 9274 10512 13174 10568
rect 13230 10512 13235 10568
rect 9213 10510 13235 10512
rect 9213 10507 9279 10510
rect 13169 10507 13235 10510
rect 2589 10434 2655 10437
rect 3141 10434 3207 10437
rect 2589 10432 3207 10434
rect 2589 10376 2594 10432
rect 2650 10376 3146 10432
rect 3202 10376 3207 10432
rect 2589 10374 3207 10376
rect 2589 10371 2655 10374
rect 3141 10371 3207 10374
rect 7598 10372 7604 10436
rect 7668 10434 7674 10436
rect 7833 10434 7899 10437
rect 7668 10432 7899 10434
rect 7668 10376 7838 10432
rect 7894 10376 7899 10432
rect 7668 10374 7899 10376
rect 7668 10372 7674 10374
rect 7833 10371 7899 10374
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 3734 10236 3740 10300
rect 3804 10298 3810 10300
rect 3969 10298 4035 10301
rect 3804 10296 4035 10298
rect 3804 10240 3974 10296
rect 4030 10240 4035 10296
rect 3804 10238 4035 10240
rect 3804 10236 3810 10238
rect 3969 10235 4035 10238
rect 10041 10298 10107 10301
rect 10358 10298 10364 10300
rect 10041 10296 10364 10298
rect 10041 10240 10046 10296
rect 10102 10240 10364 10296
rect 10041 10238 10364 10240
rect 10041 10235 10107 10238
rect 10358 10236 10364 10238
rect 10428 10236 10434 10300
rect 11973 10298 12039 10301
rect 15101 10298 15167 10301
rect 11973 10296 15167 10298
rect 11973 10240 11978 10296
rect 12034 10240 15106 10296
rect 15162 10240 15167 10296
rect 11973 10238 15167 10240
rect 11973 10235 12039 10238
rect 15101 10235 15167 10238
rect 11605 10162 11671 10165
rect 12157 10162 12223 10165
rect 16297 10164 16363 10165
rect 5904 10102 11346 10162
rect 5904 10029 5964 10102
rect 5022 9964 5028 10028
rect 5092 10026 5098 10028
rect 5901 10026 5967 10029
rect 11094 10026 11100 10028
rect 5092 10024 5967 10026
rect 5092 9968 5906 10024
rect 5962 9968 5967 10024
rect 5092 9966 5967 9968
rect 5092 9964 5098 9966
rect 5901 9963 5967 9966
rect 7606 9966 11100 10026
rect 0 9890 400 9920
rect 7606 9893 7666 9966
rect 11094 9964 11100 9966
rect 11164 9964 11170 10028
rect 11286 10026 11346 10102
rect 11605 10160 12223 10162
rect 11605 10104 11610 10160
rect 11666 10104 12162 10160
rect 12218 10104 12223 10160
rect 11605 10102 12223 10104
rect 11605 10099 11671 10102
rect 12157 10099 12223 10102
rect 15694 10100 15700 10164
rect 15764 10162 15770 10164
rect 16246 10162 16252 10164
rect 15764 10102 16252 10162
rect 16316 10162 16363 10164
rect 16316 10160 16408 10162
rect 16358 10104 16408 10160
rect 15764 10100 15770 10102
rect 16246 10100 16252 10102
rect 16316 10102 16408 10104
rect 16316 10100 16363 10102
rect 16297 10099 16363 10100
rect 13169 10026 13235 10029
rect 16757 10026 16823 10029
rect 17217 10026 17283 10029
rect 11286 10024 13235 10026
rect 11286 9968 13174 10024
rect 13230 9968 13235 10024
rect 11286 9966 13235 9968
rect 13169 9963 13235 9966
rect 14644 10024 17283 10026
rect 14644 9968 16762 10024
rect 16818 9968 17222 10024
rect 17278 9968 17283 10024
rect 14644 9966 17283 9968
rect 473 9890 539 9893
rect 5993 9892 6059 9893
rect 5942 9890 5948 9892
rect 0 9888 539 9890
rect 0 9832 478 9888
rect 534 9832 539 9888
rect 0 9830 539 9832
rect 5902 9830 5948 9890
rect 6012 9888 6059 9892
rect 6054 9832 6059 9888
rect 0 9800 400 9830
rect 473 9827 539 9830
rect 5942 9828 5948 9830
rect 6012 9828 6059 9832
rect 7606 9888 7715 9893
rect 7606 9832 7654 9888
rect 7710 9832 7715 9888
rect 7606 9830 7715 9832
rect 5993 9827 6059 9828
rect 7649 9827 7715 9830
rect 11973 9890 12039 9893
rect 14644 9890 14704 9966
rect 16757 9963 16823 9966
rect 17217 9963 17283 9966
rect 11973 9888 14704 9890
rect 11973 9832 11978 9888
rect 12034 9832 14704 9888
rect 11973 9830 14704 9832
rect 11973 9827 12039 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 1853 9754 1919 9757
rect 6545 9754 6611 9757
rect 1853 9752 6611 9754
rect 1853 9696 1858 9752
rect 1914 9696 6550 9752
rect 6606 9696 6611 9752
rect 1853 9694 6611 9696
rect 1853 9691 1919 9694
rect 6545 9691 6611 9694
rect 8518 9692 8524 9756
rect 8588 9754 8594 9756
rect 8937 9754 9003 9757
rect 9581 9754 9647 9757
rect 8588 9752 9647 9754
rect 8588 9696 8942 9752
rect 8998 9696 9586 9752
rect 9642 9696 9647 9752
rect 8588 9694 9647 9696
rect 8588 9692 8594 9694
rect 8937 9691 9003 9694
rect 9581 9691 9647 9694
rect 14365 9754 14431 9757
rect 22829 9754 22895 9757
rect 26509 9754 26575 9757
rect 14365 9752 14658 9754
rect 14365 9696 14370 9752
rect 14426 9696 14658 9752
rect 14365 9694 14658 9696
rect 14365 9691 14431 9694
rect 790 9556 796 9620
rect 860 9618 866 9620
rect 1393 9618 1459 9621
rect 860 9616 1459 9618
rect 860 9560 1398 9616
rect 1454 9560 1459 9616
rect 860 9558 1459 9560
rect 860 9556 866 9558
rect 1393 9555 1459 9558
rect 1761 9618 1827 9621
rect 3141 9618 3207 9621
rect 1761 9616 3207 9618
rect 1761 9560 1766 9616
rect 1822 9560 3146 9616
rect 3202 9560 3207 9616
rect 1761 9558 3207 9560
rect 1761 9555 1827 9558
rect 3141 9555 3207 9558
rect 7925 9618 7991 9621
rect 9397 9618 9463 9621
rect 7925 9616 9463 9618
rect 7925 9560 7930 9616
rect 7986 9560 9402 9616
rect 9458 9560 9463 9616
rect 7925 9558 9463 9560
rect 7925 9555 7991 9558
rect 9397 9555 9463 9558
rect 11237 9618 11303 9621
rect 11237 9616 13370 9618
rect 11237 9560 11242 9616
rect 11298 9560 13370 9616
rect 11237 9558 13370 9560
rect 11237 9555 11303 9558
rect 11605 9482 11671 9485
rect 12893 9482 12959 9485
rect 13118 9482 13124 9484
rect 11605 9480 12220 9482
rect 11605 9424 11610 9480
rect 11666 9424 12220 9480
rect 11605 9422 12220 9424
rect 11605 9419 11671 9422
rect 12160 9349 12220 9422
rect 12893 9480 13124 9482
rect 12893 9424 12898 9480
rect 12954 9424 13124 9480
rect 12893 9422 13124 9424
rect 12893 9419 12959 9422
rect 13118 9420 13124 9422
rect 13188 9420 13194 9484
rect 13310 9482 13370 9558
rect 14222 9556 14228 9620
rect 14292 9618 14298 9620
rect 14598 9618 14658 9694
rect 22829 9752 26575 9754
rect 22829 9696 22834 9752
rect 22890 9696 26514 9752
rect 26570 9696 26575 9752
rect 22829 9694 26575 9696
rect 22829 9691 22895 9694
rect 26509 9691 26575 9694
rect 15101 9618 15167 9621
rect 16481 9618 16547 9621
rect 14292 9616 16547 9618
rect 14292 9560 15106 9616
rect 15162 9560 16486 9616
rect 16542 9560 16547 9616
rect 14292 9558 16547 9560
rect 14292 9556 14298 9558
rect 15101 9555 15167 9558
rect 16481 9555 16547 9558
rect 15009 9482 15075 9485
rect 13310 9480 15075 9482
rect 13310 9424 15014 9480
rect 15070 9424 15075 9480
rect 13310 9422 15075 9424
rect 15009 9419 15075 9422
rect 15285 9482 15351 9485
rect 16113 9482 16179 9485
rect 17033 9482 17099 9485
rect 18137 9482 18203 9485
rect 15285 9480 18203 9482
rect 15285 9424 15290 9480
rect 15346 9424 16118 9480
rect 16174 9424 17038 9480
rect 17094 9424 18142 9480
rect 18198 9424 18203 9480
rect 15285 9422 18203 9424
rect 15285 9419 15351 9422
rect 16113 9419 16179 9422
rect 17033 9419 17099 9422
rect 18137 9419 18203 9422
rect 18873 9482 18939 9485
rect 24761 9482 24827 9485
rect 18873 9480 24827 9482
rect 18873 9424 18878 9480
rect 18934 9424 24766 9480
rect 24822 9424 24827 9480
rect 18873 9422 24827 9424
rect 18873 9419 18939 9422
rect 24761 9419 24827 9422
rect 12157 9344 12223 9349
rect 12157 9288 12162 9344
rect 12218 9288 12223 9344
rect 12157 9283 12223 9288
rect 13670 9284 13676 9348
rect 13740 9346 13746 9348
rect 15745 9346 15811 9349
rect 13740 9344 15811 9346
rect 13740 9288 15750 9344
rect 15806 9288 15811 9344
rect 13740 9286 15811 9288
rect 13740 9284 13746 9286
rect 15745 9283 15811 9286
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 1761 9210 1827 9213
rect 1894 9210 1900 9212
rect 1761 9208 1900 9210
rect 1761 9152 1766 9208
rect 1822 9152 1900 9208
rect 1761 9150 1900 9152
rect 1761 9147 1827 9150
rect 1894 9148 1900 9150
rect 1964 9148 1970 9212
rect 7230 9148 7236 9212
rect 7300 9210 7306 9212
rect 7649 9210 7715 9213
rect 7300 9208 7715 9210
rect 7300 9152 7654 9208
rect 7710 9152 7715 9208
rect 7300 9150 7715 9152
rect 7300 9148 7306 9150
rect 7649 9147 7715 9150
rect 15469 9210 15535 9213
rect 16481 9210 16547 9213
rect 15469 9208 16547 9210
rect 15469 9152 15474 9208
rect 15530 9152 16486 9208
rect 16542 9152 16547 9208
rect 15469 9150 16547 9152
rect 15469 9147 15535 9150
rect 16481 9147 16547 9150
rect 2262 9012 2268 9076
rect 2332 9074 2338 9076
rect 3233 9074 3299 9077
rect 27245 9074 27311 9077
rect 2332 9072 27311 9074
rect 2332 9016 3238 9072
rect 3294 9016 27250 9072
rect 27306 9016 27311 9072
rect 2332 9014 27311 9016
rect 2332 9012 2338 9014
rect 3233 9011 3299 9014
rect 27245 9011 27311 9014
rect 14457 8938 14523 8941
rect 16297 8938 16363 8941
rect 14457 8936 16363 8938
rect 14457 8880 14462 8936
rect 14518 8880 16302 8936
rect 16358 8880 16363 8936
rect 14457 8878 16363 8880
rect 14457 8875 14523 8878
rect 16297 8875 16363 8878
rect 22001 8938 22067 8941
rect 25221 8938 25287 8941
rect 22001 8936 25287 8938
rect 22001 8880 22006 8936
rect 22062 8880 25226 8936
rect 25282 8880 25287 8936
rect 22001 8878 25287 8880
rect 22001 8875 22067 8878
rect 25221 8875 25287 8878
rect 11329 8802 11395 8805
rect 12893 8802 12959 8805
rect 11329 8800 12959 8802
rect 11329 8744 11334 8800
rect 11390 8744 12898 8800
rect 12954 8744 12959 8800
rect 11329 8742 12959 8744
rect 11329 8739 11395 8742
rect 12893 8739 12959 8742
rect 22369 8802 22435 8805
rect 27153 8802 27219 8805
rect 22369 8800 27219 8802
rect 22369 8744 22374 8800
rect 22430 8744 27158 8800
rect 27214 8744 27219 8800
rect 22369 8742 27219 8744
rect 22369 8739 22435 8742
rect 27153 8739 27219 8742
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 9581 8666 9647 8669
rect 13445 8666 13511 8669
rect 14222 8666 14228 8668
rect 9581 8664 14228 8666
rect 9581 8608 9586 8664
rect 9642 8608 13450 8664
rect 13506 8608 14228 8664
rect 9581 8606 14228 8608
rect 9581 8603 9647 8606
rect 13445 8603 13511 8606
rect 14222 8604 14228 8606
rect 14292 8604 14298 8668
rect 17902 8604 17908 8668
rect 17972 8666 17978 8668
rect 20437 8666 20503 8669
rect 17972 8664 20503 8666
rect 17972 8608 20442 8664
rect 20498 8608 20503 8664
rect 17972 8606 20503 8608
rect 17972 8604 17978 8606
rect 20437 8603 20503 8606
rect 5533 8530 5599 8533
rect 16113 8530 16179 8533
rect 5533 8528 16179 8530
rect 5533 8472 5538 8528
rect 5594 8472 16118 8528
rect 16174 8472 16179 8528
rect 5533 8470 16179 8472
rect 5533 8467 5599 8470
rect 16113 8467 16179 8470
rect 18689 8530 18755 8533
rect 19517 8530 19583 8533
rect 21909 8530 21975 8533
rect 22093 8530 22159 8533
rect 18689 8528 19994 8530
rect 18689 8472 18694 8528
rect 18750 8472 19522 8528
rect 19578 8472 19994 8528
rect 18689 8470 19994 8472
rect 18689 8467 18755 8470
rect 19517 8467 19583 8470
rect 5533 8394 5599 8397
rect 6494 8394 6500 8396
rect 5533 8392 6500 8394
rect 5533 8336 5538 8392
rect 5594 8336 6500 8392
rect 5533 8334 6500 8336
rect 5533 8331 5599 8334
rect 6494 8332 6500 8334
rect 6564 8332 6570 8396
rect 9581 8394 9647 8397
rect 10777 8394 10843 8397
rect 9581 8392 10843 8394
rect 9581 8336 9586 8392
rect 9642 8336 10782 8392
rect 10838 8336 10843 8392
rect 9581 8334 10843 8336
rect 9581 8331 9647 8334
rect 10777 8331 10843 8334
rect 13118 8332 13124 8396
rect 13188 8394 13194 8396
rect 13445 8394 13511 8397
rect 13188 8392 13511 8394
rect 13188 8336 13450 8392
rect 13506 8336 13511 8392
rect 13188 8334 13511 8336
rect 13188 8332 13194 8334
rect 13445 8331 13511 8334
rect 14641 8394 14707 8397
rect 18689 8394 18755 8397
rect 14641 8392 18755 8394
rect 14641 8336 14646 8392
rect 14702 8336 18694 8392
rect 18750 8336 18755 8392
rect 14641 8334 18755 8336
rect 19934 8394 19994 8470
rect 21909 8528 22159 8530
rect 21909 8472 21914 8528
rect 21970 8472 22098 8528
rect 22154 8472 22159 8528
rect 21909 8470 22159 8472
rect 21909 8467 21975 8470
rect 22093 8467 22159 8470
rect 26325 8394 26391 8397
rect 19934 8392 26391 8394
rect 19934 8336 26330 8392
rect 26386 8336 26391 8392
rect 19934 8334 26391 8336
rect 14641 8331 14707 8334
rect 18689 8331 18755 8334
rect 26325 8331 26391 8334
rect 2313 8258 2379 8261
rect 2630 8258 2636 8260
rect 2313 8256 2636 8258
rect 2313 8200 2318 8256
rect 2374 8200 2636 8256
rect 2313 8198 2636 8200
rect 2313 8195 2379 8198
rect 2630 8196 2636 8198
rect 2700 8196 2706 8260
rect 14406 8196 14412 8260
rect 14476 8258 14482 8260
rect 15101 8258 15167 8261
rect 14476 8256 15167 8258
rect 14476 8200 15106 8256
rect 15162 8200 15167 8256
rect 14476 8198 15167 8200
rect 14476 8196 14482 8198
rect 15101 8195 15167 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 11838 8062 17234 8122
rect 3049 7986 3115 7989
rect 3918 7986 3924 7988
rect 3049 7984 3924 7986
rect 3049 7928 3054 7984
rect 3110 7928 3924 7984
rect 3049 7926 3924 7928
rect 3049 7923 3115 7926
rect 3918 7924 3924 7926
rect 3988 7924 3994 7988
rect 6177 7986 6243 7989
rect 7373 7986 7439 7989
rect 11838 7986 11898 8062
rect 6177 7984 11898 7986
rect 6177 7928 6182 7984
rect 6238 7928 7378 7984
rect 7434 7928 11898 7984
rect 6177 7926 11898 7928
rect 12341 7986 12407 7989
rect 12525 7986 12591 7989
rect 12341 7984 12591 7986
rect 12341 7928 12346 7984
rect 12402 7928 12530 7984
rect 12586 7928 12591 7984
rect 12341 7926 12591 7928
rect 17174 7986 17234 8062
rect 22921 7986 22987 7989
rect 17174 7984 22987 7986
rect 17174 7928 22926 7984
rect 22982 7928 22987 7984
rect 17174 7926 22987 7928
rect 6177 7923 6243 7926
rect 7373 7923 7439 7926
rect 12341 7923 12407 7926
rect 12525 7923 12591 7926
rect 22921 7923 22987 7926
rect 0 7850 400 7880
rect 13670 7850 13676 7852
rect 0 7790 13676 7850
rect 0 7760 400 7790
rect 13670 7788 13676 7790
rect 13740 7788 13746 7852
rect 19885 7850 19951 7853
rect 26601 7850 26667 7853
rect 19885 7848 26667 7850
rect 19885 7792 19890 7848
rect 19946 7792 26606 7848
rect 26662 7792 26667 7848
rect 19885 7790 26667 7792
rect 19885 7787 19951 7790
rect 26601 7787 26667 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 6913 7442 6979 7445
rect 7598 7442 7604 7444
rect 6913 7440 7604 7442
rect 6913 7384 6918 7440
rect 6974 7384 7604 7440
rect 6913 7382 7604 7384
rect 6913 7379 6979 7382
rect 7598 7380 7604 7382
rect 7668 7442 7674 7444
rect 17166 7442 17172 7444
rect 7668 7382 17172 7442
rect 7668 7380 7674 7382
rect 17166 7380 17172 7382
rect 17236 7380 17242 7444
rect 4705 7306 4771 7309
rect 5022 7306 5028 7308
rect 4705 7304 5028 7306
rect 4705 7248 4710 7304
rect 4766 7248 5028 7304
rect 4705 7246 5028 7248
rect 4705 7243 4771 7246
rect 5022 7244 5028 7246
rect 5092 7244 5098 7308
rect 6913 7306 6979 7309
rect 7414 7306 7420 7308
rect 6913 7304 7420 7306
rect 6913 7248 6918 7304
rect 6974 7248 7420 7304
rect 6913 7246 7420 7248
rect 6913 7243 6979 7246
rect 7414 7244 7420 7246
rect 7484 7306 7490 7308
rect 8109 7306 8175 7309
rect 7484 7304 8175 7306
rect 7484 7248 8114 7304
rect 8170 7248 8175 7304
rect 7484 7246 8175 7248
rect 7484 7244 7490 7246
rect 8109 7243 8175 7246
rect 11973 7306 12039 7309
rect 14733 7306 14799 7309
rect 11973 7304 14799 7306
rect 11973 7248 11978 7304
rect 12034 7248 14738 7304
rect 14794 7248 14799 7304
rect 11973 7246 14799 7248
rect 11973 7243 12039 7246
rect 14733 7243 14799 7246
rect 17861 7306 17927 7309
rect 19977 7306 20043 7309
rect 25681 7306 25747 7309
rect 17861 7304 25747 7306
rect 17861 7248 17866 7304
rect 17922 7248 19982 7304
rect 20038 7248 25686 7304
rect 25742 7248 25747 7304
rect 17861 7246 25747 7248
rect 17861 7243 17927 7246
rect 19977 7243 20043 7246
rect 25681 7243 25747 7246
rect 17217 7170 17283 7173
rect 17350 7170 17356 7172
rect 17217 7168 17356 7170
rect 17217 7112 17222 7168
rect 17278 7112 17356 7168
rect 17217 7110 17356 7112
rect 17217 7107 17283 7110
rect 17350 7108 17356 7110
rect 17420 7108 17426 7172
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 15469 7034 15535 7037
rect 17902 7034 17908 7036
rect 15469 7032 17908 7034
rect 15469 6976 15474 7032
rect 15530 6976 17908 7032
rect 15469 6974 17908 6976
rect 15469 6971 15535 6974
rect 17902 6972 17908 6974
rect 17972 6972 17978 7036
rect 12157 6898 12223 6901
rect 15326 6898 15332 6900
rect 12157 6896 15332 6898
rect 12157 6840 12162 6896
rect 12218 6840 15332 6896
rect 12157 6838 15332 6840
rect 12157 6835 12223 6838
rect 15326 6836 15332 6838
rect 15396 6836 15402 6900
rect 16481 6898 16547 6901
rect 17534 6898 17540 6900
rect 16481 6896 17540 6898
rect 16481 6840 16486 6896
rect 16542 6840 17540 6896
rect 16481 6838 17540 6840
rect 16481 6835 16547 6838
rect 17534 6836 17540 6838
rect 17604 6898 17610 6900
rect 24025 6898 24091 6901
rect 17604 6896 24091 6898
rect 17604 6840 24030 6896
rect 24086 6840 24091 6896
rect 17604 6838 24091 6840
rect 17604 6836 17610 6838
rect 24025 6835 24091 6838
rect 1158 6700 1164 6764
rect 1228 6762 1234 6764
rect 2957 6762 3023 6765
rect 1228 6760 3023 6762
rect 1228 6704 2962 6760
rect 3018 6704 3023 6760
rect 1228 6702 3023 6704
rect 1228 6700 1234 6702
rect 2957 6699 3023 6702
rect 9765 6762 9831 6765
rect 9990 6762 9996 6764
rect 9765 6760 9996 6762
rect 9765 6704 9770 6760
rect 9826 6704 9996 6760
rect 9765 6702 9996 6704
rect 9765 6699 9831 6702
rect 9990 6700 9996 6702
rect 10060 6700 10066 6764
rect 11237 6762 11303 6765
rect 12433 6762 12499 6765
rect 11237 6760 12499 6762
rect 11237 6704 11242 6760
rect 11298 6704 12438 6760
rect 12494 6704 12499 6760
rect 11237 6702 12499 6704
rect 11237 6699 11303 6702
rect 12433 6699 12499 6702
rect 15469 6762 15535 6765
rect 15694 6762 15700 6764
rect 15469 6760 15700 6762
rect 15469 6704 15474 6760
rect 15530 6704 15700 6760
rect 15469 6702 15700 6704
rect 15469 6699 15535 6702
rect 15694 6700 15700 6702
rect 15764 6700 15770 6764
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4613 6490 4679 6493
rect 5758 6490 5764 6492
rect 4613 6488 5764 6490
rect 4613 6432 4618 6488
rect 4674 6432 5764 6488
rect 4613 6430 5764 6432
rect 4613 6427 4679 6430
rect 5758 6428 5764 6430
rect 5828 6428 5834 6492
rect 15469 6490 15535 6493
rect 15745 6490 15811 6493
rect 15469 6488 15811 6490
rect 15469 6432 15474 6488
rect 15530 6432 15750 6488
rect 15806 6432 15811 6488
rect 15469 6430 15811 6432
rect 15469 6427 15535 6430
rect 15745 6427 15811 6430
rect 5942 6292 5948 6356
rect 6012 6354 6018 6356
rect 6177 6354 6243 6357
rect 19057 6354 19123 6357
rect 6012 6352 19123 6354
rect 6012 6296 6182 6352
rect 6238 6296 19062 6352
rect 19118 6296 19123 6352
rect 6012 6294 19123 6296
rect 6012 6292 6018 6294
rect 6177 6291 6243 6294
rect 19057 6291 19123 6294
rect 23381 6354 23447 6357
rect 26417 6354 26483 6357
rect 23381 6352 26483 6354
rect 23381 6296 23386 6352
rect 23442 6296 26422 6352
rect 26478 6296 26483 6352
rect 23381 6294 26483 6296
rect 23381 6291 23447 6294
rect 26417 6291 26483 6294
rect 4153 6220 4219 6221
rect 4102 6218 4108 6220
rect 4062 6158 4108 6218
rect 4172 6218 4219 6220
rect 5441 6218 5507 6221
rect 4172 6216 5507 6218
rect 4214 6160 5446 6216
rect 5502 6160 5507 6216
rect 4102 6156 4108 6158
rect 4172 6158 5507 6160
rect 4172 6156 4219 6158
rect 4153 6155 4219 6156
rect 5441 6155 5507 6158
rect 15193 6218 15259 6221
rect 15837 6218 15903 6221
rect 15193 6216 15903 6218
rect 15193 6160 15198 6216
rect 15254 6160 15842 6216
rect 15898 6160 15903 6216
rect 15193 6158 15903 6160
rect 15193 6155 15259 6158
rect 15837 6155 15903 6158
rect 16021 6218 16087 6221
rect 20989 6218 21055 6221
rect 16021 6216 21055 6218
rect 16021 6160 16026 6216
rect 16082 6160 20994 6216
rect 21050 6160 21055 6216
rect 16021 6158 21055 6160
rect 16021 6155 16087 6158
rect 20989 6155 21055 6158
rect 4797 6082 4863 6085
rect 9397 6082 9463 6085
rect 4797 6080 9463 6082
rect 4797 6024 4802 6080
rect 4858 6024 9402 6080
rect 9458 6024 9463 6080
rect 4797 6022 9463 6024
rect 4797 6019 4863 6022
rect 9397 6019 9463 6022
rect 13169 6082 13235 6085
rect 13813 6082 13879 6085
rect 13169 6080 13879 6082
rect 13169 6024 13174 6080
rect 13230 6024 13818 6080
rect 13874 6024 13879 6080
rect 13169 6022 13879 6024
rect 13169 6019 13235 6022
rect 13813 6019 13879 6022
rect 14273 6082 14339 6085
rect 16021 6082 16087 6085
rect 14273 6080 16087 6082
rect 14273 6024 14278 6080
rect 14334 6024 16026 6080
rect 16082 6024 16087 6080
rect 14273 6022 16087 6024
rect 14273 6019 14339 6022
rect 16021 6019 16087 6022
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 7005 5946 7071 5949
rect 7230 5946 7236 5948
rect 7005 5944 7236 5946
rect 7005 5888 7010 5944
rect 7066 5888 7236 5944
rect 7005 5886 7236 5888
rect 7005 5883 7071 5886
rect 7230 5884 7236 5886
rect 7300 5884 7306 5948
rect 13353 5946 13419 5949
rect 16573 5946 16639 5949
rect 13353 5944 16639 5946
rect 13353 5888 13358 5944
rect 13414 5888 16578 5944
rect 16634 5888 16639 5944
rect 13353 5886 16639 5888
rect 13353 5883 13419 5886
rect 16573 5883 16639 5886
rect 0 5810 400 5840
rect 473 5810 539 5813
rect 0 5808 539 5810
rect 0 5752 478 5808
rect 534 5752 539 5808
rect 0 5750 539 5752
rect 0 5720 400 5750
rect 473 5747 539 5750
rect 1853 5810 1919 5813
rect 4981 5810 5047 5813
rect 5206 5810 5212 5812
rect 1853 5808 2790 5810
rect 1853 5752 1858 5808
rect 1914 5752 2790 5808
rect 1853 5750 2790 5752
rect 1853 5747 1919 5750
rect 2730 5674 2790 5750
rect 4981 5808 5212 5810
rect 4981 5752 4986 5808
rect 5042 5752 5212 5808
rect 4981 5750 5212 5752
rect 4981 5747 5047 5750
rect 5206 5748 5212 5750
rect 5276 5748 5282 5812
rect 5758 5748 5764 5812
rect 5828 5810 5834 5812
rect 18689 5810 18755 5813
rect 5828 5808 18755 5810
rect 5828 5752 18694 5808
rect 18750 5752 18755 5808
rect 5828 5750 18755 5752
rect 5828 5748 5834 5750
rect 18689 5747 18755 5750
rect 15193 5674 15259 5677
rect 22318 5674 22324 5676
rect 2730 5672 22324 5674
rect 2730 5616 15198 5672
rect 15254 5616 22324 5672
rect 2730 5614 22324 5616
rect 15193 5611 15259 5614
rect 22318 5612 22324 5614
rect 22388 5612 22394 5676
rect 3509 5538 3575 5541
rect 6729 5538 6795 5541
rect 3509 5536 6795 5538
rect 3509 5480 3514 5536
rect 3570 5480 6734 5536
rect 6790 5480 6795 5536
rect 3509 5478 6795 5480
rect 3509 5475 3575 5478
rect 6729 5475 6795 5478
rect 12985 5538 13051 5541
rect 13721 5538 13787 5541
rect 14273 5538 14339 5541
rect 12985 5536 14339 5538
rect 12985 5480 12990 5536
rect 13046 5480 13726 5536
rect 13782 5480 14278 5536
rect 14334 5480 14339 5536
rect 12985 5478 14339 5480
rect 12985 5475 13051 5478
rect 13721 5475 13787 5478
rect 14273 5475 14339 5478
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 6637 5266 6703 5269
rect 27705 5266 27771 5269
rect 6637 5264 27771 5266
rect 6637 5208 6642 5264
rect 6698 5208 27710 5264
rect 27766 5208 27771 5264
rect 6637 5206 27771 5208
rect 6637 5203 6703 5206
rect 27705 5203 27771 5206
rect 5809 5130 5875 5133
rect 24117 5130 24183 5133
rect 5809 5128 24183 5130
rect 5809 5072 5814 5128
rect 5870 5072 24122 5128
rect 24178 5072 24183 5128
rect 5809 5070 24183 5072
rect 5809 5067 5875 5070
rect 24117 5067 24183 5070
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 4838 4796 4844 4860
rect 4908 4858 4914 4860
rect 4981 4858 5047 4861
rect 4908 4856 5047 4858
rect 4908 4800 4986 4856
rect 5042 4800 5047 4856
rect 4908 4798 5047 4800
rect 4908 4796 4914 4798
rect 4981 4795 5047 4798
rect 7373 4722 7439 4725
rect 27613 4722 27679 4725
rect 7373 4720 27679 4722
rect 7373 4664 7378 4720
rect 7434 4664 27618 4720
rect 27674 4664 27679 4720
rect 7373 4662 27679 4664
rect 7373 4659 7439 4662
rect 27613 4659 27679 4662
rect 17166 4524 17172 4588
rect 17236 4586 17242 4588
rect 27337 4586 27403 4589
rect 17236 4584 27403 4586
rect 17236 4528 27342 4584
rect 27398 4528 27403 4584
rect 17236 4526 27403 4528
rect 17236 4524 17242 4526
rect 27337 4523 27403 4526
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 17902 4116 17908 4180
rect 17972 4178 17978 4180
rect 22369 4178 22435 4181
rect 23381 4178 23447 4181
rect 17972 4176 23447 4178
rect 17972 4120 22374 4176
rect 22430 4120 23386 4176
rect 23442 4120 23447 4176
rect 17972 4118 23447 4120
rect 17972 4116 17978 4118
rect 22369 4115 22435 4118
rect 23381 4115 23447 4118
rect 5073 4042 5139 4045
rect 27337 4042 27403 4045
rect 5073 4040 27403 4042
rect 5073 3984 5078 4040
rect 5134 3984 27342 4040
rect 27398 3984 27403 4040
rect 5073 3982 27403 3984
rect 5073 3979 5139 3982
rect 27337 3979 27403 3982
rect 5625 3908 5691 3909
rect 5574 3906 5580 3908
rect 5534 3846 5580 3906
rect 5644 3904 5691 3908
rect 5686 3848 5691 3904
rect 5574 3844 5580 3846
rect 5644 3844 5691 3848
rect 5625 3843 5691 3844
rect 20437 3906 20503 3909
rect 23381 3906 23447 3909
rect 20437 3904 23447 3906
rect 20437 3848 20442 3904
rect 20498 3848 23386 3904
rect 23442 3848 23447 3904
rect 20437 3846 23447 3848
rect 20437 3843 20503 3846
rect 23381 3843 23447 3846
rect 4419 3840 4735 3841
rect 0 3770 400 3800
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 473 3770 539 3773
rect 0 3768 539 3770
rect 0 3712 478 3768
rect 534 3712 539 3768
rect 0 3710 539 3712
rect 0 3680 400 3710
rect 473 3707 539 3710
rect 19793 3634 19859 3637
rect 25773 3634 25839 3637
rect 19793 3632 25839 3634
rect 19793 3576 19798 3632
rect 19854 3576 25778 3632
rect 25834 3576 25839 3632
rect 19793 3574 25839 3576
rect 19793 3571 19859 3574
rect 25773 3571 25839 3574
rect 5717 3500 5783 3501
rect 5717 3498 5764 3500
rect 5672 3496 5764 3498
rect 5672 3440 5722 3496
rect 5672 3438 5764 3440
rect 5717 3436 5764 3438
rect 5828 3436 5834 3500
rect 20437 3498 20503 3501
rect 21909 3498 21975 3501
rect 20437 3496 21975 3498
rect 20437 3440 20442 3496
rect 20498 3440 21914 3496
rect 21970 3440 21975 3496
rect 20437 3438 21975 3440
rect 5717 3435 5783 3436
rect 20437 3435 20503 3438
rect 21909 3435 21975 3438
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 5349 3090 5415 3093
rect 18781 3090 18847 3093
rect 5349 3088 18847 3090
rect 5349 3032 5354 3088
rect 5410 3032 18786 3088
rect 18842 3032 18847 3088
rect 5349 3030 18847 3032
rect 5349 3027 5415 3030
rect 18781 3027 18847 3030
rect 13445 2954 13511 2957
rect 26233 2954 26299 2957
rect 13445 2952 26299 2954
rect 13445 2896 13450 2952
rect 13506 2896 26238 2952
rect 26294 2896 26299 2952
rect 13445 2894 26299 2896
rect 13445 2891 13511 2894
rect 26233 2891 26299 2894
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 19425 2682 19491 2685
rect 21909 2682 21975 2685
rect 19425 2680 21975 2682
rect 19425 2624 19430 2680
rect 19486 2624 21914 2680
rect 21970 2624 21975 2680
rect 19425 2622 21975 2624
rect 19425 2619 19491 2622
rect 21909 2619 21975 2622
rect 974 2484 980 2548
rect 1044 2546 1050 2548
rect 1669 2546 1735 2549
rect 1044 2544 1735 2546
rect 1044 2488 1674 2544
rect 1730 2488 1735 2544
rect 1044 2486 1735 2488
rect 1044 2484 1050 2486
rect 1669 2483 1735 2486
rect 8201 2546 8267 2549
rect 25681 2546 25747 2549
rect 8201 2544 25747 2546
rect 8201 2488 8206 2544
rect 8262 2488 25686 2544
rect 25742 2488 25747 2544
rect 8201 2486 25747 2488
rect 8201 2483 8267 2486
rect 25681 2483 25747 2486
rect 4797 2410 4863 2413
rect 26509 2410 26575 2413
rect 4797 2408 26575 2410
rect 4797 2352 4802 2408
rect 4858 2352 26514 2408
rect 26570 2352 26575 2408
rect 4797 2350 26575 2352
rect 4797 2347 4863 2350
rect 26509 2347 26575 2350
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 21173 2138 21239 2141
rect 21541 2138 21607 2141
rect 21173 2136 21607 2138
rect 21173 2080 21178 2136
rect 21234 2080 21546 2136
rect 21602 2080 21607 2136
rect 21173 2078 21607 2080
rect 21173 2075 21239 2078
rect 21541 2075 21607 2078
rect 54 1940 60 2004
rect 124 2002 130 2004
rect 2589 2002 2655 2005
rect 26325 2002 26391 2005
rect 124 1942 536 2002
rect 124 1940 130 1942
rect 0 1730 400 1760
rect 476 1730 536 1942
rect 2589 2000 26391 2002
rect 2589 1944 2594 2000
rect 2650 1944 26330 2000
rect 26386 1944 26391 2000
rect 2589 1942 26391 1944
rect 2589 1939 2655 1942
rect 26325 1939 26391 1942
rect 0 1670 536 1730
rect 0 1640 400 1670
rect 4419 1664 4735 1665
rect 4419 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4735 1664
rect 4419 1599 4735 1600
rect 11365 1664 11681 1665
rect 11365 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11681 1664
rect 11365 1599 11681 1600
rect 18311 1664 18627 1665
rect 18311 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18627 1664
rect 18311 1599 18627 1600
rect 25257 1664 25573 1665
rect 25257 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25573 1664
rect 25257 1599 25573 1600
rect 17309 1594 17375 1597
rect 17861 1594 17927 1597
rect 17309 1592 17927 1594
rect 17309 1536 17314 1592
rect 17370 1536 17866 1592
rect 17922 1536 17927 1592
rect 17309 1534 17927 1536
rect 17309 1531 17375 1534
rect 17861 1531 17927 1534
rect 8201 1322 8267 1325
rect 13486 1322 13492 1324
rect 8201 1320 13492 1322
rect 8201 1264 8206 1320
rect 8262 1264 13492 1320
rect 8201 1262 13492 1264
rect 8201 1259 8267 1262
rect 13486 1260 13492 1262
rect 13556 1260 13562 1324
rect 7892 1120 8208 1121
rect 7892 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8208 1120
rect 7892 1055 8208 1056
rect 14838 1120 15154 1121
rect 14838 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15154 1120
rect 14838 1055 15154 1056
rect 21784 1120 22100 1121
rect 21784 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22100 1120
rect 21784 1055 22100 1056
rect 28730 1120 29046 1121
rect 28730 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29046 1120
rect 28730 1055 29046 1056
<< via3 >>
rect 7898 32668 7962 32672
rect 7898 32612 7902 32668
rect 7902 32612 7958 32668
rect 7958 32612 7962 32668
rect 7898 32608 7962 32612
rect 7978 32668 8042 32672
rect 7978 32612 7982 32668
rect 7982 32612 8038 32668
rect 8038 32612 8042 32668
rect 7978 32608 8042 32612
rect 8058 32668 8122 32672
rect 8058 32612 8062 32668
rect 8062 32612 8118 32668
rect 8118 32612 8122 32668
rect 8058 32608 8122 32612
rect 8138 32668 8202 32672
rect 8138 32612 8142 32668
rect 8142 32612 8198 32668
rect 8198 32612 8202 32668
rect 8138 32608 8202 32612
rect 14844 32668 14908 32672
rect 14844 32612 14848 32668
rect 14848 32612 14904 32668
rect 14904 32612 14908 32668
rect 14844 32608 14908 32612
rect 14924 32668 14988 32672
rect 14924 32612 14928 32668
rect 14928 32612 14984 32668
rect 14984 32612 14988 32668
rect 14924 32608 14988 32612
rect 15004 32668 15068 32672
rect 15004 32612 15008 32668
rect 15008 32612 15064 32668
rect 15064 32612 15068 32668
rect 15004 32608 15068 32612
rect 15084 32668 15148 32672
rect 15084 32612 15088 32668
rect 15088 32612 15144 32668
rect 15144 32612 15148 32668
rect 15084 32608 15148 32612
rect 21790 32668 21854 32672
rect 21790 32612 21794 32668
rect 21794 32612 21850 32668
rect 21850 32612 21854 32668
rect 21790 32608 21854 32612
rect 21870 32668 21934 32672
rect 21870 32612 21874 32668
rect 21874 32612 21930 32668
rect 21930 32612 21934 32668
rect 21870 32608 21934 32612
rect 21950 32668 22014 32672
rect 21950 32612 21954 32668
rect 21954 32612 22010 32668
rect 22010 32612 22014 32668
rect 21950 32608 22014 32612
rect 22030 32668 22094 32672
rect 22030 32612 22034 32668
rect 22034 32612 22090 32668
rect 22090 32612 22094 32668
rect 22030 32608 22094 32612
rect 28736 32668 28800 32672
rect 28736 32612 28740 32668
rect 28740 32612 28796 32668
rect 28796 32612 28800 32668
rect 28736 32608 28800 32612
rect 28816 32668 28880 32672
rect 28816 32612 28820 32668
rect 28820 32612 28876 32668
rect 28876 32612 28880 32668
rect 28816 32608 28880 32612
rect 28896 32668 28960 32672
rect 28896 32612 28900 32668
rect 28900 32612 28956 32668
rect 28956 32612 28960 32668
rect 28896 32608 28960 32612
rect 28976 32668 29040 32672
rect 28976 32612 28980 32668
rect 28980 32612 29036 32668
rect 29036 32612 29040 32668
rect 28976 32608 29040 32612
rect 4425 32124 4489 32128
rect 4425 32068 4429 32124
rect 4429 32068 4485 32124
rect 4485 32068 4489 32124
rect 4425 32064 4489 32068
rect 4505 32124 4569 32128
rect 4505 32068 4509 32124
rect 4509 32068 4565 32124
rect 4565 32068 4569 32124
rect 4505 32064 4569 32068
rect 4585 32124 4649 32128
rect 4585 32068 4589 32124
rect 4589 32068 4645 32124
rect 4645 32068 4649 32124
rect 4585 32064 4649 32068
rect 4665 32124 4729 32128
rect 4665 32068 4669 32124
rect 4669 32068 4725 32124
rect 4725 32068 4729 32124
rect 4665 32064 4729 32068
rect 11371 32124 11435 32128
rect 11371 32068 11375 32124
rect 11375 32068 11431 32124
rect 11431 32068 11435 32124
rect 11371 32064 11435 32068
rect 11451 32124 11515 32128
rect 11451 32068 11455 32124
rect 11455 32068 11511 32124
rect 11511 32068 11515 32124
rect 11451 32064 11515 32068
rect 11531 32124 11595 32128
rect 11531 32068 11535 32124
rect 11535 32068 11591 32124
rect 11591 32068 11595 32124
rect 11531 32064 11595 32068
rect 11611 32124 11675 32128
rect 11611 32068 11615 32124
rect 11615 32068 11671 32124
rect 11671 32068 11675 32124
rect 11611 32064 11675 32068
rect 18317 32124 18381 32128
rect 18317 32068 18321 32124
rect 18321 32068 18377 32124
rect 18377 32068 18381 32124
rect 18317 32064 18381 32068
rect 18397 32124 18461 32128
rect 18397 32068 18401 32124
rect 18401 32068 18457 32124
rect 18457 32068 18461 32124
rect 18397 32064 18461 32068
rect 18477 32124 18541 32128
rect 18477 32068 18481 32124
rect 18481 32068 18537 32124
rect 18537 32068 18541 32124
rect 18477 32064 18541 32068
rect 18557 32124 18621 32128
rect 18557 32068 18561 32124
rect 18561 32068 18617 32124
rect 18617 32068 18621 32124
rect 18557 32064 18621 32068
rect 25263 32124 25327 32128
rect 25263 32068 25267 32124
rect 25267 32068 25323 32124
rect 25323 32068 25327 32124
rect 25263 32064 25327 32068
rect 25343 32124 25407 32128
rect 25343 32068 25347 32124
rect 25347 32068 25403 32124
rect 25403 32068 25407 32124
rect 25343 32064 25407 32068
rect 25423 32124 25487 32128
rect 25423 32068 25427 32124
rect 25427 32068 25483 32124
rect 25483 32068 25487 32124
rect 25423 32064 25487 32068
rect 25503 32124 25567 32128
rect 25503 32068 25507 32124
rect 25507 32068 25563 32124
rect 25563 32068 25567 32124
rect 25503 32064 25567 32068
rect 14596 31724 14660 31788
rect 15884 31588 15948 31652
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 17172 30772 17236 30836
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 10548 29956 10612 30020
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 17908 28596 17972 28660
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 5212 28460 5276 28524
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 17356 28188 17420 28252
rect 17172 28052 17236 28116
rect 5580 27780 5644 27844
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 19380 27780 19444 27844
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 14412 27704 14476 27708
rect 14412 27648 14426 27704
rect 14426 27648 14476 27704
rect 14412 27644 14476 27648
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 13308 26692 13372 26756
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 5212 26556 5276 26620
rect 14044 26616 14108 26620
rect 14044 26560 14058 26616
rect 14058 26560 14108 26616
rect 14044 26556 14108 26560
rect 6684 26480 6748 26484
rect 6684 26424 6698 26480
rect 6698 26424 6748 26480
rect 6684 26420 6748 26424
rect 5212 26344 5276 26348
rect 5212 26288 5262 26344
rect 5262 26288 5276 26344
rect 5212 26284 5276 26288
rect 9260 26284 9324 26348
rect 8340 26148 8404 26212
rect 10364 26148 10428 26212
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 4108 26012 4172 26076
rect 22324 26148 22388 26212
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 17908 26012 17972 26076
rect 19380 25876 19444 25940
rect 9812 25800 9876 25804
rect 9812 25744 9826 25800
rect 9826 25744 9876 25800
rect 9812 25740 9876 25744
rect 7604 25604 7668 25668
rect 18828 25604 18892 25668
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 14596 25468 14660 25532
rect 3188 25332 3252 25396
rect 22324 25196 22388 25260
rect 15332 25060 15396 25124
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 5396 24984 5460 24988
rect 5396 24928 5410 24984
rect 5410 24928 5460 24984
rect 5396 24924 5460 24928
rect 13124 24984 13188 24988
rect 13124 24928 13174 24984
rect 13174 24928 13188 24984
rect 13124 24924 13188 24928
rect 16068 24924 16132 24988
rect 18828 24924 18892 24988
rect 15884 24652 15948 24716
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 6316 23972 6380 24036
rect 10364 23972 10428 24036
rect 13124 23972 13188 24036
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 7052 23836 7116 23900
rect 12020 23836 12084 23900
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 19012 24032 19076 24036
rect 19012 23976 19062 24032
rect 19062 23976 19076 24032
rect 19012 23972 19076 23976
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4292 23624 4356 23628
rect 4292 23568 4342 23624
rect 4342 23568 4356 23624
rect 4292 23564 4356 23568
rect 8340 23564 8404 23628
rect 9444 23564 9508 23628
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 10548 23216 10612 23220
rect 10548 23160 10562 23216
rect 10562 23160 10612 23216
rect 10548 23156 10612 23160
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 6684 23020 6748 23084
rect 16436 22884 16500 22948
rect 19380 22884 19444 22948
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 5580 22612 5644 22676
rect 17356 22612 17420 22676
rect 18092 22612 18156 22676
rect 7604 22476 7668 22540
rect 19196 22340 19260 22404
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 14596 22204 14660 22268
rect 16068 21932 16132 21996
rect 6316 21796 6380 21860
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 19012 21660 19076 21724
rect 3188 21524 3252 21588
rect 15332 21388 15396 21452
rect 18828 21388 18892 21452
rect 20300 21388 20364 21452
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 5212 21116 5276 21180
rect 5212 21040 5276 21044
rect 5212 20984 5226 21040
rect 5226 20984 5276 21040
rect 5212 20980 5276 20984
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 6684 21040 6748 21044
rect 6684 20984 6698 21040
rect 6698 20984 6748 21040
rect 6684 20980 6748 20984
rect 19196 20980 19260 21044
rect 8524 20768 8588 20772
rect 8524 20712 8538 20768
rect 8538 20712 8588 20768
rect 8524 20708 8588 20712
rect 12020 20708 12084 20772
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 19380 20572 19444 20636
rect 9260 20436 9324 20500
rect 1164 20300 1228 20364
rect 4108 20224 4172 20228
rect 4108 20168 4158 20224
rect 4158 20168 4172 20224
rect 4108 20164 4172 20168
rect 7052 20224 7116 20228
rect 7052 20168 7102 20224
rect 7102 20168 7116 20224
rect 7052 20164 7116 20168
rect 20484 20164 20548 20228
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 13676 20028 13740 20092
rect 5396 19892 5460 19956
rect 14228 19892 14292 19956
rect 14596 19892 14660 19956
rect 15516 19892 15580 19956
rect 796 19620 860 19684
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 5396 19484 5460 19548
rect 14596 19756 14660 19820
rect 17908 19680 17972 19684
rect 17908 19624 17958 19680
rect 17958 19624 17972 19680
rect 17908 19620 17972 19624
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 6500 19484 6564 19548
rect 12204 19484 12268 19548
rect 13492 19348 13556 19412
rect 14412 19348 14476 19412
rect 16620 19408 16684 19412
rect 16620 19352 16670 19408
rect 16670 19352 16684 19408
rect 16620 19348 16684 19352
rect 13308 19272 13372 19276
rect 13308 19216 13322 19272
rect 13322 19216 13372 19272
rect 13308 19212 13372 19216
rect 17908 19076 17972 19140
rect 19380 19136 19444 19140
rect 19380 19080 19430 19136
rect 19430 19080 19444 19136
rect 19380 19076 19444 19080
rect 20116 19136 20180 19140
rect 20116 19080 20166 19136
rect 20166 19080 20180 19136
rect 20116 19076 20180 19080
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 16068 18940 16132 19004
rect 22324 18804 22388 18868
rect 15884 18668 15948 18732
rect 20300 18668 20364 18732
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4292 18260 4356 18324
rect 7604 18124 7668 18188
rect 1900 17988 1964 18052
rect 11836 18048 11900 18052
rect 11836 17992 11886 18048
rect 11886 17992 11900 18048
rect 11836 17988 11900 17992
rect 14412 17988 14476 18052
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 5028 17912 5092 17916
rect 5028 17856 5042 17912
rect 5042 17856 5092 17912
rect 5028 17852 5092 17856
rect 5212 17852 5276 17916
rect 13124 17852 13188 17916
rect 14044 17912 14108 17916
rect 14044 17856 14058 17912
rect 14058 17856 14108 17912
rect 14044 17852 14108 17856
rect 16252 17852 16316 17916
rect 16436 17912 16500 17916
rect 19748 17988 19812 18052
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 16436 17856 16450 17912
rect 16450 17856 16500 17912
rect 16436 17852 16500 17856
rect 9996 17716 10060 17780
rect 18092 17716 18156 17780
rect 12204 17444 12268 17508
rect 19564 17504 19628 17508
rect 19564 17448 19614 17504
rect 19614 17448 19628 17504
rect 19564 17444 19628 17448
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 2268 17172 2332 17236
rect 13124 17172 13188 17236
rect 19380 16900 19444 16964
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 3740 16688 3804 16692
rect 3740 16632 3754 16688
rect 3754 16632 3804 16688
rect 3740 16628 3804 16632
rect 4292 16628 4356 16692
rect 6684 16492 6748 16556
rect 18828 16356 18892 16420
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 7420 16220 7484 16284
rect 6500 16144 6564 16148
rect 6500 16088 6514 16144
rect 6514 16088 6564 16144
rect 6500 16084 6564 16088
rect 9812 16084 9876 16148
rect 11836 16084 11900 16148
rect 19380 16144 19444 16148
rect 19380 16088 19394 16144
rect 19394 16088 19444 16144
rect 19380 16084 19444 16088
rect 13492 16008 13556 16012
rect 13492 15952 13542 16008
rect 13542 15952 13556 16008
rect 13492 15948 13556 15952
rect 15332 15812 15396 15876
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7052 15404 7116 15468
rect 16620 15404 16684 15468
rect 2636 15268 2700 15332
rect 13676 15268 13740 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 7236 15132 7300 15196
rect 20484 15132 20548 15196
rect 16068 14860 16132 14924
rect 14412 14724 14476 14788
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 19932 14512 19996 14516
rect 19932 14456 19982 14512
rect 19982 14456 19996 14512
rect 19932 14452 19996 14456
rect 980 14316 1044 14380
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 11100 13908 11164 13972
rect 14228 13908 14292 13972
rect 9444 13772 9508 13836
rect 13492 13832 13556 13836
rect 13492 13776 13542 13832
rect 13542 13776 13556 13832
rect 13492 13772 13556 13776
rect 12020 13636 12084 13700
rect 20116 13636 20180 13700
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 9260 13500 9324 13564
rect 15516 13500 15580 13564
rect 14412 13364 14476 13428
rect 19564 13364 19628 13428
rect 17356 13092 17420 13156
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4292 12880 4356 12884
rect 4292 12824 4342 12880
rect 4342 12824 4356 12880
rect 4292 12820 4356 12824
rect 5212 12820 5276 12884
rect 14596 12820 14660 12884
rect 7604 12744 7668 12748
rect 7604 12688 7618 12744
rect 7618 12688 7668 12744
rect 7604 12684 7668 12688
rect 10180 12744 10244 12748
rect 10180 12688 10230 12744
rect 10230 12688 10244 12744
rect 10180 12684 10244 12688
rect 17908 12684 17972 12748
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 60 12412 124 12476
rect 5396 12412 5460 12476
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 17540 12472 17604 12476
rect 17540 12416 17554 12472
rect 17554 12416 17604 12472
rect 17540 12412 17604 12416
rect 15332 12276 15396 12340
rect 19748 12336 19812 12340
rect 19748 12280 19798 12336
rect 19798 12280 19812 12336
rect 19748 12276 19812 12280
rect 3924 12140 3988 12204
rect 2268 12004 2332 12068
rect 10364 12004 10428 12068
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 5580 11868 5644 11932
rect 16068 11732 16132 11796
rect 5764 11460 5828 11524
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 9260 11188 9324 11252
rect 15332 11248 15396 11252
rect 15332 11192 15382 11248
rect 15382 11192 15396 11248
rect 15332 11188 15396 11192
rect 15884 11248 15948 11252
rect 15884 11192 15934 11248
rect 15934 11192 15948 11248
rect 15884 11188 15948 11192
rect 2268 11052 2332 11116
rect 4108 11112 4172 11116
rect 4108 11056 4158 11112
rect 4158 11056 4172 11112
rect 4108 11052 4172 11056
rect 4844 11052 4908 11116
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 16068 10840 16132 10844
rect 16068 10784 16118 10840
rect 16118 10784 16132 10840
rect 16068 10780 16132 10784
rect 19932 10840 19996 10844
rect 19932 10784 19982 10840
rect 19982 10784 19996 10840
rect 19932 10780 19996 10784
rect 7052 10644 7116 10708
rect 10180 10644 10244 10708
rect 7604 10372 7668 10436
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 3740 10236 3804 10300
rect 10364 10236 10428 10300
rect 5028 9964 5092 10028
rect 11100 9964 11164 10028
rect 15700 10100 15764 10164
rect 16252 10160 16316 10164
rect 16252 10104 16302 10160
rect 16302 10104 16316 10160
rect 16252 10100 16316 10104
rect 5948 9888 6012 9892
rect 5948 9832 5998 9888
rect 5998 9832 6012 9888
rect 5948 9828 6012 9832
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 8524 9692 8588 9756
rect 796 9556 860 9620
rect 13124 9420 13188 9484
rect 14228 9556 14292 9620
rect 13676 9284 13740 9348
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 1900 9148 1964 9212
rect 7236 9148 7300 9212
rect 2268 9012 2332 9076
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 14228 8604 14292 8668
rect 17908 8604 17972 8668
rect 6500 8332 6564 8396
rect 13124 8332 13188 8396
rect 2636 8196 2700 8260
rect 14412 8196 14476 8260
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 3924 7924 3988 7988
rect 13676 7788 13740 7852
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 7604 7380 7668 7444
rect 17172 7380 17236 7444
rect 5028 7244 5092 7308
rect 7420 7244 7484 7308
rect 17356 7108 17420 7172
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 17908 6972 17972 7036
rect 15332 6836 15396 6900
rect 17540 6836 17604 6900
rect 1164 6700 1228 6764
rect 9996 6700 10060 6764
rect 15700 6700 15764 6764
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 5764 6428 5828 6492
rect 5948 6292 6012 6356
rect 4108 6216 4172 6220
rect 4108 6160 4158 6216
rect 4158 6160 4172 6216
rect 4108 6156 4172 6160
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7236 5884 7300 5948
rect 5212 5748 5276 5812
rect 5764 5748 5828 5812
rect 22324 5612 22388 5676
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 4844 4796 4908 4860
rect 17172 4524 17236 4588
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 17908 4116 17972 4180
rect 5580 3904 5644 3908
rect 5580 3848 5630 3904
rect 5630 3848 5644 3904
rect 5580 3844 5644 3848
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 5764 3496 5828 3500
rect 5764 3440 5778 3496
rect 5778 3440 5828 3496
rect 5764 3436 5828 3440
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 980 2484 1044 2548
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
rect 60 1940 124 2004
rect 4425 1660 4489 1664
rect 4425 1604 4429 1660
rect 4429 1604 4485 1660
rect 4485 1604 4489 1660
rect 4425 1600 4489 1604
rect 4505 1660 4569 1664
rect 4505 1604 4509 1660
rect 4509 1604 4565 1660
rect 4565 1604 4569 1660
rect 4505 1600 4569 1604
rect 4585 1660 4649 1664
rect 4585 1604 4589 1660
rect 4589 1604 4645 1660
rect 4645 1604 4649 1660
rect 4585 1600 4649 1604
rect 4665 1660 4729 1664
rect 4665 1604 4669 1660
rect 4669 1604 4725 1660
rect 4725 1604 4729 1660
rect 4665 1600 4729 1604
rect 11371 1660 11435 1664
rect 11371 1604 11375 1660
rect 11375 1604 11431 1660
rect 11431 1604 11435 1660
rect 11371 1600 11435 1604
rect 11451 1660 11515 1664
rect 11451 1604 11455 1660
rect 11455 1604 11511 1660
rect 11511 1604 11515 1660
rect 11451 1600 11515 1604
rect 11531 1660 11595 1664
rect 11531 1604 11535 1660
rect 11535 1604 11591 1660
rect 11591 1604 11595 1660
rect 11531 1600 11595 1604
rect 11611 1660 11675 1664
rect 11611 1604 11615 1660
rect 11615 1604 11671 1660
rect 11671 1604 11675 1660
rect 11611 1600 11675 1604
rect 18317 1660 18381 1664
rect 18317 1604 18321 1660
rect 18321 1604 18377 1660
rect 18377 1604 18381 1660
rect 18317 1600 18381 1604
rect 18397 1660 18461 1664
rect 18397 1604 18401 1660
rect 18401 1604 18457 1660
rect 18457 1604 18461 1660
rect 18397 1600 18461 1604
rect 18477 1660 18541 1664
rect 18477 1604 18481 1660
rect 18481 1604 18537 1660
rect 18537 1604 18541 1660
rect 18477 1600 18541 1604
rect 18557 1660 18621 1664
rect 18557 1604 18561 1660
rect 18561 1604 18617 1660
rect 18617 1604 18621 1660
rect 18557 1600 18621 1604
rect 25263 1660 25327 1664
rect 25263 1604 25267 1660
rect 25267 1604 25323 1660
rect 25323 1604 25327 1660
rect 25263 1600 25327 1604
rect 25343 1660 25407 1664
rect 25343 1604 25347 1660
rect 25347 1604 25403 1660
rect 25403 1604 25407 1660
rect 25343 1600 25407 1604
rect 25423 1660 25487 1664
rect 25423 1604 25427 1660
rect 25427 1604 25483 1660
rect 25483 1604 25487 1660
rect 25423 1600 25487 1604
rect 25503 1660 25567 1664
rect 25503 1604 25507 1660
rect 25507 1604 25563 1660
rect 25563 1604 25567 1660
rect 25503 1600 25567 1604
rect 13492 1260 13556 1324
rect 7898 1116 7962 1120
rect 7898 1060 7902 1116
rect 7902 1060 7958 1116
rect 7958 1060 7962 1116
rect 7898 1056 7962 1060
rect 7978 1116 8042 1120
rect 7978 1060 7982 1116
rect 7982 1060 8038 1116
rect 8038 1060 8042 1116
rect 7978 1056 8042 1060
rect 8058 1116 8122 1120
rect 8058 1060 8062 1116
rect 8062 1060 8118 1116
rect 8118 1060 8122 1116
rect 8058 1056 8122 1060
rect 8138 1116 8202 1120
rect 8138 1060 8142 1116
rect 8142 1060 8198 1116
rect 8198 1060 8202 1116
rect 8138 1056 8202 1060
rect 14844 1116 14908 1120
rect 14844 1060 14848 1116
rect 14848 1060 14904 1116
rect 14904 1060 14908 1116
rect 14844 1056 14908 1060
rect 14924 1116 14988 1120
rect 14924 1060 14928 1116
rect 14928 1060 14984 1116
rect 14984 1060 14988 1116
rect 14924 1056 14988 1060
rect 15004 1116 15068 1120
rect 15004 1060 15008 1116
rect 15008 1060 15064 1116
rect 15064 1060 15068 1116
rect 15004 1056 15068 1060
rect 15084 1116 15148 1120
rect 15084 1060 15088 1116
rect 15088 1060 15144 1116
rect 15144 1060 15148 1116
rect 15084 1056 15148 1060
rect 21790 1116 21854 1120
rect 21790 1060 21794 1116
rect 21794 1060 21850 1116
rect 21850 1060 21854 1116
rect 21790 1056 21854 1060
rect 21870 1116 21934 1120
rect 21870 1060 21874 1116
rect 21874 1060 21930 1116
rect 21930 1060 21934 1116
rect 21870 1056 21934 1060
rect 21950 1116 22014 1120
rect 21950 1060 21954 1116
rect 21954 1060 22010 1116
rect 22010 1060 22014 1116
rect 21950 1056 22014 1060
rect 22030 1116 22094 1120
rect 22030 1060 22034 1116
rect 22034 1060 22090 1116
rect 22090 1060 22094 1116
rect 22030 1056 22094 1060
rect 28736 1116 28800 1120
rect 28736 1060 28740 1116
rect 28740 1060 28796 1116
rect 28796 1060 28800 1116
rect 28736 1056 28800 1060
rect 28816 1116 28880 1120
rect 28816 1060 28820 1116
rect 28820 1060 28876 1116
rect 28876 1060 28880 1116
rect 28816 1056 28880 1060
rect 28896 1116 28960 1120
rect 28896 1060 28900 1116
rect 28900 1060 28956 1116
rect 28956 1060 28960 1116
rect 28896 1056 28960 1060
rect 28976 1116 29040 1120
rect 28976 1060 28980 1116
rect 28980 1060 29036 1116
rect 29036 1060 29040 1116
rect 28976 1056 29040 1060
<< metal4 >>
rect 4417 32128 4737 32688
rect 4417 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4737 32128
rect 4417 31040 4737 32064
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 7890 32672 8210 32688
rect 7890 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8210 32672
rect 7890 31584 8210 32608
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 11363 32128 11683 32688
rect 11363 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11683 32128
rect 11363 31040 11683 32064
rect 14836 32672 15156 32688
rect 14836 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15156 32672
rect 14595 31788 14661 31789
rect 14595 31724 14596 31788
rect 14660 31724 14661 31788
rect 14595 31723 14661 31724
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 10547 30020 10613 30021
rect 10547 29956 10548 30020
rect 10612 29956 10613 30020
rect 10547 29955 10613 29956
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 5211 28524 5277 28525
rect 5211 28460 5212 28524
rect 5276 28460 5277 28524
rect 5211 28459 5277 28460
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4107 26076 4173 26077
rect 4107 26012 4108 26076
rect 4172 26012 4173 26076
rect 4107 26011 4173 26012
rect 3187 25396 3253 25397
rect 3187 25332 3188 25396
rect 3252 25332 3253 25396
rect 3187 25331 3253 25332
rect 3190 21589 3250 25331
rect 3187 21588 3253 21589
rect 3187 21524 3188 21588
rect 3252 21524 3253 21588
rect 3187 21523 3253 21524
rect 1163 20364 1229 20365
rect 1163 20300 1164 20364
rect 1228 20300 1229 20364
rect 1163 20299 1229 20300
rect 795 19684 861 19685
rect 795 19620 796 19684
rect 860 19620 861 19684
rect 795 19619 861 19620
rect 59 12476 125 12477
rect 59 12412 60 12476
rect 124 12412 125 12476
rect 59 12411 125 12412
rect 62 2005 122 12411
rect 798 9621 858 19619
rect 979 14380 1045 14381
rect 979 14316 980 14380
rect 1044 14316 1045 14380
rect 979 14315 1045 14316
rect 795 9620 861 9621
rect 795 9556 796 9620
rect 860 9556 861 9620
rect 795 9555 861 9556
rect 982 2549 1042 14315
rect 1166 6765 1226 20299
rect 4110 20229 4170 26011
rect 4417 25600 4737 26624
rect 5214 26621 5274 28459
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 5579 27844 5645 27845
rect 5579 27780 5580 27844
rect 5644 27780 5645 27844
rect 5579 27779 5645 27780
rect 5211 26620 5277 26621
rect 5211 26556 5212 26620
rect 5276 26556 5277 26620
rect 5211 26555 5277 26556
rect 5214 26349 5274 26555
rect 5211 26348 5277 26349
rect 5211 26284 5212 26348
rect 5276 26284 5277 26348
rect 5211 26283 5277 26284
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4291 23628 4357 23629
rect 4291 23564 4292 23628
rect 4356 23564 4357 23628
rect 4291 23563 4357 23564
rect 4107 20228 4173 20229
rect 4107 20164 4108 20228
rect 4172 20164 4173 20228
rect 4107 20163 4173 20164
rect 4294 18325 4354 23563
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 5214 21181 5274 26283
rect 5395 24988 5461 24989
rect 5395 24924 5396 24988
rect 5460 24924 5461 24988
rect 5395 24923 5461 24924
rect 5211 21180 5277 21181
rect 5211 21116 5212 21180
rect 5276 21116 5277 21180
rect 5211 21115 5277 21116
rect 5211 21044 5277 21045
rect 5211 20980 5212 21044
rect 5276 20980 5277 21044
rect 5211 20979 5277 20980
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4291 18324 4357 18325
rect 4291 18260 4292 18324
rect 4356 18260 4357 18324
rect 4291 18259 4357 18260
rect 1899 18052 1965 18053
rect 1899 17988 1900 18052
rect 1964 17988 1965 18052
rect 1899 17987 1965 17988
rect 1902 9213 1962 17987
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 2267 17236 2333 17237
rect 2267 17172 2268 17236
rect 2332 17172 2333 17236
rect 2267 17171 2333 17172
rect 2270 12069 2330 17171
rect 4417 16896 4737 17920
rect 5214 17917 5274 20979
rect 5398 19957 5458 24923
rect 5582 22677 5642 27779
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 6683 26484 6749 26485
rect 6683 26420 6684 26484
rect 6748 26420 6749 26484
rect 6683 26419 6749 26420
rect 6315 24036 6381 24037
rect 6315 23972 6316 24036
rect 6380 23972 6381 24036
rect 6315 23971 6381 23972
rect 5579 22676 5645 22677
rect 5579 22612 5580 22676
rect 5644 22612 5645 22676
rect 5579 22611 5645 22612
rect 6318 21861 6378 23971
rect 6686 23085 6746 26419
rect 7890 26144 8210 27168
rect 9259 26348 9325 26349
rect 9259 26284 9260 26348
rect 9324 26284 9325 26348
rect 9259 26283 9325 26284
rect 8339 26212 8405 26213
rect 8339 26148 8340 26212
rect 8404 26148 8405 26212
rect 8339 26147 8405 26148
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7603 25668 7669 25669
rect 7603 25604 7604 25668
rect 7668 25604 7669 25668
rect 7603 25603 7669 25604
rect 7051 23900 7117 23901
rect 7051 23836 7052 23900
rect 7116 23836 7117 23900
rect 7051 23835 7117 23836
rect 6683 23084 6749 23085
rect 6683 23020 6684 23084
rect 6748 23020 6749 23084
rect 6683 23019 6749 23020
rect 6315 21860 6381 21861
rect 6315 21796 6316 21860
rect 6380 21796 6381 21860
rect 6315 21795 6381 21796
rect 6686 21045 6746 23019
rect 6683 21044 6749 21045
rect 6683 20980 6684 21044
rect 6748 20980 6749 21044
rect 6683 20979 6749 20980
rect 5395 19956 5461 19957
rect 5395 19892 5396 19956
rect 5460 19892 5461 19956
rect 5395 19891 5461 19892
rect 5395 19548 5461 19549
rect 5395 19484 5396 19548
rect 5460 19484 5461 19548
rect 5395 19483 5461 19484
rect 6499 19548 6565 19549
rect 6499 19484 6500 19548
rect 6564 19484 6565 19548
rect 6499 19483 6565 19484
rect 5027 17916 5093 17917
rect 5027 17852 5028 17916
rect 5092 17852 5093 17916
rect 5027 17851 5093 17852
rect 5211 17916 5277 17917
rect 5211 17852 5212 17916
rect 5276 17852 5277 17916
rect 5211 17851 5277 17852
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 3739 16692 3805 16693
rect 3739 16628 3740 16692
rect 3804 16628 3805 16692
rect 3739 16627 3805 16628
rect 4291 16692 4357 16693
rect 4291 16628 4292 16692
rect 4356 16628 4357 16692
rect 4291 16627 4357 16628
rect 2635 15332 2701 15333
rect 2635 15268 2636 15332
rect 2700 15268 2701 15332
rect 2635 15267 2701 15268
rect 2267 12068 2333 12069
rect 2267 12004 2268 12068
rect 2332 12004 2333 12068
rect 2267 12003 2333 12004
rect 2267 11116 2333 11117
rect 2267 11052 2268 11116
rect 2332 11052 2333 11116
rect 2267 11051 2333 11052
rect 1899 9212 1965 9213
rect 1899 9148 1900 9212
rect 1964 9148 1965 9212
rect 1899 9147 1965 9148
rect 2270 9077 2330 11051
rect 2267 9076 2333 9077
rect 2267 9012 2268 9076
rect 2332 9012 2333 9076
rect 2267 9011 2333 9012
rect 2638 8261 2698 15267
rect 3742 10301 3802 16627
rect 4294 12885 4354 16627
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4291 12884 4357 12885
rect 4291 12820 4292 12884
rect 4356 12820 4357 12884
rect 4291 12819 4357 12820
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 3923 12204 3989 12205
rect 3923 12140 3924 12204
rect 3988 12140 3989 12204
rect 3923 12139 3989 12140
rect 3739 10300 3805 10301
rect 3739 10236 3740 10300
rect 3804 10236 3805 10300
rect 3739 10235 3805 10236
rect 2635 8260 2701 8261
rect 2635 8196 2636 8260
rect 2700 8196 2701 8260
rect 2635 8195 2701 8196
rect 3926 7989 3986 12139
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4107 11116 4173 11117
rect 4107 11052 4108 11116
rect 4172 11052 4173 11116
rect 4107 11051 4173 11052
rect 3923 7988 3989 7989
rect 3923 7924 3924 7988
rect 3988 7924 3989 7988
rect 3923 7923 3989 7924
rect 1163 6764 1229 6765
rect 1163 6700 1164 6764
rect 1228 6700 1229 6764
rect 1163 6699 1229 6700
rect 4110 6221 4170 11051
rect 4417 10368 4737 11392
rect 4843 11116 4909 11117
rect 4843 11052 4844 11116
rect 4908 11052 4909 11116
rect 4843 11051 4909 11052
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4107 6220 4173 6221
rect 4107 6156 4108 6220
rect 4172 6156 4173 6220
rect 4107 6155 4173 6156
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4846 4861 4906 11051
rect 5030 10029 5090 17851
rect 5211 12884 5277 12885
rect 5211 12820 5212 12884
rect 5276 12820 5277 12884
rect 5211 12819 5277 12820
rect 5027 10028 5093 10029
rect 5027 9964 5028 10028
rect 5092 9964 5093 10028
rect 5027 9963 5093 9964
rect 5030 7309 5090 9963
rect 5027 7308 5093 7309
rect 5027 7244 5028 7308
rect 5092 7244 5093 7308
rect 5027 7243 5093 7244
rect 5214 5813 5274 12819
rect 5398 12477 5458 19483
rect 6502 16149 6562 19483
rect 6686 16557 6746 20979
rect 7054 20229 7114 23835
rect 7606 22541 7666 25603
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 8342 23629 8402 26147
rect 8339 23628 8405 23629
rect 8339 23564 8340 23628
rect 8404 23564 8405 23628
rect 8339 23563 8405 23564
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7603 22540 7669 22541
rect 7603 22476 7604 22540
rect 7668 22476 7669 22540
rect 7603 22475 7669 22476
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 8523 20772 8589 20773
rect 8523 20708 8524 20772
rect 8588 20708 8589 20772
rect 8523 20707 8589 20708
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7051 20228 7117 20229
rect 7051 20164 7052 20228
rect 7116 20226 7117 20228
rect 7116 20166 7298 20226
rect 7116 20164 7117 20166
rect 7051 20163 7117 20164
rect 6683 16556 6749 16557
rect 6683 16492 6684 16556
rect 6748 16492 6749 16556
rect 6683 16491 6749 16492
rect 6499 16148 6565 16149
rect 6499 16084 6500 16148
rect 6564 16084 6565 16148
rect 6499 16083 6565 16084
rect 5395 12476 5461 12477
rect 5395 12412 5396 12476
rect 5460 12412 5461 12476
rect 5395 12411 5461 12412
rect 5579 11932 5645 11933
rect 5579 11868 5580 11932
rect 5644 11868 5645 11932
rect 5579 11867 5645 11868
rect 5211 5812 5277 5813
rect 5211 5748 5212 5812
rect 5276 5748 5277 5812
rect 5211 5747 5277 5748
rect 4843 4860 4909 4861
rect 4843 4796 4844 4860
rect 4908 4796 4909 4860
rect 4843 4795 4909 4796
rect 5582 3909 5642 11867
rect 5763 11524 5829 11525
rect 5763 11460 5764 11524
rect 5828 11460 5829 11524
rect 5763 11459 5829 11460
rect 5766 6493 5826 11459
rect 5947 9892 6013 9893
rect 5947 9828 5948 9892
rect 6012 9828 6013 9892
rect 5947 9827 6013 9828
rect 5763 6492 5829 6493
rect 5763 6428 5764 6492
rect 5828 6428 5829 6492
rect 5763 6427 5829 6428
rect 5766 5813 5826 6427
rect 5950 6357 6010 9827
rect 6502 8397 6562 16083
rect 7051 15468 7117 15469
rect 7051 15404 7052 15468
rect 7116 15404 7117 15468
rect 7051 15403 7117 15404
rect 7054 10709 7114 15403
rect 7238 15197 7298 20166
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7603 18188 7669 18189
rect 7603 18124 7604 18188
rect 7668 18124 7669 18188
rect 7603 18123 7669 18124
rect 7419 16284 7485 16285
rect 7419 16220 7420 16284
rect 7484 16220 7485 16284
rect 7419 16219 7485 16220
rect 7235 15196 7301 15197
rect 7235 15132 7236 15196
rect 7300 15132 7301 15196
rect 7235 15131 7301 15132
rect 7051 10708 7117 10709
rect 7051 10644 7052 10708
rect 7116 10644 7117 10708
rect 7051 10643 7117 10644
rect 7235 9212 7301 9213
rect 7235 9148 7236 9212
rect 7300 9148 7301 9212
rect 7235 9147 7301 9148
rect 6499 8396 6565 8397
rect 6499 8332 6500 8396
rect 6564 8332 6565 8396
rect 6499 8331 6565 8332
rect 5947 6356 6013 6357
rect 5947 6292 5948 6356
rect 6012 6292 6013 6356
rect 5947 6291 6013 6292
rect 7238 5949 7298 9147
rect 7422 7309 7482 16219
rect 7606 12749 7666 18123
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7603 12748 7669 12749
rect 7603 12684 7604 12748
rect 7668 12684 7669 12748
rect 7603 12683 7669 12684
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7603 10436 7669 10437
rect 7603 10372 7604 10436
rect 7668 10372 7669 10436
rect 7603 10371 7669 10372
rect 7606 7445 7666 10371
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 8526 9757 8586 20707
rect 9262 20501 9322 26283
rect 10363 26212 10429 26213
rect 10363 26148 10364 26212
rect 10428 26148 10429 26212
rect 10363 26147 10429 26148
rect 9811 25804 9877 25805
rect 9811 25740 9812 25804
rect 9876 25740 9877 25804
rect 9811 25739 9877 25740
rect 9443 23628 9509 23629
rect 9443 23564 9444 23628
rect 9508 23564 9509 23628
rect 9443 23563 9509 23564
rect 9259 20500 9325 20501
rect 9259 20436 9260 20500
rect 9324 20436 9325 20500
rect 9259 20435 9325 20436
rect 9446 13837 9506 23563
rect 9814 16149 9874 25739
rect 10366 24037 10426 26147
rect 10363 24036 10429 24037
rect 10363 23972 10364 24036
rect 10428 23972 10429 24036
rect 10363 23971 10429 23972
rect 10550 23221 10610 29955
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 14411 27708 14477 27709
rect 14411 27644 14412 27708
rect 14476 27644 14477 27708
rect 14411 27643 14477 27644
rect 13307 26756 13373 26757
rect 13307 26692 13308 26756
rect 13372 26692 13373 26756
rect 13307 26691 13373 26692
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 13123 24988 13189 24989
rect 13123 24924 13124 24988
rect 13188 24924 13189 24988
rect 13123 24923 13189 24924
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 13126 24037 13186 24923
rect 13123 24036 13189 24037
rect 13123 23972 13124 24036
rect 13188 23972 13189 24036
rect 13123 23971 13189 23972
rect 12019 23900 12085 23901
rect 12019 23836 12020 23900
rect 12084 23836 12085 23900
rect 12019 23835 12085 23836
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 10547 23220 10613 23221
rect 10547 23156 10548 23220
rect 10612 23156 10613 23220
rect 10547 23155 10613 23156
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 12022 20773 12082 23835
rect 12019 20772 12085 20773
rect 12019 20708 12020 20772
rect 12084 20708 12085 20772
rect 12019 20707 12085 20708
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11835 18052 11901 18053
rect 11835 17988 11836 18052
rect 11900 17988 11901 18052
rect 11835 17987 11901 17988
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 9995 17780 10061 17781
rect 9995 17716 9996 17780
rect 10060 17716 10061 17780
rect 9995 17715 10061 17716
rect 9811 16148 9877 16149
rect 9811 16084 9812 16148
rect 9876 16084 9877 16148
rect 9811 16083 9877 16084
rect 9443 13836 9509 13837
rect 9443 13772 9444 13836
rect 9508 13772 9509 13836
rect 9443 13771 9509 13772
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 9262 11253 9322 13499
rect 9259 11252 9325 11253
rect 9259 11188 9260 11252
rect 9324 11188 9325 11252
rect 9259 11187 9325 11188
rect 8523 9756 8589 9757
rect 8523 9692 8524 9756
rect 8588 9692 8589 9756
rect 8523 9691 8589 9692
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7603 7444 7669 7445
rect 7603 7380 7604 7444
rect 7668 7380 7669 7444
rect 7603 7379 7669 7380
rect 7419 7308 7485 7309
rect 7419 7244 7420 7308
rect 7484 7244 7485 7308
rect 7419 7243 7485 7244
rect 7890 6560 8210 7584
rect 9998 6765 10058 17715
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11838 16149 11898 17987
rect 11835 16148 11901 16149
rect 11835 16084 11836 16148
rect 11900 16084 11901 16148
rect 11835 16083 11901 16084
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11099 13972 11165 13973
rect 11099 13908 11100 13972
rect 11164 13908 11165 13972
rect 11099 13907 11165 13908
rect 10179 12748 10245 12749
rect 10179 12684 10180 12748
rect 10244 12684 10245 12748
rect 10179 12683 10245 12684
rect 10182 10709 10242 12683
rect 10363 12068 10429 12069
rect 10363 12004 10364 12068
rect 10428 12004 10429 12068
rect 10363 12003 10429 12004
rect 10179 10708 10245 10709
rect 10179 10644 10180 10708
rect 10244 10644 10245 10708
rect 10179 10643 10245 10644
rect 10366 10301 10426 12003
rect 10363 10300 10429 10301
rect 10363 10236 10364 10300
rect 10428 10236 10429 10300
rect 10363 10235 10429 10236
rect 11102 10029 11162 13907
rect 11363 13632 11683 14656
rect 12022 13701 12082 20707
rect 12203 19548 12269 19549
rect 12203 19484 12204 19548
rect 12268 19484 12269 19548
rect 12203 19483 12269 19484
rect 12206 17509 12266 19483
rect 13126 17917 13186 23971
rect 13310 19277 13370 26691
rect 14043 26620 14109 26621
rect 14043 26556 14044 26620
rect 14108 26556 14109 26620
rect 14043 26555 14109 26556
rect 13675 20092 13741 20093
rect 13675 20028 13676 20092
rect 13740 20028 13741 20092
rect 13675 20027 13741 20028
rect 13491 19412 13557 19413
rect 13491 19348 13492 19412
rect 13556 19348 13557 19412
rect 13491 19347 13557 19348
rect 13307 19276 13373 19277
rect 13307 19212 13308 19276
rect 13372 19212 13373 19276
rect 13307 19211 13373 19212
rect 13123 17916 13189 17917
rect 13123 17852 13124 17916
rect 13188 17852 13189 17916
rect 13123 17851 13189 17852
rect 12203 17508 12269 17509
rect 12203 17444 12204 17508
rect 12268 17444 12269 17508
rect 12203 17443 12269 17444
rect 13123 17236 13189 17237
rect 13123 17172 13124 17236
rect 13188 17172 13189 17236
rect 13123 17171 13189 17172
rect 12019 13700 12085 13701
rect 12019 13636 12020 13700
rect 12084 13636 12085 13700
rect 12019 13635 12085 13636
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11099 10028 11165 10029
rect 11099 9964 11100 10028
rect 11164 9964 11165 10028
rect 11099 9963 11165 9964
rect 11363 9280 11683 10304
rect 13126 9485 13186 17171
rect 13494 16013 13554 19347
rect 13491 16012 13557 16013
rect 13491 15948 13492 16012
rect 13556 15948 13557 16012
rect 13491 15947 13557 15948
rect 13678 15333 13738 20027
rect 14046 17917 14106 26555
rect 14227 19956 14293 19957
rect 14227 19892 14228 19956
rect 14292 19892 14293 19956
rect 14227 19891 14293 19892
rect 14043 17916 14109 17917
rect 14043 17852 14044 17916
rect 14108 17852 14109 17916
rect 14043 17851 14109 17852
rect 13675 15332 13741 15333
rect 13675 15268 13676 15332
rect 13740 15268 13741 15332
rect 13675 15267 13741 15268
rect 14230 13973 14290 19891
rect 14414 19413 14474 27643
rect 14598 25533 14658 31723
rect 14836 31584 15156 32608
rect 18309 32128 18629 32688
rect 18309 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18629 32128
rect 15883 31652 15949 31653
rect 15883 31588 15884 31652
rect 15948 31588 15949 31652
rect 15883 31587 15949 31588
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14595 25532 14661 25533
rect 14595 25468 14596 25532
rect 14660 25468 14661 25532
rect 14595 25467 14661 25468
rect 14836 25056 15156 26080
rect 15331 25124 15397 25125
rect 15331 25060 15332 25124
rect 15396 25060 15397 25124
rect 15331 25059 15397 25060
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14595 22268 14661 22269
rect 14595 22204 14596 22268
rect 14660 22204 14661 22268
rect 14595 22203 14661 22204
rect 14598 19957 14658 22203
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 15334 21453 15394 25059
rect 15886 24717 15946 31587
rect 18309 31040 18629 32064
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 17171 30836 17237 30837
rect 17171 30772 17172 30836
rect 17236 30772 17237 30836
rect 17171 30771 17237 30772
rect 17174 28117 17234 30771
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 17907 28660 17973 28661
rect 17907 28596 17908 28660
rect 17972 28596 17973 28660
rect 17907 28595 17973 28596
rect 17355 28252 17421 28253
rect 17355 28188 17356 28252
rect 17420 28188 17421 28252
rect 17355 28187 17421 28188
rect 17171 28116 17237 28117
rect 17171 28052 17172 28116
rect 17236 28052 17237 28116
rect 17171 28051 17237 28052
rect 16067 24988 16133 24989
rect 16067 24924 16068 24988
rect 16132 24924 16133 24988
rect 16067 24923 16133 24924
rect 15883 24716 15949 24717
rect 15883 24652 15884 24716
rect 15948 24652 15949 24716
rect 15883 24651 15949 24652
rect 16070 21997 16130 24923
rect 16435 22948 16501 22949
rect 16435 22884 16436 22948
rect 16500 22884 16501 22948
rect 16435 22883 16501 22884
rect 16067 21996 16133 21997
rect 16067 21932 16068 21996
rect 16132 21932 16133 21996
rect 16067 21931 16133 21932
rect 15331 21452 15397 21453
rect 15331 21388 15332 21452
rect 15396 21388 15397 21452
rect 15331 21387 15397 21388
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14595 19956 14661 19957
rect 14595 19892 14596 19956
rect 14660 19892 14661 19956
rect 14595 19891 14661 19892
rect 14595 19820 14661 19821
rect 14595 19756 14596 19820
rect 14660 19756 14661 19820
rect 14595 19755 14661 19756
rect 14411 19412 14477 19413
rect 14411 19348 14412 19412
rect 14476 19348 14477 19412
rect 14411 19347 14477 19348
rect 14411 18052 14477 18053
rect 14411 17988 14412 18052
rect 14476 17988 14477 18052
rect 14411 17987 14477 17988
rect 14414 14789 14474 17987
rect 14411 14788 14477 14789
rect 14411 14724 14412 14788
rect 14476 14724 14477 14788
rect 14411 14723 14477 14724
rect 14227 13972 14293 13973
rect 14227 13908 14228 13972
rect 14292 13908 14293 13972
rect 14227 13907 14293 13908
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 13123 9484 13189 9485
rect 13123 9420 13124 9484
rect 13188 9420 13189 9484
rect 13123 9419 13189 9420
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 13126 8397 13186 9419
rect 13123 8396 13189 8397
rect 13123 8332 13124 8396
rect 13188 8332 13189 8396
rect 13123 8331 13189 8332
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 9995 6764 10061 6765
rect 9995 6700 9996 6764
rect 10060 6700 10061 6764
rect 9995 6699 10061 6700
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7235 5948 7301 5949
rect 7235 5884 7236 5948
rect 7300 5884 7301 5948
rect 7235 5883 7301 5884
rect 5763 5812 5829 5813
rect 5763 5748 5764 5812
rect 5828 5748 5829 5812
rect 5763 5747 5829 5748
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 5766 3501 5826 5747
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 5763 3500 5829 3501
rect 5763 3436 5764 3500
rect 5828 3436 5829 3500
rect 5763 3435 5829 3436
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 979 2548 1045 2549
rect 979 2484 980 2548
rect 1044 2484 1045 2548
rect 979 2483 1045 2484
rect 59 2004 125 2005
rect 59 1940 60 2004
rect 124 1940 125 2004
rect 59 1939 125 1940
rect 4417 1664 4737 2688
rect 4417 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4737 1664
rect 4417 1040 4737 1600
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 1120 8210 2144
rect 7890 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8210 1120
rect 7890 1040 8210 1056
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 1664 11683 2688
rect 11363 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11683 1664
rect 11363 1040 11683 1600
rect 13494 1325 13554 13771
rect 14411 13428 14477 13429
rect 14411 13364 14412 13428
rect 14476 13364 14477 13428
rect 14411 13363 14477 13364
rect 14227 9620 14293 9621
rect 14227 9556 14228 9620
rect 14292 9556 14293 9620
rect 14227 9555 14293 9556
rect 13675 9348 13741 9349
rect 13675 9284 13676 9348
rect 13740 9284 13741 9348
rect 13675 9283 13741 9284
rect 13678 7853 13738 9283
rect 14230 8669 14290 9555
rect 14227 8668 14293 8669
rect 14227 8604 14228 8668
rect 14292 8604 14293 8668
rect 14227 8603 14293 8604
rect 14414 8261 14474 13363
rect 14598 12885 14658 19755
rect 14836 19616 15156 20640
rect 15515 19956 15581 19957
rect 15515 19892 15516 19956
rect 15580 19892 15581 19956
rect 15515 19891 15581 19892
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 15331 15876 15397 15877
rect 15331 15812 15332 15876
rect 15396 15812 15397 15876
rect 15331 15811 15397 15812
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14595 12884 14661 12885
rect 14595 12820 14596 12884
rect 14660 12820 14661 12884
rect 14595 12819 14661 12820
rect 14836 12000 15156 13024
rect 15334 12341 15394 15811
rect 15518 13565 15578 19891
rect 16070 19005 16130 21931
rect 16067 19004 16133 19005
rect 16067 18940 16068 19004
rect 16132 18940 16133 19004
rect 16067 18939 16133 18940
rect 15883 18732 15949 18733
rect 15883 18668 15884 18732
rect 15948 18668 15949 18732
rect 15883 18667 15949 18668
rect 15515 13564 15581 13565
rect 15515 13500 15516 13564
rect 15580 13500 15581 13564
rect 15515 13499 15581 13500
rect 15331 12340 15397 12341
rect 15331 12276 15332 12340
rect 15396 12276 15397 12340
rect 15331 12275 15397 12276
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 15886 11253 15946 18667
rect 16438 17917 16498 22883
rect 17358 22677 17418 28187
rect 17910 26077 17970 28595
rect 18309 27776 18629 28800
rect 21782 32672 22102 32688
rect 21782 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22102 32672
rect 21782 31584 22102 32608
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 19379 27844 19445 27845
rect 19379 27780 19380 27844
rect 19444 27780 19445 27844
rect 19379 27779 19445 27780
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 17907 26076 17973 26077
rect 17907 26012 17908 26076
rect 17972 26012 17973 26076
rect 17907 26011 17973 26012
rect 18309 25600 18629 26624
rect 19382 25941 19442 27779
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 25255 32128 25575 32688
rect 25255 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25575 32128
rect 25255 31040 25575 32064
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 22323 26212 22389 26213
rect 22323 26148 22324 26212
rect 22388 26148 22389 26212
rect 22323 26147 22389 26148
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 19379 25940 19445 25941
rect 19379 25876 19380 25940
rect 19444 25876 19445 25940
rect 19379 25875 19445 25876
rect 18827 25668 18893 25669
rect 18827 25604 18828 25668
rect 18892 25604 18893 25668
rect 18827 25603 18893 25604
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18830 24989 18890 25603
rect 21782 25056 22102 26080
rect 22326 25261 22386 26147
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 22323 25260 22389 25261
rect 22323 25196 22324 25260
rect 22388 25196 22389 25260
rect 22323 25195 22389 25196
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 18827 24988 18893 24989
rect 18827 24924 18828 24988
rect 18892 24924 18893 24988
rect 18827 24923 18893 24924
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 19011 24036 19077 24037
rect 19011 23972 19012 24036
rect 19076 23972 19077 24036
rect 19011 23971 19077 23972
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 17355 22676 17421 22677
rect 17355 22612 17356 22676
rect 17420 22612 17421 22676
rect 17355 22611 17421 22612
rect 18091 22676 18157 22677
rect 18091 22612 18092 22676
rect 18156 22612 18157 22676
rect 18091 22611 18157 22612
rect 17907 19684 17973 19685
rect 17907 19620 17908 19684
rect 17972 19620 17973 19684
rect 17907 19619 17973 19620
rect 16619 19412 16685 19413
rect 16619 19348 16620 19412
rect 16684 19348 16685 19412
rect 16619 19347 16685 19348
rect 16251 17916 16317 17917
rect 16251 17852 16252 17916
rect 16316 17852 16317 17916
rect 16251 17851 16317 17852
rect 16435 17916 16501 17917
rect 16435 17852 16436 17916
rect 16500 17852 16501 17916
rect 16435 17851 16501 17852
rect 16067 14924 16133 14925
rect 16067 14860 16068 14924
rect 16132 14860 16133 14924
rect 16067 14859 16133 14860
rect 16070 11797 16130 14859
rect 16067 11796 16133 11797
rect 16067 11732 16068 11796
rect 16132 11732 16133 11796
rect 16067 11731 16133 11732
rect 15331 11252 15397 11253
rect 15331 11188 15332 11252
rect 15396 11188 15397 11252
rect 15331 11187 15397 11188
rect 15883 11252 15949 11253
rect 15883 11188 15884 11252
rect 15948 11188 15949 11252
rect 15883 11187 15949 11188
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14411 8260 14477 8261
rect 14411 8196 14412 8260
rect 14476 8196 14477 8260
rect 14411 8195 14477 8196
rect 13675 7852 13741 7853
rect 13675 7788 13676 7852
rect 13740 7788 13741 7852
rect 13675 7787 13741 7788
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 15334 6901 15394 11187
rect 16070 10845 16130 11731
rect 16067 10844 16133 10845
rect 16067 10780 16068 10844
rect 16132 10780 16133 10844
rect 16067 10779 16133 10780
rect 16254 10165 16314 17851
rect 16622 15469 16682 19347
rect 17910 19141 17970 19619
rect 17907 19140 17973 19141
rect 17907 19076 17908 19140
rect 17972 19076 17973 19140
rect 17907 19075 17973 19076
rect 18094 17781 18154 22611
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 19014 21725 19074 23971
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 19379 22948 19445 22949
rect 19379 22884 19380 22948
rect 19444 22884 19445 22948
rect 19379 22883 19445 22884
rect 19195 22404 19261 22405
rect 19195 22340 19196 22404
rect 19260 22340 19261 22404
rect 19195 22339 19261 22340
rect 19011 21724 19077 21725
rect 19011 21660 19012 21724
rect 19076 21660 19077 21724
rect 19011 21659 19077 21660
rect 18827 21452 18893 21453
rect 18827 21388 18828 21452
rect 18892 21388 18893 21452
rect 18827 21387 18893 21388
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18091 17780 18157 17781
rect 18091 17716 18092 17780
rect 18156 17716 18157 17780
rect 18091 17715 18157 17716
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18830 16421 18890 21387
rect 19198 21045 19258 22339
rect 19195 21044 19261 21045
rect 19195 20980 19196 21044
rect 19260 20980 19261 21044
rect 19195 20979 19261 20980
rect 19382 20637 19442 22883
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 20299 21452 20365 21453
rect 20299 21388 20300 21452
rect 20364 21388 20365 21452
rect 20299 21387 20365 21388
rect 19379 20636 19445 20637
rect 19379 20572 19380 20636
rect 19444 20572 19445 20636
rect 19379 20571 19445 20572
rect 19379 19140 19445 19141
rect 19379 19076 19380 19140
rect 19444 19076 19445 19140
rect 19379 19075 19445 19076
rect 20115 19140 20181 19141
rect 20115 19076 20116 19140
rect 20180 19076 20181 19140
rect 20115 19075 20181 19076
rect 19382 16965 19442 19075
rect 19747 18052 19813 18053
rect 19747 17988 19748 18052
rect 19812 17988 19813 18052
rect 19747 17987 19813 17988
rect 19563 17508 19629 17509
rect 19563 17444 19564 17508
rect 19628 17444 19629 17508
rect 19563 17443 19629 17444
rect 19379 16964 19445 16965
rect 19379 16900 19380 16964
rect 19444 16900 19445 16964
rect 19379 16899 19445 16900
rect 18827 16420 18893 16421
rect 18827 16356 18828 16420
rect 18892 16356 18893 16420
rect 18827 16355 18893 16356
rect 19382 16149 19442 16899
rect 19379 16148 19445 16149
rect 19379 16084 19380 16148
rect 19444 16084 19445 16148
rect 19379 16083 19445 16084
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 16619 15468 16685 15469
rect 16619 15404 16620 15468
rect 16684 15404 16685 15468
rect 16619 15403 16685 15404
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 17355 13156 17421 13157
rect 17355 13092 17356 13156
rect 17420 13092 17421 13156
rect 17355 13091 17421 13092
rect 15699 10164 15765 10165
rect 15699 10100 15700 10164
rect 15764 10100 15765 10164
rect 15699 10099 15765 10100
rect 16251 10164 16317 10165
rect 16251 10100 16252 10164
rect 16316 10100 16317 10164
rect 16251 10099 16317 10100
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 15702 6765 15762 10099
rect 17171 7444 17237 7445
rect 17171 7380 17172 7444
rect 17236 7380 17237 7444
rect 17171 7379 17237 7380
rect 15699 6764 15765 6765
rect 15699 6700 15700 6764
rect 15764 6700 15765 6764
rect 15699 6699 15765 6700
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 17174 4589 17234 7379
rect 17358 7173 17418 13091
rect 17907 12748 17973 12749
rect 17907 12684 17908 12748
rect 17972 12684 17973 12748
rect 17907 12683 17973 12684
rect 17539 12476 17605 12477
rect 17539 12412 17540 12476
rect 17604 12412 17605 12476
rect 17539 12411 17605 12412
rect 17355 7172 17421 7173
rect 17355 7108 17356 7172
rect 17420 7108 17421 7172
rect 17355 7107 17421 7108
rect 17542 6901 17602 12411
rect 17910 8669 17970 12683
rect 18309 12544 18629 13568
rect 19566 13429 19626 17443
rect 19563 13428 19629 13429
rect 19563 13364 19564 13428
rect 19628 13364 19629 13428
rect 19563 13363 19629 13364
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 19750 12341 19810 17987
rect 19931 14516 19997 14517
rect 19931 14452 19932 14516
rect 19996 14452 19997 14516
rect 19931 14451 19997 14452
rect 19747 12340 19813 12341
rect 19747 12276 19748 12340
rect 19812 12276 19813 12340
rect 19747 12275 19813 12276
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 19934 10845 19994 14451
rect 20118 13701 20178 19075
rect 20302 18733 20362 21387
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 20483 20228 20549 20229
rect 20483 20164 20484 20228
rect 20548 20164 20549 20228
rect 20483 20163 20549 20164
rect 20299 18732 20365 18733
rect 20299 18668 20300 18732
rect 20364 18668 20365 18732
rect 20299 18667 20365 18668
rect 20486 15197 20546 20163
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 22323 18868 22389 18869
rect 22323 18804 22324 18868
rect 22388 18804 22389 18868
rect 22323 18803 22389 18804
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 20483 15196 20549 15197
rect 20483 15132 20484 15196
rect 20548 15132 20549 15196
rect 20483 15131 20549 15132
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 20115 13700 20181 13701
rect 20115 13636 20116 13700
rect 20180 13636 20181 13700
rect 20115 13635 20181 13636
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 19931 10844 19997 10845
rect 19931 10780 19932 10844
rect 19996 10780 19997 10844
rect 19931 10779 19997 10780
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 17907 8668 17973 8669
rect 17907 8604 17908 8668
rect 17972 8604 17973 8668
rect 17907 8603 17973 8604
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 17907 7036 17973 7037
rect 17907 6972 17908 7036
rect 17972 6972 17973 7036
rect 17907 6971 17973 6972
rect 17539 6900 17605 6901
rect 17539 6836 17540 6900
rect 17604 6836 17605 6900
rect 17539 6835 17605 6836
rect 17171 4588 17237 4589
rect 17171 4524 17172 4588
rect 17236 4524 17237 4588
rect 17171 4523 17237 4524
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 17910 4181 17970 6971
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 17907 4180 17973 4181
rect 17907 4116 17908 4180
rect 17972 4116 17973 4180
rect 17907 4115 17973 4116
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 13491 1324 13557 1325
rect 13491 1260 13492 1324
rect 13556 1260 13557 1324
rect 13491 1259 13557 1260
rect 14836 1120 15156 2144
rect 14836 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15156 1120
rect 14836 1040 15156 1056
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 1664 18629 2688
rect 18309 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18629 1664
rect 18309 1040 18629 1600
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 22326 5677 22386 18803
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 22323 5676 22389 5677
rect 22323 5612 22324 5676
rect 22388 5612 22389 5676
rect 22323 5611 22389 5612
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 1120 22102 2144
rect 21782 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22102 1120
rect 21782 1040 22102 1056
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 1664 25575 2688
rect 25255 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25575 1664
rect 25255 1040 25575 1600
rect 28728 32672 29048 32688
rect 28728 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29048 32672
rect 28728 31584 29048 32608
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 1120 29048 2144
rect 28728 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29048 1120
rect 28728 1040 29048 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 10304 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 27600 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 2760 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1676037725
transform 1 0 10856 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1676037725
transform 1 0 14996 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1676037725
transform 1 0 15824 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_271
timestamp 1676037725
transform 1 0 26036 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_286
timestamp 1676037725
transform 1 0 27416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_290
timestamp 1676037725
transform 1 0 27784 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1676037725
transform 1 0 28520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1676037725
transform 1 0 5428 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1676037725
transform 1 0 6900 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1676037725
transform 1 0 7544 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1676037725
transform 1 0 9384 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1676037725
transform 1 0 11960 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1676037725
transform 1 0 14720 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1676037725
transform 1 0 15088 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1676037725
transform 1 0 15732 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1676037725
transform 1 0 20792 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1676037725
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_263
timestamp 1676037725
transform 1 0 25300 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1676037725
transform 1 0 25944 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1676037725
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1676037725
transform 1 0 13432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1676037725
transform 1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1676037725
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1676037725
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_227
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1676037725
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1676037725
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_41
timestamp 1676037725
transform 1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1676037725
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_73
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1676037725
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1676037725
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_179
timestamp 1676037725
transform 1 0 17572 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_251
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_269
timestamp 1676037725
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1676037725
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_35
timestamp 1676037725
transform 1 0 4324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1676037725
transform 1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1676037725
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1676037725
transform 1 0 12604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1676037725
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_148
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_156
timestamp 1676037725
transform 1 0 15456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1676037725
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1676037725
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_225
timestamp 1676037725
transform 1 0 21804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1676037725
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1676037725
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1676037725
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1676037725
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1676037725
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_126
timestamp 1676037725
transform 1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1676037725
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 1676037725
transform 1 0 13984 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1676037725
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_176
timestamp 1676037725
transform 1 0 17296 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1676037725
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_202
timestamp 1676037725
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1676037725
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_253
timestamp 1676037725
transform 1 0 24380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_286
timestamp 1676037725
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1676037725
transform 1 0 28520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_37
timestamp 1676037725
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1676037725
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1676037725
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1676037725
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1676037725
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1676037725
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_103
timestamp 1676037725
transform 1 0 10580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1676037725
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_119
timestamp 1676037725
transform 1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1676037725
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_169
timestamp 1676037725
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1676037725
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_202
timestamp 1676037725
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_206
timestamp 1676037725
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_258
timestamp 1676037725
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1676037725
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_291
timestamp 1676037725
transform 1 0 27876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_29
timestamp 1676037725
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1676037725
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_72
timestamp 1676037725
transform 1 0 7728 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1676037725
transform 1 0 8280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_85
timestamp 1676037725
transform 1 0 8924 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1676037725
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1676037725
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1676037725
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1676037725
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_190
timestamp 1676037725
transform 1 0 18584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1676037725
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_208
timestamp 1676037725
transform 1 0 20240 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1676037725
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1676037725
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_257
timestamp 1676037725
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_286
timestamp 1676037725
transform 1 0 27416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1676037725
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1676037725
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_35
timestamp 1676037725
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1676037725
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_54
timestamp 1676037725
transform 1 0 6072 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1676037725
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_70
timestamp 1676037725
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1676037725
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1676037725
transform 1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1676037725
transform 1 0 11592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_120
timestamp 1676037725
transform 1 0 12144 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1676037725
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1676037725
transform 1 0 15456 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_168
timestamp 1676037725
transform 1 0 16560 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_180
timestamp 1676037725
transform 1 0 17664 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1676037725
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_240
timestamp 1676037725
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_279
timestamp 1676037725
transform 1 0 26772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1676037725
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1676037725
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1676037725
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1676037725
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1676037725
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1676037725
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1676037725
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1676037725
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1676037725
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1676037725
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1676037725
transform 1 0 14628 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_196
timestamp 1676037725
transform 1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1676037725
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1676037725
transform 1 0 23644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_252
timestamp 1676037725
transform 1 0 24288 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1676037725
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_63
timestamp 1676037725
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_75
timestamp 1676037725
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_98
timestamp 1676037725
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_110
timestamp 1676037725
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1676037725
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1676037725
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_173
timestamp 1676037725
transform 1 0 17020 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1676037725
transform 1 0 17664 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1676037725
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_240
timestamp 1676037725
transform 1 0 23184 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1676037725
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1676037725
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_291
timestamp 1676037725
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1676037725
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_44
timestamp 1676037725
transform 1 0 5152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1676037725
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1676037725
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_83
timestamp 1676037725
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1676037725
transform 1 0 11960 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1676037725
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1676037725
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 1676037725
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1676037725
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_214
timestamp 1676037725
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_231
timestamp 1676037725
transform 1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_238
timestamp 1676037725
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1676037725
transform 1 0 23644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1676037725
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1676037725
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_42
timestamp 1676037725
transform 1 0 4968 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1676037725
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1676037725
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_68
timestamp 1676037725
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_104
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_111
timestamp 1676037725
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1676037725
transform 1 0 12880 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_148
timestamp 1676037725
transform 1 0 14720 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_156
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_167
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1676037725
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_182
timestamp 1676037725
transform 1 0 17848 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_188
timestamp 1676037725
transform 1 0 18400 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_204
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_210
timestamp 1676037725
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_227
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_237
timestamp 1676037725
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1676037725
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_266
timestamp 1676037725
transform 1 0 25576 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_284
timestamp 1676037725
transform 1 0 27232 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1676037725
transform 1 0 28336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_29
timestamp 1676037725
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_45
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1676037725
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_67
timestamp 1676037725
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1676037725
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_88
timestamp 1676037725
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1676037725
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1676037725
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1676037725
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_238
timestamp 1676037725
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_255
timestamp 1676037725
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 1676037725
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1676037725
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_52
timestamp 1676037725
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1676037725
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1676037725
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_116
timestamp 1676037725
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1676037725
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1676037725
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1676037725
transform 1 0 19872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_220
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_227
timestamp 1676037725
transform 1 0 21988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_271
timestamp 1676037725
transform 1 0 26036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_294
timestamp 1676037725
transform 1 0 28152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1676037725
transform 1 0 28520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_22
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_34
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_41
timestamp 1676037725
transform 1 0 4876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1676037725
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1676037725
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1676037725
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1676037725
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1676037725
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_179
timestamp 1676037725
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_200
timestamp 1676037725
transform 1 0 19504 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1676037725
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1676037725
transform 1 0 23276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_270
timestamp 1676037725
transform 1 0 25944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 1676037725
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_43
timestamp 1676037725
transform 1 0 5060 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1676037725
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_63
timestamp 1676037725
transform 1 0 6900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1676037725
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1676037725
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1676037725
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1676037725
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1676037725
transform 1 0 21528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1676037725
transform 1 0 23092 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1676037725
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_36
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_42
timestamp 1676037725
transform 1 0 4968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1676037725
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1676037725
transform 1 0 7636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1676037725
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_99
timestamp 1676037725
transform 1 0 10212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1676037725
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1676037725
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_176
timestamp 1676037725
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_190
timestamp 1676037725
transform 1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_208
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_233
timestamp 1676037725
transform 1 0 22540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_241
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1676037725
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1676037725
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_43
timestamp 1676037725
transform 1 0 5060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1676037725
transform 1 0 5796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1676037725
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_66
timestamp 1676037725
transform 1 0 7176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_72
timestamp 1676037725
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1676037725
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_104
timestamp 1676037725
transform 1 0 10672 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_113
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1676037725
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_130
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_204
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1676037725
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_274
timestamp 1676037725
transform 1 0 26312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1676037725
transform 1 0 28336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1676037725
transform 1 0 2208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_32
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_40
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1676037725
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_77
timestamp 1676037725
transform 1 0 8188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1676037725
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1676037725
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1676037725
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1676037725
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1676037725
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_14
timestamp 1676037725
transform 1 0 2392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_22
timestamp 1676037725
transform 1 0 3128 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_35
timestamp 1676037725
transform 1 0 4324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_42
timestamp 1676037725
transform 1 0 4968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1676037725
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_90
timestamp 1676037725
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1676037725
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_113
timestamp 1676037725
transform 1 0 11500 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1676037725
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1676037725
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_204
timestamp 1676037725
transform 1 0 19872 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1676037725
transform 1 0 21988 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1676037725
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_270
timestamp 1676037725
transform 1 0 25944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_28
timestamp 1676037725
transform 1 0 3680 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp 1676037725
transform 1 0 4232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_49
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1676037725
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1676037725
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1676037725
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1676037725
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1676037725
transform 1 0 12144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_289
timestamp 1676037725
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_296
timestamp 1676037725
transform 1 0 28336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1676037725
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1676037725
transform 1 0 4968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_50
timestamp 1676037725
transform 1 0 5704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1676037725
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_101
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1676037725
transform 1 0 11316 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_149
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_157
timestamp 1676037725
transform 1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1676037725
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1676037725
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_243
timestamp 1676037725
transform 1 0 23460 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_13
timestamp 1676037725
transform 1 0 2300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_30
timestamp 1676037725
transform 1 0 3864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_66
timestamp 1676037725
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1676037725
transform 1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1676037725
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_212
timestamp 1676037725
transform 1 0 20608 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_252
timestamp 1676037725
transform 1 0 24288 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_260
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_296
timestamp 1676037725
transform 1 0 28336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_12
timestamp 1676037725
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_20
timestamp 1676037725
transform 1 0 2944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1676037725
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_49
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1676037725
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_92
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1676037725
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_224
timestamp 1676037725
transform 1 0 21712 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1676037725
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1676037725
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_18
timestamp 1676037725
transform 1 0 2760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_120
timestamp 1676037725
transform 1 0 12144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_127
timestamp 1676037725
transform 1 0 12788 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1676037725
transform 1 0 14260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1676037725
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_242
timestamp 1676037725
transform 1 0 23368 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1676037725
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_294
timestamp 1676037725
transform 1 0 28152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1676037725
transform 1 0 28520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_13
timestamp 1676037725
transform 1 0 2300 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1676037725
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_45
timestamp 1676037725
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_56
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1676037725
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1676037725
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_99
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1676037725
transform 1 0 10948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1676037725
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1676037725
transform 1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_184
timestamp 1676037725
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_234
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1676037725
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_10
timestamp 1676037725
transform 1 0 2024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_44
timestamp 1676037725
transform 1 0 5152 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1676037725
transform 1 0 5704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1676037725
transform 1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_74
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_88
timestamp 1676037725
transform 1 0 9200 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1676037725
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_134
timestamp 1676037725
transform 1 0 13432 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_140
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1676037725
transform 1 0 25668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_288
timestamp 1676037725
transform 1 0 27600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1676037725
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_13
timestamp 1676037725
transform 1 0 2300 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1676037725
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_35
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1676037725
transform 1 0 5244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1676037725
transform 1 0 7912 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_115
timestamp 1676037725
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1676037725
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1676037725
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1676037725
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1676037725
transform 1 0 26220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_293
timestamp 1676037725
transform 1 0 28060 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_8
timestamp 1676037725
transform 1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_20
timestamp 1676037725
transform 1 0 2944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_28
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_37
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1676037725
transform 1 0 7084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_77
timestamp 1676037725
transform 1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_90
timestamp 1676037725
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_128
timestamp 1676037725
transform 1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_197
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1676037725
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_256
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1676037725
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_290
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1676037725
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_18
timestamp 1676037725
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_45
timestamp 1676037725
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_51
timestamp 1676037725
transform 1 0 5796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1676037725
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1676037725
transform 1 0 6808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_66
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1676037725
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1676037725
transform 1 0 12972 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_148
timestamp 1676037725
transform 1 0 14720 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1676037725
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_291
timestamp 1676037725
transform 1 0 27876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1676037725
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1676037725
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1676037725
transform 1 0 13340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_141
timestamp 1676037725
transform 1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1676037725
transform 1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_230
timestamp 1676037725
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_269
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1676037725
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_12
timestamp 1676037725
transform 1 0 2208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_18
timestamp 1676037725
transform 1 0 2760 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1676037725
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_52
timestamp 1676037725
transform 1 0 5888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1676037725
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_94
timestamp 1676037725
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1676037725
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_158
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_164
timestamp 1676037725
transform 1 0 16192 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_280
timestamp 1676037725
transform 1 0 26864 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1676037725
transform 1 0 2392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_26
timestamp 1676037725
transform 1 0 3496 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_36
timestamp 1676037725
transform 1 0 4416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_46
timestamp 1676037725
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_77
timestamp 1676037725
transform 1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1676037725
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1676037725
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1676037725
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_189
timestamp 1676037725
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 1676037725
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_10
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_37
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_55
timestamp 1676037725
transform 1 0 6164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1676037725
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_116
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_122
timestamp 1676037725
transform 1 0 12328 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_126
timestamp 1676037725
transform 1 0 12696 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_171
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1676037725
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_240
timestamp 1676037725
transform 1 0 23184 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_246
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_8
timestamp 1676037725
transform 1 0 1840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_12
timestamp 1676037725
transform 1 0 2208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_17
timestamp 1676037725
transform 1 0 2668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_30
timestamp 1676037725
transform 1 0 3864 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_43
timestamp 1676037725
transform 1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1676037725
transform 1 0 7176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1676037725
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1676037725
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_145
timestamp 1676037725
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1676037725
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_185
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_252
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_260
timestamp 1676037725
transform 1 0 25024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1676037725
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1676037725
transform 1 0 2668 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_37
timestamp 1676037725
transform 1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_49
timestamp 1676037725
transform 1 0 5612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_68
timestamp 1676037725
transform 1 0 7360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_101
timestamp 1676037725
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1676037725
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_130
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_157
timestamp 1676037725
transform 1 0 15548 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_168
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_176
timestamp 1676037725
transform 1 0 17296 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_188
timestamp 1676037725
transform 1 0 18400 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1676037725
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_271
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_22
timestamp 1676037725
transform 1 0 3128 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1676037725
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_68
timestamp 1676037725
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_78
timestamp 1676037725
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_84
timestamp 1676037725
transform 1 0 8832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1676037725
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_102
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_122
timestamp 1676037725
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1676037725
transform 1 0 12972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_176
timestamp 1676037725
transform 1 0 17296 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1676037725
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1676037725
transform 1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_207
timestamp 1676037725
transform 1 0 20148 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1676037725
transform 1 0 22540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_244
timestamp 1676037725
transform 1 0 23552 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_268
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_12
timestamp 1676037725
transform 1 0 2208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1676037725
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_40
timestamp 1676037725
transform 1 0 4784 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_67
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_75
timestamp 1676037725
transform 1 0 8004 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_94
timestamp 1676037725
transform 1 0 9752 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_116
timestamp 1676037725
transform 1 0 11776 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1676037725
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_187
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1676037725
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1676037725
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_31
timestamp 1676037725
transform 1 0 3956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1676037725
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1676037725
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_78
timestamp 1676037725
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1676037725
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1676037725
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_130
timestamp 1676037725
transform 1 0 13064 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_176
timestamp 1676037725
transform 1 0 17296 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_185
timestamp 1676037725
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_194
timestamp 1676037725
transform 1 0 18952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_203
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_234
timestamp 1676037725
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1676037725
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_10
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1676037725
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1676037725
transform 1 0 4784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_50
timestamp 1676037725
transform 1 0 5704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_60
timestamp 1676037725
transform 1 0 6624 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_68
timestamp 1676037725
transform 1 0 7360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_76
timestamp 1676037725
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_96
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_126
timestamp 1676037725
transform 1 0 12696 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_132
timestamp 1676037725
transform 1 0 13248 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1676037725
transform 1 0 14812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1676037725
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_183
timestamp 1676037725
transform 1 0 17940 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_227
timestamp 1676037725
transform 1 0 21988 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1676037725
transform 1 0 23092 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_270
timestamp 1676037725
transform 1 0 25944 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_12
timestamp 1676037725
transform 1 0 2208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_36
timestamp 1676037725
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_74
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_78
timestamp 1676037725
transform 1 0 8280 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_88
timestamp 1676037725
transform 1 0 9200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_101
timestamp 1676037725
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1676037725
transform 1 0 12880 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1676037725
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_152
timestamp 1676037725
transform 1 0 15088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1676037725
transform 1 0 17204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_182
timestamp 1676037725
transform 1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_190
timestamp 1676037725
transform 1 0 18584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1676037725
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1676037725
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_231
timestamp 1676037725
transform 1 0 22356 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_239
timestamp 1676037725
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_256
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_40
timestamp 1676037725
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1676037725
transform 1 0 6992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_73
timestamp 1676037725
transform 1 0 7820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1676037725
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_93
timestamp 1676037725
transform 1 0 9660 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_116
timestamp 1676037725
transform 1 0 11776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1676037725
transform 1 0 12880 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_132
timestamp 1676037725
transform 1 0 13248 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_152
timestamp 1676037725
transform 1 0 15088 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1676037725
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_187
timestamp 1676037725
transform 1 0 18308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_211
timestamp 1676037725
transform 1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_229
timestamp 1676037725
transform 1 0 22172 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1676037725
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_291
timestamp 1676037725
transform 1 0 27876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_10
timestamp 1676037725
transform 1 0 2024 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_33
timestamp 1676037725
transform 1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_46
timestamp 1676037725
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1676037725
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_64
timestamp 1676037725
transform 1 0 6992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_68
timestamp 1676037725
transform 1 0 7360 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_75
timestamp 1676037725
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_84
timestamp 1676037725
transform 1 0 8832 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1676037725
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_132
timestamp 1676037725
transform 1 0 13248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1676037725
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_192
timestamp 1676037725
transform 1 0 18768 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_198
timestamp 1676037725
transform 1 0 19320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_212
timestamp 1676037725
transform 1 0 20608 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1676037725
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_250
timestamp 1676037725
transform 1 0 24104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1676037725
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_47
timestamp 1676037725
transform 1 0 5428 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_61
timestamp 1676037725
transform 1 0 6716 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_71
timestamp 1676037725
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1676037725
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1676037725
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_104
timestamp 1676037725
transform 1 0 10672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_128
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_154
timestamp 1676037725
transform 1 0 15272 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_170
timestamp 1676037725
transform 1 0 16744 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1676037725
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1676037725
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_204
timestamp 1676037725
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_211
timestamp 1676037725
transform 1 0 20516 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_217
timestamp 1676037725
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_229
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1676037725
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1676037725
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_258
timestamp 1676037725
transform 1 0 24840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_270
timestamp 1676037725
transform 1 0 25944 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1676037725
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_45
timestamp 1676037725
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1676037725
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_68
timestamp 1676037725
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1676037725
transform 1 0 8188 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1676037725
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1676037725
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_103
timestamp 1676037725
transform 1 0 10580 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_119
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_139
timestamp 1676037725
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1676037725
transform 1 0 14536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_176
timestamp 1676037725
transform 1 0 17296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1676037725
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_197
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_204
timestamp 1676037725
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_211
timestamp 1676037725
transform 1 0 20516 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_243
timestamp 1676037725
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1676037725
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_270
timestamp 1676037725
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1676037725
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_50
timestamp 1676037725
transform 1 0 5704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_58
timestamp 1676037725
transform 1 0 6440 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_66
timestamp 1676037725
transform 1 0 7176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1676037725
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1676037725
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_92
timestamp 1676037725
transform 1 0 9568 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_105
timestamp 1676037725
transform 1 0 10764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_113
timestamp 1676037725
transform 1 0 11500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_128
timestamp 1676037725
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_157
timestamp 1676037725
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1676037725
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1676037725
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_235
timestamp 1676037725
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_242
timestamp 1676037725
transform 1 0 23368 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1676037725
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1676037725
transform 1 0 2208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_36
timestamp 1676037725
transform 1 0 4416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_45
timestamp 1676037725
transform 1 0 5244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1676037725
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_66
timestamp 1676037725
transform 1 0 7176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_76
timestamp 1676037725
transform 1 0 8096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_84
timestamp 1676037725
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_90
timestamp 1676037725
transform 1 0 9384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_103
timestamp 1676037725
transform 1 0 10580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1676037725
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1676037725
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1676037725
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_140
timestamp 1676037725
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_146
timestamp 1676037725
transform 1 0 14536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1676037725
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1676037725
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_178
timestamp 1676037725
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1676037725
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_195
timestamp 1676037725
transform 1 0 19044 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_202
timestamp 1676037725
transform 1 0 19688 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_211
timestamp 1676037725
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1676037725
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_250
timestamp 1676037725
transform 1 0 24104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_257
timestamp 1676037725
transform 1 0 24748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_286
timestamp 1676037725
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_9
timestamp 1676037725
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1676037725
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_50
timestamp 1676037725
transform 1 0 5704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_59
timestamp 1676037725
transform 1 0 6532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_68
timestamp 1676037725
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1676037725
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_91
timestamp 1676037725
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_117
timestamp 1676037725
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_127
timestamp 1676037725
transform 1 0 12788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1676037725
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_151
timestamp 1676037725
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1676037725
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_167
timestamp 1676037725
transform 1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_173
timestamp 1676037725
transform 1 0 17020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_183
timestamp 1676037725
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1676037725
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_202
timestamp 1676037725
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_216
timestamp 1676037725
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1676037725
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1676037725
transform 1 0 22264 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_271
timestamp 1676037725
transform 1 0 26036 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_279
timestamp 1676037725
transform 1 0 26772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1676037725
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1676037725
transform 1 0 2116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_33
timestamp 1676037725
transform 1 0 4140 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_37
timestamp 1676037725
transform 1 0 4508 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_43
timestamp 1676037725
transform 1 0 5060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1676037725
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_67
timestamp 1676037725
transform 1 0 7268 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_79
timestamp 1676037725
transform 1 0 8372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_88
timestamp 1676037725
transform 1 0 9200 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1676037725
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_119
timestamp 1676037725
transform 1 0 12052 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_133
timestamp 1676037725
transform 1 0 13340 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1676037725
transform 1 0 14536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_157
timestamp 1676037725
transform 1 0 15548 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_187
timestamp 1676037725
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_198
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_229
timestamp 1676037725
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_246
timestamp 1676037725
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_267
timestamp 1676037725
transform 1 0 25668 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1676037725
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1676037725
transform 1 0 27416 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1676037725
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_36
timestamp 1676037725
transform 1 0 4416 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_44
timestamp 1676037725
transform 1 0 5152 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_76
timestamp 1676037725
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_91
timestamp 1676037725
transform 1 0 9476 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_100
timestamp 1676037725
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_118
timestamp 1676037725
transform 1 0 11960 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1676037725
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_154
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_178
timestamp 1676037725
transform 1 0 17480 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_186
timestamp 1676037725
transform 1 0 18216 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1676037725
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1676037725
transform 1 0 21712 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_231
timestamp 1676037725
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1676037725
transform 1 0 23000 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_271
timestamp 1676037725
transform 1 0 26036 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_279
timestamp 1676037725
transform 1 0 26772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_296
timestamp 1676037725
transform 1 0 28336 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_25
timestamp 1676037725
transform 1 0 3404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_35
timestamp 1676037725
transform 1 0 4324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_44
timestamp 1676037725
transform 1 0 5152 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_48
timestamp 1676037725
transform 1 0 5520 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1676037725
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_65
timestamp 1676037725
transform 1 0 7084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_73
timestamp 1676037725
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_82
timestamp 1676037725
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_91
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_127
timestamp 1676037725
transform 1 0 12788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_136
timestamp 1676037725
transform 1 0 13616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_142
timestamp 1676037725
transform 1 0 14168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_157
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_175
timestamp 1676037725
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_192
timestamp 1676037725
transform 1 0 18768 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1676037725
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_264
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_271
timestamp 1676037725
transform 1 0 26036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1676037725
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_286
timestamp 1676037725
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1676037725
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_37
timestamp 1676037725
transform 1 0 4508 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_46
timestamp 1676037725
transform 1 0 5336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_55
timestamp 1676037725
transform 1 0 6164 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_64
timestamp 1676037725
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_73
timestamp 1676037725
transform 1 0 7820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1676037725
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_108
timestamp 1676037725
transform 1 0 11040 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_114
timestamp 1676037725
transform 1 0 11592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_131
timestamp 1676037725
transform 1 0 13156 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_147
timestamp 1676037725
transform 1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_167
timestamp 1676037725
transform 1 0 16468 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_173
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1676037725
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_215
timestamp 1676037725
transform 1 0 20884 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_223
timestamp 1676037725
transform 1 0 21620 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_241
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1676037725
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1676037725
transform 1 0 27232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_291
timestamp 1676037725
transform 1 0 27876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1676037725
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1676037725
transform 1 0 6808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_72
timestamp 1676037725
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_86
timestamp 1676037725
transform 1 0 9016 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_120
timestamp 1676037725
transform 1 0 12144 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_142
timestamp 1676037725
transform 1 0 14168 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_152
timestamp 1676037725
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1676037725
transform 1 0 18308 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_191
timestamp 1676037725
transform 1 0 18676 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_202
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_209
timestamp 1676037725
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1676037725
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_230
timestamp 1676037725
transform 1 0 22264 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_259
timestamp 1676037725
transform 1 0 24932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_266
timestamp 1676037725
transform 1 0 25576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1676037725
transform 1 0 27416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 1676037725
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_40
timestamp 1676037725
transform 1 0 4784 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_48
timestamp 1676037725
transform 1 0 5520 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_55
timestamp 1676037725
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_64
timestamp 1676037725
transform 1 0 6992 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1676037725
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1676037725
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_129
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_159
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1676037725
transform 1 0 16560 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_184
timestamp 1676037725
transform 1 0 18032 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp 1676037725
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_216
timestamp 1676037725
transform 1 0 20976 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_236
timestamp 1676037725
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_243
timestamp 1676037725
transform 1 0 23460 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_258
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_272
timestamp 1676037725
transform 1 0 26128 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_279
timestamp 1676037725
transform 1 0 26772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1676037725
transform 1 0 27416 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_293
timestamp 1676037725
transform 1 0 28060 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_11
timestamp 1676037725
transform 1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_65
timestamp 1676037725
transform 1 0 7084 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_74
timestamp 1676037725
transform 1 0 7912 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_83
timestamp 1676037725
transform 1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_103
timestamp 1676037725
transform 1 0 10580 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_126
timestamp 1676037725
transform 1 0 12696 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_146
timestamp 1676037725
transform 1 0 14536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_174
timestamp 1676037725
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_194
timestamp 1676037725
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1676037725
transform 1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1676037725
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_250
timestamp 1676037725
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_257
timestamp 1676037725
transform 1 0 24748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_271
timestamp 1676037725
transform 1 0 26036 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1676037725
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_19
timestamp 1676037725
transform 1 0 2852 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1676037725
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_37
timestamp 1676037725
transform 1 0 4508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_46
timestamp 1676037725
transform 1 0 5336 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_55
timestamp 1676037725
transform 1 0 6164 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_64
timestamp 1676037725
transform 1 0 6992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_74
timestamp 1676037725
transform 1 0 7912 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1676037725
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1676037725
transform 1 0 9476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_98
timestamp 1676037725
transform 1 0 10120 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_102
timestamp 1676037725
transform 1 0 10488 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_120
timestamp 1676037725
transform 1 0 12144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_124
timestamp 1676037725
transform 1 0 12512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_128
timestamp 1676037725
transform 1 0 12880 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_163
timestamp 1676037725
transform 1 0 16100 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 1676037725
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1676037725
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_215
timestamp 1676037725
transform 1 0 20884 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_238
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1676037725
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_278
timestamp 1676037725
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_285
timestamp 1676037725
transform 1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_292
timestamp 1676037725
transform 1 0 27968 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_298
timestamp 1676037725
transform 1 0 28520 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_16
timestamp 1676037725
transform 1 0 2576 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_20
timestamp 1676037725
transform 1 0 2944 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_26
timestamp 1676037725
transform 1 0 3496 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_29
timestamp 1676037725
transform 1 0 3772 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_36
timestamp 1676037725
transform 1 0 4416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1676037725
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_64
timestamp 1676037725
transform 1 0 6992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_73
timestamp 1676037725
transform 1 0 7820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_82
timestamp 1676037725
transform 1 0 8648 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1676037725
transform 1 0 8924 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 1676037725
transform 1 0 9568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_101
timestamp 1676037725
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1676037725
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1676037725
transform 1 0 11960 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_128
timestamp 1676037725
transform 1 0 12880 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_138
timestamp 1676037725
transform 1 0 13800 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1676037725
transform 1 0 14076 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_146
timestamp 1676037725
transform 1 0 14536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_174
timestamp 1676037725
transform 1 0 17112 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_194
timestamp 1676037725
transform 1 0 18952 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_197
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1676037725
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_244
timestamp 1676037725
transform 1 0 23552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_258
timestamp 1676037725
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_265
timestamp 1676037725
transform 1 0 25484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_272
timestamp 1676037725
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1676037725
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 28888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 28888 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0903_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0905_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6072 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0909_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0912_
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0914_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0915_
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0917_
timestamp 1676037725
transform 1 0 2944 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__or3b_4  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8372 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0920_
timestamp 1676037725
transform 1 0 7728 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1676037725
transform 1 0 24472 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_4  _0924_
timestamp 1676037725
transform 1 0 10396 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_1  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0926_
timestamp 1676037725
transform 1 0 5060 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0927_
timestamp 1676037725
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0928_
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0932_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0933_
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0936_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0937_
timestamp 1676037725
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0940_
timestamp 1676037725
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0941_
timestamp 1676037725
transform 1 0 6808 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0942_
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _0943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1676037725
transform 1 0 18400 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0945_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11500 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _0948_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_2  _0950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1676037725
transform 1 0 15272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0955_
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0957_
timestamp 1676037725
transform 1 0 14536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1676037725
transform 1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0959_
timestamp 1676037725
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0960_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1676037725
transform 1 0 16652 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0962_
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1676037725
transform 1 0 17480 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0966_
timestamp 1676037725
transform 1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_4  _0967_
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1676037725
transform 1 0 17664 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0969_
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1676037725
transform 1 0 17940 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0971_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _0972_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0975_
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_4  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _0977_
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0978_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0979_
timestamp 1676037725
transform 1 0 10672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _0980_
timestamp 1676037725
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0981_
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0983_
timestamp 1676037725
transform 1 0 10120 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0984_
timestamp 1676037725
transform 1 0 12144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0985_
timestamp 1676037725
transform 1 0 15548 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9936 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0987_
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0988_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0989_
timestamp 1676037725
transform 1 0 9844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0990_
timestamp 1676037725
transform 1 0 8280 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0992_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0994_
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0997_
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0998_
timestamp 1676037725
transform 1 0 17020 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0999_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1676037725
transform 1 0 18492 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1002_
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1003_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1004_
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1006_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1007_
timestamp 1676037725
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1010_
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9936 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1012_
timestamp 1676037725
transform 1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1676037725
transform 1 0 10580 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1014_
timestamp 1676037725
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1016_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1018_
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1019_
timestamp 1676037725
transform 1 0 15456 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1020_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1676037725
transform 1 0 17664 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1023_
timestamp 1676037725
transform 1 0 17388 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1024_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1676037725
transform 1 0 14720 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1027_
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1028_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1029_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1030_
timestamp 1676037725
transform 1 0 14352 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1032_
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1033_
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_2  _1034_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1035_
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1036_
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 1676037725
transform 1 0 16008 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1038_
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1039_
timestamp 1676037725
transform 1 0 12880 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1040_
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1041_
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1042_
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1043_
timestamp 1676037725
transform 1 0 12144 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1045_
timestamp 1676037725
transform 1 0 11868 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1047_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1048_
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1049_
timestamp 1676037725
transform 1 0 17756 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_2  _1050_
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1051_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1052_
timestamp 1676037725
transform 1 0 8004 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1053_
timestamp 1676037725
transform 1 0 14628 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1054_
timestamp 1676037725
transform 1 0 15824 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1055_
timestamp 1676037725
transform 1 0 13340 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1056_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1058_
timestamp 1676037725
transform 1 0 9568 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1059_
timestamp 1676037725
transform 1 0 15272 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1060_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1061_
timestamp 1676037725
transform 1 0 18768 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1062_
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1063_
timestamp 1676037725
transform 1 0 14444 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1064_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1066_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1067_
timestamp 1676037725
transform 1 0 11684 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1068_
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1676037725
transform 1 0 17112 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12420 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1072_
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1073_
timestamp 1676037725
transform 1 0 16192 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1074_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1075_
timestamp 1676037725
transform 1 0 17664 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1076_
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1077_
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1078_
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1080_
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1081_
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1082_
timestamp 1676037725
transform 1 0 14352 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1086_
timestamp 1676037725
transform 1 0 6992 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1676037725
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1088_
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1089_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1090_
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1091_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1093_
timestamp 1676037725
transform 1 0 17940 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1094_
timestamp 1676037725
transform 1 0 12880 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1095_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1096_
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1097_
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1098_
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1099_
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1100_
timestamp 1676037725
transform 1 0 14720 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1102_
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1103_
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1104_
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1105_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1106_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1107_
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1108_
timestamp 1676037725
transform 1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1109_
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1110_
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1112_
timestamp 1676037725
transform 1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1113_
timestamp 1676037725
transform 1 0 17204 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 1676037725
transform 1 0 13616 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1115_
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1116_
timestamp 1676037725
transform 1 0 14996 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1117_
timestamp 1676037725
transform 1 0 11776 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1118_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1119_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1120_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_2  _1121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1124_
timestamp 1676037725
transform 1 0 8740 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1125_
timestamp 1676037725
transform 1 0 6624 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6716 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1127_
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1128_
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1129_
timestamp 1676037725
transform 1 0 19780 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1130_
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1131_
timestamp 1676037725
transform 1 0 15456 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 1676037725
transform 1 0 14812 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1133_
timestamp 1676037725
transform 1 0 17388 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1134_
timestamp 1676037725
transform 1 0 17480 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1136_
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1137_
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1138_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1139_
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1140_
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1141_
timestamp 1676037725
transform 1 0 11868 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1142_
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1143_
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 1676037725
transform 1 0 9660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1145_
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1146_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1147_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1148_
timestamp 1676037725
transform 1 0 11684 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1149_
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1150_
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1151_
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1152_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1154_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1155_
timestamp 1676037725
transform 1 0 16836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1156_
timestamp 1676037725
transform 1 0 13524 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1157_
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1160_
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1161_
timestamp 1676037725
transform 1 0 6440 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1162_
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1163_
timestamp 1676037725
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1168_
timestamp 1676037725
transform 1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1676037725
transform 1 0 4416 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1170_
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1676037725
transform 1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4416 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1173_
timestamp 1676037725
transform 1 0 5520 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o22ai_2  _1175_
timestamp 1676037725
transform 1 0 7912 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1176_
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1178_
timestamp 1676037725
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1179_
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1180_
timestamp 1676037725
transform 1 0 14904 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1181_
timestamp 1676037725
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1183_
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1185_
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1186_
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1188_
timestamp 1676037725
transform 1 0 8832 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1189_
timestamp 1676037725
transform 1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1190_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1191_
timestamp 1676037725
transform 1 0 19872 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1192_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1193_
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1194_
timestamp 1676037725
transform 1 0 12880 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1195_
timestamp 1676037725
transform 1 0 15824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1198_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1676037725
transform 1 0 9384 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1201_
timestamp 1676037725
transform 1 0 1748 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1676037725
transform 1 0 27600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1204_
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _1207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1676037725
transform 1 0 1748 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1209_
timestamp 1676037725
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1676037725
transform 1 0 5244 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1211_
timestamp 1676037725
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1213_
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1676037725
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1215_
timestamp 1676037725
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1216_
timestamp 1676037725
transform 1 0 4416 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1217_
timestamp 1676037725
transform 1 0 4968 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1218_
timestamp 1676037725
transform 1 0 6992 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2392 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1223_
timestamp 1676037725
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1224_
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 1676037725
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_2  _1229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_1  _1230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2760 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _1232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1676037725
transform 1 0 8280 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1234_
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1235_
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_4  _1236_
timestamp 1676037725
transform 1 0 10396 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1676037725
transform 1 0 2576 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1238_
timestamp 1676037725
transform 1 0 7452 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1239_
timestamp 1676037725
transform 1 0 4324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1240_
timestamp 1676037725
transform 1 0 3220 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1242_
timestamp 1676037725
transform 1 0 5060 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1676037725
transform 1 0 3220 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _1245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o32ai_1  _1246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1247_
timestamp 1676037725
transform 1 0 1748 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4692 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1250_
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1251_
timestamp 1676037725
transform 1 0 5152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1253_
timestamp 1676037725
transform 1 0 5336 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1254_
timestamp 1676037725
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1255_
timestamp 1676037725
transform 1 0 7728 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1258_
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1259_
timestamp 1676037725
transform 1 0 6532 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_4  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _1261_
timestamp 1676037725
transform 1 0 7544 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1262_
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1264_
timestamp 1676037725
transform 1 0 4968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1265_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1266_
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1267_
timestamp 1676037725
transform 1 0 4324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1268_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1270_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1272_
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1273_
timestamp 1676037725
transform 1 0 7452 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1274_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1275_
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1276_
timestamp 1676037725
transform 1 0 4784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1277_
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1278_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1279_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1280_
timestamp 1676037725
transform 1 0 5704 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1282_
timestamp 1676037725
transform 1 0 6072 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1283_
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1284_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1285_
timestamp 1676037725
transform 1 0 4784 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1286_
timestamp 1676037725
transform 1 0 6532 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1676037725
transform 1 0 26036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1288_
timestamp 1676037725
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1289_
timestamp 1676037725
transform 1 0 5612 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1290_
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1291_
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1676037725
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1294_
timestamp 1676037725
transform 1 0 5152 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _1295_
timestamp 1676037725
transform 1 0 4140 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1676037725
transform 1 0 1748 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1297_
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 1676037725
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1299_
timestamp 1676037725
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1300_
timestamp 1676037725
transform 1 0 2852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1301_
timestamp 1676037725
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1302_
timestamp 1676037725
transform 1 0 4416 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1303_
timestamp 1676037725
transform 1 0 5060 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1304_
timestamp 1676037725
transform 1 0 6532 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1305_
timestamp 1676037725
transform 1 0 5612 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1306_
timestamp 1676037725
transform 1 0 6624 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1307_
timestamp 1676037725
transform 1 0 5152 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1310_
timestamp 1676037725
transform 1 0 5704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1311_
timestamp 1676037725
transform 1 0 2392 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1314_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1315_
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1317_
timestamp 1676037725
transform 1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1320_
timestamp 1676037725
transform 1 0 3680 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1321_
timestamp 1676037725
transform 1 0 5520 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1322_
timestamp 1676037725
transform 1 0 5244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1323_
timestamp 1676037725
transform 1 0 3128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1324_
timestamp 1676037725
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1325_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1326_
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1327_
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1328_
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1330_
timestamp 1676037725
transform 1 0 3956 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1331_
timestamp 1676037725
transform 1 0 21344 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1676037725
transform 1 0 21988 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1333_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1334_
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1335_
timestamp 1676037725
transform 1 0 9568 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1676037725
transform 1 0 9384 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1337_
timestamp 1676037725
transform 1 0 1748 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1676037725
transform 1 0 27784 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1676037725
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1340_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1676037725
transform 1 0 23828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1676037725
transform 1 0 25760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1343_
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1676037725
transform 1 0 26404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_
timestamp 1676037725
transform 1 0 7728 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1348_
timestamp 1676037725
transform 1 0 9844 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1349_
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1350_
timestamp 1676037725
transform 1 0 5244 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 1676037725
transform 1 0 26956 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1353_
timestamp 1676037725
transform 1 0 26404 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1354_
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1676037725
transform 1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1357_
timestamp 1676037725
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1358_
timestamp 1676037725
transform 1 0 7360 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1359_
timestamp 1676037725
transform 1 0 8188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1676037725
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1361_
timestamp 1676037725
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1362_
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1364_
timestamp 1676037725
transform 1 0 8648 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1676037725
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1676037725
transform 1 0 4692 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1676037725
transform 1 0 5520 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1676037725
transform 1 0 5796 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1676037725
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1372_
timestamp 1676037725
transform 1 0 6808 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1676037725
transform 1 0 7544 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1374_
timestamp 1676037725
transform 1 0 8648 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1376_
timestamp 1676037725
transform 1 0 11776 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1676037725
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1378_
timestamp 1676037725
transform 1 0 12788 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1379_
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1380_
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1381_
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1382_
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1384_
timestamp 1676037725
transform 1 0 20792 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1385_
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1386_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1387_
timestamp 1676037725
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1388_
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1390_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1391_
timestamp 1676037725
transform 1 0 21620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1676037725
transform 1 0 21620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1397_
timestamp 1676037725
transform 1 0 18032 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1398_
timestamp 1676037725
transform 1 0 15272 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1400_
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1676037725
transform 1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1402_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1403_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1404_
timestamp 1676037725
transform 1 0 20976 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1406_
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1411_
timestamp 1676037725
transform 1 0 19964 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1412_
timestamp 1676037725
transform 1 0 23276 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1413_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1676037725
transform 1 0 20332 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1415_
timestamp 1676037725
transform 1 0 18216 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1417_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1418_
timestamp 1676037725
transform 1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1419_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1420_
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1421_
timestamp 1676037725
transform 1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1676037725
transform 1 0 12420 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1423_
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1424_
timestamp 1676037725
transform 1 0 15732 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1425_
timestamp 1676037725
transform 1 0 18400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1426_
timestamp 1676037725
transform 1 0 18032 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1676037725
transform 1 0 20056 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1428_
timestamp 1676037725
transform 1 0 18032 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1676037725
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1676037725
transform 1 0 12972 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1431_
timestamp 1676037725
transform 1 0 14260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1432_
timestamp 1676037725
transform 1 0 10120 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1434_
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1435_
timestamp 1676037725
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1436_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1438_
timestamp 1676037725
transform 1 0 12052 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1676037725
transform 1 0 11224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1440_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1676037725
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1442_
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1444_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1676037725
transform 1 0 7728 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1676037725
transform 1 0 9200 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1448_
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1449_
timestamp 1676037725
transform 1 0 6716 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1676037725
transform 1 0 27784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1451_
timestamp 1676037725
transform 1 0 7360 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1452_
timestamp 1676037725
transform 1 0 27784 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1453_
timestamp 1676037725
transform 1 0 10212 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1676037725
transform 1 0 25392 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1455_
timestamp 1676037725
transform 1 0 6900 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1676037725
transform 1 0 27784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1457_
timestamp 1676037725
transform 1 0 10672 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1676037725
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1459_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1676037725
transform 1 0 13248 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1676037725
transform 1 0 17848 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1462_
timestamp 1676037725
transform 1 0 7176 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1676037725
transform 1 0 27600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1464_
timestamp 1676037725
transform 1 0 9568 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1676037725
transform 1 0 27140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1466_
timestamp 1676037725
transform 1 0 14260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1676037725
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1676037725
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1676037725
transform 1 0 14076 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1676037725
transform 1 0 17756 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1472_
timestamp 1676037725
transform 1 0 14076 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1676037725
transform 1 0 12604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1474_
timestamp 1676037725
transform 1 0 13248 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1676037725
transform 1 0 23368 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1476_
timestamp 1676037725
transform 1 0 12328 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1676037725
transform 1 0 23276 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1478_
timestamp 1676037725
transform 1 0 14536 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1676037725
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1676037725
transform 1 0 14536 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1676037725
transform 1 0 20056 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1676037725
transform 1 0 19136 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1676037725
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1486_
timestamp 1676037725
transform 1 0 13248 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1676037725
transform 1 0 21160 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1488_
timestamp 1676037725
transform 1 0 12788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1489_
timestamp 1676037725
transform 1 0 18400 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1491_
timestamp 1676037725
transform 1 0 18400 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1676037725
transform 1 0 20700 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1676037725
transform 1 0 17020 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1676037725
transform 1 0 19412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1495_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1676037725
transform 1 0 19596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 1676037725
transform 1 0 18492 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1499_
timestamp 1676037725
transform 1 0 20792 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1501_
timestamp 1676037725
transform 1 0 19872 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1676037725
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1503_
timestamp 1676037725
transform 1 0 21620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1676037725
transform 1 0 24472 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1505_
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1676037725
transform 1 0 19596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1676037725
transform 1 0 23828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1676037725
transform 1 0 20240 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1509_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 1676037725
transform 1 0 20700 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1511_
timestamp 1676037725
transform 1 0 21160 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1512_
timestamp 1676037725
transform 1 0 20148 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1513_
timestamp 1676037725
transform 1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1514_
timestamp 1676037725
transform 1 0 21344 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1515_
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1516_
timestamp 1676037725
transform 1 0 20516 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1518_
timestamp 1676037725
transform 1 0 20884 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1519_
timestamp 1676037725
transform 1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1521_
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1676037725
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1524_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1526_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1528_
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1529_
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1530_
timestamp 1676037725
transform 1 0 19412 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1676037725
transform 1 0 20240 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1532_
timestamp 1676037725
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1533_
timestamp 1676037725
transform 1 0 17480 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1534_
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1535_
timestamp 1676037725
transform 1 0 18492 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1676037725
transform 1 0 20240 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1537_
timestamp 1676037725
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1538_
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1539_
timestamp 1676037725
transform 1 0 14720 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1541_
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1676037725
transform 1 0 16192 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1543_
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1544_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1676037725
transform 1 0 11408 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1676037725
transform 1 0 9200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1548_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1676037725
transform 1 0 8372 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1676037725
transform 1 0 24748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1676037725
transform 1 0 7360 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1676037725
transform 1 0 20884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1554_
timestamp 1676037725
transform 1 0 7728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1676037725
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1556_
timestamp 1676037725
transform 1 0 7820 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1557_
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1558_
timestamp 1676037725
transform 1 0 10120 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1676037725
transform 1 0 10120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1560_
timestamp 1676037725
transform 1 0 9384 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1676037725
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1562_
timestamp 1676037725
transform 1 0 7912 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1676037725
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1564_
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1676037725
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1566_
timestamp 1676037725
transform 1 0 8372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 1676037725
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1568_
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1572_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1676037725
transform 1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1576_
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1577_
timestamp 1676037725
transform 1 0 20608 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1579_
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 1676037725
transform 1 0 18492 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1676037725
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1583_
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1587_
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1676037725
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1589_
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1590_
timestamp 1676037725
transform 1 0 20608 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1591_
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1592_
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1593_
timestamp 1676037725
transform 1 0 23552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1594_
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1595_
timestamp 1676037725
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1596_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1676037725
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1676037725
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1676037725
transform 1 0 20240 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1601_
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1602_
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1603_
timestamp 1676037725
transform 1 0 23276 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1604_
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1605_
timestamp 1676037725
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1606_
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1607_
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1608_
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1609_
timestamp 1676037725
transform 1 0 16100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1611_
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1613_
timestamp 1676037725
transform 1 0 10396 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1615_
timestamp 1676037725
transform 1 0 9476 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1676037725
transform 1 0 26404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1617_
timestamp 1676037725
transform 1 0 11500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1676037725
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1619_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1620_
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1621_
timestamp 1676037725
transform 1 0 14076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1622_
timestamp 1676037725
transform 1 0 15088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1623_
timestamp 1676037725
transform 1 0 12420 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1676037725
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1625_
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1676037725
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1627_
timestamp 1676037725
transform 1 0 15364 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1628_
timestamp 1676037725
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1629_
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1630_
timestamp 1676037725
transform 1 0 20516 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1631_
timestamp 1676037725
transform 1 0 17020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1633_
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1635_
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1636_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1637_
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1638_
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1639_
timestamp 1676037725
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1640_
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1676037725
transform 1 0 16836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1642_
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1643_
timestamp 1676037725
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1644_
timestamp 1676037725
transform 1 0 14444 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1676037725
transform 1 0 13524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1646_
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1676037725
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1648_
timestamp 1676037725
transform 1 0 7636 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1650_
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1676037725
transform 1 0 26312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1652_
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1676037725
transform 1 0 27140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1654_
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1655_
timestamp 1676037725
transform 1 0 25668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1656_
timestamp 1676037725
transform 1 0 6992 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1657_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1658_
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1676037725
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1660_
timestamp 1676037725
transform 1 0 12144 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1662_
timestamp 1676037725
transform 1 0 12328 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1676037725
transform 1 0 11684 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1664_
timestamp 1676037725
transform 1 0 15180 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1665_
timestamp 1676037725
transform 1 0 16100 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1666_
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1667_
timestamp 1676037725
transform 1 0 18032 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1671_
timestamp 1676037725
transform 1 0 20792 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1673_
timestamp 1676037725
transform 1 0 20700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1675_
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1677_
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1676037725
transform 1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1679_
timestamp 1676037725
transform 1 0 22356 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1676037725
transform 1 0 23000 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1681_
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1676037725
transform 1 0 23368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1683_
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1685_
timestamp 1676037725
transform 1 0 23552 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1688_
timestamp 1676037725
transform 1 0 20884 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1690_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1676037725
transform 1 0 22080 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1692_
timestamp 1676037725
transform 1 0 23460 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1693_
timestamp 1676037725
transform 1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1694_
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1696_
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1697_
timestamp 1676037725
transform 1 0 23460 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1698_
timestamp 1676037725
transform 1 0 22816 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1700_
timestamp 1676037725
transform 1 0 27876 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1676037725
transform 1 0 27324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1702_
timestamp 1676037725
transform 1 0 27416 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1703_
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1704_
timestamp 1676037725
transform 1 0 27600 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1705_
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1706_
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1708_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1709_
timestamp 1676037725
transform 1 0 22356 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1711_
timestamp 1676037725
transform 1 0 23092 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1676037725
transform 1 0 23368 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1713_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1715_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1716_
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1717_
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1719_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1720_
timestamp 1676037725
transform 1 0 25484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1721_
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1723_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1676037725
transform 1 0 23092 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1725_
timestamp 1676037725
transform 1 0 23092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1676037725
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1727_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1676037725
transform 1 0 26128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1729_
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1730_
timestamp 1676037725
transform 1 0 23552 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1676037725
transform 1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1732_
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1733_
timestamp 1676037725
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1734_
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1735_
timestamp 1676037725
transform 1 0 21252 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1736_
timestamp 1676037725
transform 1 0 20976 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1676037725
transform 1 0 23828 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1738_
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1739_
timestamp 1676037725
transform 1 0 21160 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1740_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1741_
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1742_
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1743_
timestamp 1676037725
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1744_
timestamp 1676037725
transform 1 0 19596 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1745_
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1746_
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1747_
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1748_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1750_
timestamp 1676037725
transform 1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1676037725
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1752_
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1676037725
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1754_
timestamp 1676037725
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1676037725
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1756_
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1757_
timestamp 1676037725
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1758_
timestamp 1676037725
transform 1 0 8740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1759_
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1760_
timestamp 1676037725
transform 1 0 2116 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1761_
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1762_
timestamp 1676037725
transform 1 0 5612 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1763_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1764_
timestamp 1676037725
transform 1 0 3956 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1765_
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _1766_
timestamp 1676037725
transform 1 0 4508 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1767_
timestamp 1676037725
transform 1 0 1656 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1768_
timestamp 1676037725
transform 1 0 4784 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1769_
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _1770_
timestamp 1676037725
transform 1 0 2392 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1771_
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1772_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1773_
timestamp 1676037725
transform 1 0 1748 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1774_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _1775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1776_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1777_
timestamp 1676037725
transform 1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1778_
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1779_
timestamp 1676037725
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1780_
timestamp 1676037725
transform 1 0 5612 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1781_
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1782_
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1784_
timestamp 1676037725
transform 1 0 12696 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1785_
timestamp 1676037725
transform 1 0 5336 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1786_
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1787_
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1788_
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1789_
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1790_
timestamp 1676037725
transform 1 0 8096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1792_
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1793_
timestamp 1676037725
transform 1 0 8004 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1794_
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1795_
timestamp 1676037725
transform 1 0 6256 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1796_
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1797_
timestamp 1676037725
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1798_
timestamp 1676037725
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1799_
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1800_
timestamp 1676037725
transform 1 0 4508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1801_
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1802_
timestamp 1676037725
transform 1 0 4048 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1676037725
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1804_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1805_
timestamp 1676037725
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1806_
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1807_
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1808_
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1809_
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1810_
timestamp 1676037725
transform 1 0 6164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1676037725
transform 1 0 9108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1676037725
transform 1 0 9752 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1676037725
transform 1 0 6808 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1676037725
transform 1 0 4140 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1676037725
transform 1 0 6992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1676037725
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1676037725
transform 1 0 13432 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1676037725
transform 1 0 22172 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1676037725
transform 1 0 26772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1676037725
transform 1 0 26772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1676037725
transform 1 0 20516 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1676037725
transform 1 0 23184 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1676037725
transform 1 0 21988 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1676037725
transform 1 0 26956 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1676037725
transform 1 0 23828 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1676037725
transform 1 0 16468 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1676037725
transform 1 0 17480 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1676037725
transform 1 0 21528 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1676037725
transform 1 0 19596 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1676037725
transform 1 0 11868 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1676037725
transform 1 0 12144 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1676037725
transform 1 0 16100 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1676037725
transform 1 0 13340 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1676037725
transform 1 0 9752 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1676037725
transform 1 0 10672 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1676037725
transform 1 0 13064 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1676037725
transform 1 0 12696 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1676037725
transform 1 0 14996 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1676037725
transform 1 0 16468 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1676037725
transform 1 0 9108 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1676037725
transform 1 0 14904 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1676037725
transform 1 0 17480 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1676037725
transform 1 0 17296 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1676037725
transform 1 0 19320 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1676037725
transform 1 0 17112 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1676037725
transform 1 0 14904 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1676037725
transform 1 0 21804 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1676037725
transform 1 0 19504 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1676037725
transform 1 0 21344 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1676037725
transform 1 0 20056 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1676037725
transform 1 0 22264 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1676037725
transform 1 0 25208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1676037725
transform 1 0 26036 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1676037725
transform 1 0 25208 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1676037725
transform 1 0 25208 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1676037725
transform 1 0 26404 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1676037725
transform 1 0 26864 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1676037725
transform 1 0 26956 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1676037725
transform 1 0 26404 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1676037725
transform 1 0 25208 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1676037725
transform 1 0 22632 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1676037725
transform 1 0 19780 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1676037725
transform 1 0 14904 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1676037725
transform 1 0 12420 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1676037725
transform 1 0 11684 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1676037725
transform 1 0 9568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1676037725
transform 1 0 9752 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1676037725
transform 1 0 7912 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1676037725
transform 1 0 24932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1676037725
transform 1 0 25208 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1676037725
transform 1 0 21712 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1676037725
transform 1 0 24564 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1676037725
transform 1 0 25116 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1676037725
transform 1 0 22632 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1676037725
transform 1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1676037725
transform 1 0 11684 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1676037725
transform 1 0 9752 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1676037725
transform 1 0 18216 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1676037725
transform 1 0 14352 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1676037725
transform 1 0 16836 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1676037725
transform 1 0 23828 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1676037725
transform 1 0 21988 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1676037725
transform 1 0 20148 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1676037725
transform 1 0 20516 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1676037725
transform 1 0 19412 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1676037725
transform 1 0 18676 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1676037725
transform 1 0 3956 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1676037725
transform 1 0 2116 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1676037725
transform 1 0 2944 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1676037725
transform 1 0 9568 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1676037725
transform 1 0 13248 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1676037725
transform 1 0 17480 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1676037725
transform 1 0 21988 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1676037725
transform 1 0 24564 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1676037725
transform 1 0 26956 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1676037725
transform 1 0 26404 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1676037725
transform 1 0 23644 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1676037725
transform 1 0 26956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1676037725
transform 1 0 26036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1676037725
transform 1 0 23644 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1676037725
transform 1 0 25208 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1676037725
transform 1 0 26404 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1981_
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1982_
timestamp 1676037725
transform 1 0 25760 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1983_
timestamp 1676037725
transform 1 0 26680 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1676037725
transform 1 0 26220 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1676037725
transform 1 0 24748 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1986_
timestamp 1676037725
transform 1 0 25208 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1987_
timestamp 1676037725
transform 1 0 26956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1988_
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1989_
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1990_
timestamp 1676037725
transform 1 0 25116 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1991_
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1992_
timestamp 1676037725
transform 1 0 24380 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1993_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1994_
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1995_
timestamp 1676037725
transform 1 0 24748 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1996_
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1997_
timestamp 1676037725
transform 1 0 14352 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1998_
timestamp 1676037725
transform 1 0 11868 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1999_
timestamp 1676037725
transform 1 0 9108 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2000_
timestamp 1676037725
transform 1 0 6624 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2001_
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2002_
timestamp 1676037725
transform 1 0 14168 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2003_
timestamp 1676037725
transform 1 0 2024 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2005_
timestamp 1676037725
transform 1 0 1932 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2006_
timestamp 1676037725
transform 1 0 2576 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2007_
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2008_
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2009_
timestamp 1676037725
transform 1 0 1748 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2010_
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2011_
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2012_
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2013_
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2014_
timestamp 1676037725
transform 1 0 1656 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2015_
timestamp 1676037725
transform 1 0 1748 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2016_
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2017_
timestamp 1676037725
transform 1 0 1748 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2018_
timestamp 1676037725
transform 1 0 1748 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2019_
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2020_
timestamp 1676037725
transform 1 0 3680 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1676037725
transform 1 0 1748 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1676037725
transform 1 0 1564 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2023_
timestamp 1676037725
transform 1 0 1656 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_in[0]
timestamp 1676037725
transform 1 0 2852 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net57
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 2852 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0380_
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_io_in[0]
timestamp 1676037725
transform 1 0 2576 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net57
timestamp 1676037725
transform 1 0 2576 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 10396 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 1564 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0380_
timestamp 1676037725
transform 1 0 1656 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_io_in[0]
timestamp 1676037725
transform 1 0 2576 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net57
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 5244 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout9
timestamp 1676037725
transform 1 0 8096 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout10
timestamp 1676037725
transform 1 0 11684 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout11
timestamp 1676037725
transform 1 0 12420 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout12
timestamp 1676037725
transform 1 0 8280 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout13
timestamp 1676037725
transform 1 0 7544 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1676037725
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1676037725
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1676037725
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout19
timestamp 1676037725
transform 1 0 15732 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1676037725
transform 1 0 23276 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout21
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout23
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1676037725
transform 1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1676037725
transform 1 0 11684 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1676037725
transform 1 0 9752 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1676037725
transform 1 0 22724 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout31
timestamp 1676037725
transform 1 0 23368 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1676037725
transform 1 0 14260 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout33
timestamp 1676037725
transform 1 0 18768 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout37
timestamp 1676037725
transform 1 0 15824 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[0\].cap_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27784 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[0\].cap
timestamp 1676037725
transform 1 0 26404 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[1\].cap
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[1\].cap_46
timestamp 1676037725
transform 1 0 23828 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[2\].cap_47
timestamp 1676037725
transform 1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[2\].cap
timestamp 1676037725
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[3\].cap_48
timestamp 1676037725
transform 1 0 22724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[3\].cap
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[4\].cap
timestamp 1676037725
transform 1 0 23828 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[4\].cap_49
timestamp 1676037725
transform 1 0 26496 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[5\].cap
timestamp 1676037725
transform 1 0 25944 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[5\].cap_50
timestamp 1676037725
transform 1 0 23368 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[6\].cap_51
timestamp 1676037725
transform 1 0 27140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[6\].cap
timestamp 1676037725
transform 1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[7\].cap
timestamp 1676037725
transform 1 0 24656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[7\].cap_52
timestamp 1676037725
transform 1 0 24104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[8\].cap_53
timestamp 1676037725
transform 1 0 27048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[8\].cap
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[9\].cap
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[9\].cap_54
timestamp 1676037725
transform 1 0 22080 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[10\].cap
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[10\].cap_40
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[11\].cap
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[11\].cap_41
timestamp 1676037725
transform 1 0 25760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[12\].cap
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[12\].cap_42
timestamp 1676037725
transform 1 0 23276 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[13\].cap_43
timestamp 1676037725
transform 1 0 25208 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[13\].cap
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[14\].cap_44
timestamp 1676037725
transform 1 0 24564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[14\].cap
timestamp 1676037725
transform 1 0 27784 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[15\].cap
timestamp 1676037725
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[15\].cap_45
timestamp 1676037725
transform 1 0 25208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 5244 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 4600 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 7360 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 4784 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 9016 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 3956 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 8740 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 4784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 8188 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 6900 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 6532 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 8188 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 9568 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1676037725
transform 1 0 9936 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1676037725
transform 1 0 6532 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1676037725
transform 1 0 6624 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1676037725
transform 1 0 12236 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1676037725
transform 1 0 5612 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1676037725
transform 1 0 7360 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 5704 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 6532 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 13156 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 16100 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 13156 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 1656 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 10672 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1676037725
transform 1 0 5704 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1676037725
transform 1 0 4048 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1676037725
transform 1 0 11592 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1676037725
transform 1 0 13248 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1676037725
transform 1 0 16928 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1676037725
transform 1 0 9844 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1676037725
transform 1 0 3036 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1676037725
transform 1 0 9568 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1676037725
transform 1 0 15364 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1676037725
transform 1 0 5612 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1676037725
transform 1 0 12328 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1676037725
transform 1 0 18308 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1676037725
transform 1 0 13156 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1676037725
transform 1 0 5612 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1676037725
transform 1 0 13156 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1676037725
transform 1 0 5704 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1676037725
transform 1 0 12328 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1676037725
transform 1 0 4048 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1676037725
transform 1 0 12328 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1676037725
transform 1 0 6532 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1676037725
transform 1 0 11500 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd_56
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 8924 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].vref_55
timestamp 1676037725
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 17112 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dcdc
timestamp 1676037725
transform 1 0 15456 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  temp1.inv1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_2
timestamp 1676037725
transform 1 0 27140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_3
timestamp 1676037725
transform 1 0 27140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_4
timestamp 1676037725
transform 1 0 27784 0 -1 28288
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 1640 400 1760 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 3680 400 3800 0 FreeSans 480 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 0 5720 400 5840 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal3 s 0 7760 400 7880 0 FreeSans 480 0 0 0 io_in[3]
port 3 nsew signal input
flabel metal3 s 0 9800 400 9920 0 FreeSans 480 0 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 0 11840 400 11960 0 FreeSans 480 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal3 s 0 13880 400 14000 0 FreeSans 480 0 0 0 io_in[6]
port 6 nsew signal input
flabel metal3 s 0 15920 400 16040 0 FreeSans 480 0 0 0 io_in[7]
port 7 nsew signal input
flabel metal3 s 0 17960 400 18080 0 FreeSans 480 0 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal3 s 0 20000 400 20120 0 FreeSans 480 0 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal3 s 0 22040 400 22160 0 FreeSans 480 0 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal3 s 0 24080 400 24200 0 FreeSans 480 0 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal3 s 0 26120 400 26240 0 FreeSans 480 0 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal3 s 0 28160 400 28280 0 FreeSans 480 0 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal3 s 0 30200 400 30320 0 FreeSans 480 0 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal3 s 0 32240 400 32360 0 FreeSans 480 0 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 4417 1040 4737 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 11363 1040 11683 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 18309 1040 18629 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 25255 1040 25575 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7890 1040 8210 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 14836 1040 15156 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 21782 1040 22102 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 28728 1040 29048 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 14996 32096 14996 32096 0 vccd1
rlabel via1 15076 32640 15076 32640 0 vssd1
rlabel metal1 6389 2346 6389 2346 0 _0000_
rlabel metal2 8418 7174 8418 7174 0 _0001_
rlabel metal2 10442 8262 10442 8262 0 _0002_
rlabel metal1 6798 4114 6798 4114 0 _0003_
rlabel metal2 5934 986 5934 986 0 _0004_
rlabel metal1 6486 2074 6486 2074 0 _0005_
rlabel metal1 10948 16218 10948 16218 0 _0006_
rlabel metal1 8004 26554 8004 26554 0 _0007_
rlabel metal2 13570 24276 13570 24276 0 _0008_
rlabel metal1 16780 18258 16780 18258 0 _0009_
rlabel metal1 15640 17306 15640 17306 0 _0010_
rlabel metal1 16422 16966 16422 16966 0 _0011_
rlabel metal1 23966 20026 23966 20026 0 _0012_
rlabel metal1 26480 16490 26480 16490 0 _0013_
rlabel via1 27089 15470 27089 15470 0 _0014_
rlabel metal1 23230 17816 23230 17816 0 _0015_
rlabel metal2 22586 19176 22586 19176 0 _0016_
rlabel via2 19458 22219 19458 22219 0 _0017_
rlabel metal1 18216 21862 18216 21862 0 _0018_
rlabel metal1 18666 14994 18666 14994 0 _0019_
rlabel metal2 16054 15079 16054 15079 0 _0020_
rlabel metal2 22586 23426 22586 23426 0 _0021_
rlabel metal1 21712 23834 21712 23834 0 _0022_
rlabel metal1 19136 24378 19136 24378 0 _0023_
rlabel metal1 20332 23834 20332 23834 0 _0024_
rlabel metal1 23736 25466 23736 25466 0 _0025_
rlabel metal1 21206 24616 21206 24616 0 _0026_
rlabel metal1 20608 25466 20608 25466 0 _0027_
rlabel metal2 20470 25075 20470 25075 0 _0028_
rlabel metal2 13846 24616 13846 24616 0 _0029_
rlabel metal2 17158 25364 17158 25364 0 _0030_
rlabel metal1 21206 31790 21206 31790 0 _0031_
rlabel metal1 20424 27574 20424 27574 0 _0032_
rlabel metal2 14122 28900 14122 28900 0 _0033_
rlabel metal1 15210 24106 15210 24106 0 _0034_
rlabel metal1 12134 15402 12134 15402 0 _0035_
rlabel metal1 11628 11798 11628 11798 0 _0036_
rlabel metal2 10902 10608 10902 10608 0 _0037_
rlabel metal3 12305 9588 12305 9588 0 _0038_
rlabel metal1 12788 15130 12788 15130 0 _0039_
rlabel metal2 13018 21318 13018 21318 0 _0040_
rlabel metal1 7682 21114 7682 21114 0 _0041_
rlabel metal2 21758 31042 21758 31042 0 _0042_
rlabel metal2 14674 30481 14674 30481 0 _0043_
rlabel metal2 10442 32470 10442 32470 0 _0044_
rlabel metal2 18722 28781 18722 28781 0 _0045_
rlabel metal2 13754 29971 13754 29971 0 _0046_
rlabel metal2 12650 27200 12650 27200 0 _0047_
rlabel metal1 17388 27098 17388 27098 0 _0048_
rlabel metal2 9430 31263 9430 31263 0 _0049_
rlabel metal1 21482 31314 21482 31314 0 _0050_
rlabel metal1 12742 32232 12742 32232 0 _0051_
rlabel metal1 17188 29206 17188 29206 0 _0052_
rlabel metal1 19632 29614 19632 29614 0 _0053_
rlabel metal2 17112 32980 17112 32980 0 _0054_
rlabel metal2 16928 32538 16928 32538 0 _0055_
rlabel metal2 17112 32436 17112 32436 0 _0056_
rlabel metal2 14674 32572 14674 32572 0 _0057_
rlabel metal2 21942 29818 21942 29818 0 _0058_
rlabel metal2 21482 28934 21482 28934 0 _0059_
rlabel metal2 20746 30498 20746 30498 0 _0060_
rlabel metal1 21564 30702 21564 30702 0 _0061_
rlabel metal1 22172 29274 22172 29274 0 _0062_
rlabel metal1 20746 27336 20746 27336 0 _0063_
rlabel metal2 19458 27574 19458 27574 0 _0064_
rlabel metal1 19872 26010 19872 26010 0 _0065_
rlabel metal1 24124 21930 24124 21930 0 _0066_
rlabel metal1 22678 18088 22678 18088 0 _0067_
rlabel metal1 22724 21114 22724 21114 0 _0068_
rlabel metal2 24518 27064 24518 27064 0 _0069_
rlabel metal1 24380 24650 24380 24650 0 _0070_
rlabel metal2 22402 22780 22402 22780 0 _0071_
rlabel metal1 21574 25466 21574 25466 0 _0072_
rlabel metal2 25070 25432 25070 25432 0 _0073_
rlabel metal1 24610 21658 24610 21658 0 _0074_
rlabel metal1 25208 22950 25208 22950 0 _0075_
rlabel metal2 21022 25109 21022 25109 0 _0076_
rlabel metal1 22770 20570 22770 20570 0 _0077_
rlabel metal1 20930 21862 20930 21862 0 _0078_
rlabel metal1 26624 17646 26624 17646 0 _0079_
rlabel via1 22494 18139 22494 18139 0 _0080_
rlabel metal1 22218 21420 22218 21420 0 _0081_
rlabel metal1 20286 25772 20286 25772 0 _0082_
rlabel metal1 19182 25670 19182 25670 0 _0083_
rlabel metal1 20378 26758 20378 26758 0 _0084_
rlabel metal1 17158 31450 17158 31450 0 _0085_
rlabel metal1 18906 31790 18906 31790 0 _0086_
rlabel metal1 19120 26282 19120 26282 0 _0087_
rlabel metal1 15226 23188 15226 23188 0 _0088_
rlabel metal1 9292 24922 9292 24922 0 _0089_
rlabel via1 12737 25874 12737 25874 0 _0090_
rlabel metal3 18124 28764 18124 28764 0 _0091_
rlabel metal1 20746 26758 20746 26758 0 _0092_
rlabel metal1 10150 27370 10150 27370 0 _0093_
rlabel viali 10253 19754 10253 19754 0 _0094_
rlabel metal1 10672 13498 10672 13498 0 _0095_
rlabel metal1 11898 8534 11898 8534 0 _0096_
rlabel via1 10069 6358 10069 6358 0 _0097_
rlabel metal1 7942 2006 7942 2006 0 _0098_
rlabel metal1 10616 3502 10616 3502 0 _0099_
rlabel via1 12829 12818 12829 12818 0 _0100_
rlabel metal2 13478 10557 13478 10557 0 _0101_
rlabel metal1 18446 12750 18446 12750 0 _0102_
rlabel metal2 20746 15011 20746 15011 0 _0103_
rlabel via1 25249 8534 25249 8534 0 _0104_
rlabel metal1 22034 8568 22034 8568 0 _0105_
rlabel metal1 21104 6766 21104 6766 0 _0106_
rlabel metal2 17802 10744 17802 10744 0 _0107_
rlabel metal1 27084 11118 27084 11118 0 _0108_
rlabel metal2 22770 8194 22770 8194 0 _0109_
rlabel metal1 25474 6290 25474 6290 0 _0110_
rlabel via1 24881 5610 24881 5610 0 _0111_
rlabel metal1 19274 5338 19274 5338 0 _0112_
rlabel metal1 21643 7174 21643 7174 0 _0113_
rlabel metal1 23138 8296 23138 8296 0 _0114_
rlabel metal1 26756 9962 26756 9962 0 _0115_
rlabel metal1 24104 8058 24104 8058 0 _0116_
rlabel metal1 22586 8942 22586 8942 0 _0117_
rlabel metal1 20010 5304 20010 5304 0 _0118_
rlabel metal1 15768 3502 15768 3502 0 _0119_
rlabel metal1 11438 1258 11438 1258 0 _0120_
rlabel metal1 9149 3026 9149 3026 0 _0121_
rlabel metal2 10994 1462 10994 1462 0 _0122_
rlabel metal1 13577 3094 13577 3094 0 _0123_
rlabel metal1 14858 2618 14858 2618 0 _0124_
rlabel metal1 14715 4182 14715 4182 0 _0125_
rlabel metal1 16820 2006 16820 2006 0 _0126_
rlabel metal1 14536 2550 14536 2550 0 _0127_
rlabel metal2 21574 2023 21574 2023 0 _0128_
rlabel metal1 20562 1904 20562 1904 0 _0129_
rlabel metal1 18860 3706 18860 3706 0 _0130_
rlabel metal1 17572 5338 17572 5338 0 _0131_
rlabel metal1 22110 2346 22110 2346 0 _0132_
rlabel metal1 17618 2312 17618 2312 0 _0133_
rlabel metal1 18982 1258 18982 1258 0 _0134_
rlabel metal1 18246 2006 18246 2006 0 _0135_
rlabel metal1 13616 1190 13616 1190 0 _0136_
rlabel metal1 11628 2414 11628 2414 0 _0137_
rlabel metal1 5469 2006 5469 2006 0 _0138_
rlabel metal2 26358 2023 26358 2023 0 _0139_
rlabel metal2 27186 1020 27186 1020 0 _0140_
rlabel metal2 25714 2159 25714 2159 0 _0141_
rlabel metal1 11730 2312 11730 2312 0 _0142_
rlabel metal1 13048 2006 13048 2006 0 _0143_
rlabel metal1 12282 3060 12282 3060 0 _0144_
rlabel metal2 15134 1462 15134 1462 0 _0145_
rlabel metal1 19826 1292 19826 1292 0 _0146_
rlabel via1 24881 1326 24881 1326 0 _0147_
rlabel metal1 25330 4522 25330 4522 0 _0148_
rlabel metal1 23782 5304 23782 5304 0 _0149_
rlabel metal1 27176 3502 27176 3502 0 _0150_
rlabel metal1 26624 6766 26624 6766 0 _0151_
rlabel metal1 25571 9554 25571 9554 0 _0152_
rlabel via1 25157 11050 25157 11050 0 _0153_
rlabel metal1 23920 9418 23920 9418 0 _0154_
rlabel metal2 22034 11458 22034 11458 0 _0155_
rlabel metal1 24150 14042 24150 14042 0 _0156_
rlabel metal1 24380 19958 24380 19958 0 _0157_
rlabel via1 23961 21590 23961 21590 0 _0158_
rlabel metal2 26266 19414 26266 19414 0 _0159_
rlabel metal1 25238 18666 25238 18666 0 _0160_
rlabel metal1 24196 23290 24196 23290 0 _0161_
rlabel metal1 25019 20910 25019 20910 0 _0162_
rlabel metal1 25939 16150 25939 16150 0 _0163_
rlabel metal2 28106 14722 28106 14722 0 _0164_
rlabel metal1 27738 16218 27738 16218 0 _0165_
rlabel via1 26721 13294 26721 13294 0 _0166_
rlabel metal1 25928 12138 25928 12138 0 _0167_
rlabel metal1 23460 12682 23460 12682 0 _0168_
rlabel metal2 28106 13090 28106 13090 0 _0169_
rlabel metal1 23823 11050 23823 11050 0 _0170_
rlabel metal1 25330 7786 25330 7786 0 _0171_
rlabel metal1 26900 8942 26900 8942 0 _0172_
rlabel metal1 25560 14314 25560 14314 0 _0173_
rlabel metal1 24012 15130 24012 15130 0 _0174_
rlabel via1 25525 13974 25525 13974 0 _0175_
rlabel metal1 26710 5610 26710 5610 0 _0176_
rlabel metal1 26900 2414 26900 2414 0 _0177_
rlabel metal1 20424 3162 20424 3162 0 _0178_
rlabel metal1 23138 1258 23138 1258 0 _0179_
rlabel metal1 23874 1224 23874 1224 0 _0180_
rlabel metal1 21942 1734 21942 1734 0 _0181_
rlabel metal2 19458 2601 19458 2601 0 _0182_
rlabel metal1 24927 2346 24927 2346 0 _0183_
rlabel via1 23414 6069 23414 6069 0 _0184_
rlabel metal1 20608 7514 20608 7514 0 _0185_
rlabel metal1 14152 5270 14152 5270 0 _0186_
rlabel metal1 11530 5270 11530 5270 0 _0187_
rlabel metal1 8586 4522 8586 4522 0 _0188_
rlabel via2 8234 1275 8234 1275 0 _0189_
rlabel metal1 7130 4794 7130 4794 0 _0190_
rlabel metal1 13445 7378 13445 7378 0 _0191_
rlabel metal1 2387 27370 2387 27370 0 _0192_
rlabel metal1 3491 28050 3491 28050 0 _0193_
rlabel metal1 2152 25262 2152 25262 0 _0194_
rlabel metal1 3491 24786 3491 24786 0 _0195_
rlabel metal2 1886 25058 1886 25058 0 _0196_
rlabel metal1 2244 24174 2244 24174 0 _0197_
rlabel metal1 1968 28526 1968 28526 0 _0198_
rlabel metal1 1334 19686 1334 19686 0 _0199_
rlabel metal3 1127 9588 1127 9588 0 _0200_
rlabel metal1 2847 4590 2847 4590 0 _0201_
rlabel metal1 1594 8534 1594 8534 0 _0202_
rlabel metal3 2507 8228 2507 8228 0 _0203_
rlabel metal1 1334 7310 1334 7310 0 _0204_
rlabel metal3 1357 2516 1357 2516 0 _0205_
rlabel metal1 1968 4114 1968 4114 0 _0206_
rlabel metal1 4002 3570 4002 3570 0 _0207_
rlabel metal1 4554 3978 4554 3978 0 _0208_
rlabel metal1 3956 5338 3956 5338 0 _0209_
rlabel metal2 5474 4318 5474 4318 0 _0210_
rlabel metal1 2341 1326 2341 1326 0 _0211_
rlabel metal1 2364 13294 2364 13294 0 _0212_
rlabel metal2 9706 19924 9706 19924 0 _0213_
rlabel metal1 8970 20026 8970 20026 0 _0214_
rlabel metal3 13708 24004 13708 24004 0 _0215_
rlabel metal1 7498 31790 7498 31790 0 _0216_
rlabel metal1 15134 28696 15134 28696 0 _0217_
rlabel metal1 8096 31926 8096 31926 0 _0218_
rlabel metal3 17020 28288 17020 28288 0 _0219_
rlabel metal2 7314 25517 7314 25517 0 _0220_
rlabel metal1 11132 26010 11132 26010 0 _0221_
rlabel metal1 19090 29206 19090 29206 0 _0222_
rlabel metal1 15870 25330 15870 25330 0 _0223_
rlabel via2 7682 30141 7682 30141 0 _0224_
rlabel metal2 10074 32504 10074 32504 0 _0225_
rlabel metal1 13386 32368 13386 32368 0 _0226_
rlabel metal1 15364 27098 15364 27098 0 _0227_
rlabel metal1 15410 26826 15410 26826 0 _0228_
rlabel metal1 14352 28186 14352 28186 0 _0229_
rlabel metal2 13754 32606 13754 32606 0 _0230_
rlabel metal2 12834 32878 12834 32878 0 _0231_
rlabel metal1 14904 30158 14904 30158 0 _0232_
rlabel metal1 15134 27574 15134 27574 0 _0233_
rlabel metal2 21298 26962 21298 26962 0 _0234_
rlabel metal1 20240 29274 20240 29274 0 _0235_
rlabel metal1 16606 33082 16606 33082 0 _0236_
rlabel metal2 19918 19856 19918 19856 0 _0237_
rlabel metal1 20470 28424 20470 28424 0 _0238_
rlabel metal1 19918 26554 19918 26554 0 _0239_
rlabel metal1 18377 27030 18377 27030 0 _0240_
rlabel metal2 19826 25670 19826 25670 0 _0241_
rlabel metal2 18906 22304 18906 22304 0 _0242_
rlabel metal1 22494 18224 22494 18224 0 _0243_
rlabel metal2 22402 20196 22402 20196 0 _0244_
rlabel metal1 22954 21862 22954 21862 0 _0245_
rlabel metal1 20194 19754 20194 19754 0 _0246_
rlabel metal2 23046 24208 23046 24208 0 _0247_
rlabel metal1 21436 21658 21436 21658 0 _0248_
rlabel metal1 21252 25262 21252 25262 0 _0249_
rlabel metal2 20562 24276 20562 24276 0 _0250_
rlabel metal2 21758 21318 21758 21318 0 _0251_
rlabel metal1 22678 20978 22678 20978 0 _0252_
rlabel metal2 21390 24412 21390 24412 0 _0253_
rlabel metal1 21160 20434 21160 20434 0 _0254_
rlabel metal2 19734 21828 19734 21828 0 _0255_
rlabel metal1 22632 19482 22632 19482 0 _0256_
rlabel metal2 19826 18054 19826 18054 0 _0257_
rlabel metal1 21252 20026 21252 20026 0 _0258_
rlabel metal1 20010 24922 20010 24922 0 _0259_
rlabel via2 7958 9571 7958 9571 0 _0260_
rlabel metal2 17894 25670 17894 25670 0 _0261_
rlabel metal1 19159 26894 19159 26894 0 _0262_
rlabel metal1 16376 27098 16376 27098 0 _0263_
rlabel metal1 16560 32402 16560 32402 0 _0264_
rlabel metal1 14490 24310 14490 24310 0 _0265_
rlabel metal1 15640 11118 15640 11118 0 _0266_
rlabel metal1 15088 23086 15088 23086 0 _0267_
rlabel metal1 10764 21046 10764 21046 0 _0268_
rlabel metal1 12926 21488 12926 21488 0 _0269_
rlabel metal3 17204 24208 17204 24208 0 _0270_
rlabel metal2 20746 26299 20746 26299 0 _0271_
rlabel metal1 7682 22406 7682 22406 0 _0272_
rlabel metal2 8326 20434 8326 20434 0 _0273_
rlabel metal1 10442 13294 10442 13294 0 _0274_
rlabel metal1 9568 10642 9568 10642 0 _0275_
rlabel metal1 8464 9690 8464 9690 0 _0276_
rlabel metal1 7728 5678 7728 5678 0 _0277_
rlabel metal2 8878 4556 8878 4556 0 _0278_
rlabel metal2 10810 10812 10810 10812 0 _0279_
rlabel metal1 9338 12240 9338 12240 0 _0280_
rlabel metal1 14674 12818 14674 12818 0 _0281_
rlabel metal1 18262 15028 18262 15028 0 _0282_
rlabel metal2 19366 9010 19366 9010 0 _0283_
rlabel metal2 22310 10880 22310 10880 0 _0284_
rlabel metal1 20907 8398 20907 8398 0 _0285_
rlabel metal1 20378 8500 20378 8500 0 _0286_
rlabel metal1 18446 11118 18446 11118 0 _0287_
rlabel metal1 19872 10982 19872 10982 0 _0288_
rlabel metal1 22080 9622 22080 9622 0 _0289_
rlabel metal1 11500 1326 11500 1326 0 _0290_
rlabel metal1 21758 8942 21758 8942 0 _0291_
rlabel metal1 20654 7888 20654 7888 0 _0292_
rlabel metal2 18906 6460 18906 6460 0 _0293_
rlabel metal2 19918 7140 19918 7140 0 _0294_
rlabel metal1 20838 8466 20838 8466 0 _0295_
rlabel metal2 22862 9350 22862 9350 0 _0296_
rlabel metal1 22770 10472 22770 10472 0 _0297_
rlabel metal2 21298 9146 21298 9146 0 _0298_
rlabel metal1 10396 1326 10396 1326 0 _0299_
rlabel metal2 20194 5372 20194 5372 0 _0300_
rlabel metal1 14812 5202 14812 5202 0 _0301_
rlabel metal1 11086 3060 11086 3060 0 _0302_
rlabel metal1 10948 1326 10948 1326 0 _0303_
rlabel metal2 9982 1054 9982 1054 0 _0304_
rlabel metal2 12190 3740 12190 3740 0 _0305_
rlabel metal1 14582 2414 14582 2414 0 _0306_
rlabel metal1 14950 4590 14950 4590 0 _0307_
rlabel metal2 12926 3978 12926 3978 0 _0308_
rlabel metal2 13754 2890 13754 2890 0 _0309_
rlabel metal1 15870 1394 15870 1394 0 _0310_
rlabel metal1 20838 1938 20838 1938 0 _0311_
rlabel metal1 18400 3502 18400 3502 0 _0312_
rlabel metal2 17066 5372 17066 5372 0 _0313_
rlabel metal1 19642 4624 19642 4624 0 _0314_
rlabel metal1 17526 3910 17526 3910 0 _0315_
rlabel metal1 4370 2550 4370 2550 0 _0316_
rlabel metal1 17480 3366 17480 3366 0 _0317_
rlabel metal1 14996 3366 14996 3366 0 _0318_
rlabel metal1 13754 1258 13754 1258 0 _0319_
rlabel metal2 11178 4998 11178 4998 0 _0320_
rlabel metal1 7682 3638 7682 3638 0 _0321_
rlabel metal2 4830 2329 4830 2329 0 _0322_
rlabel metal2 27370 986 27370 986 0 _0323_
rlabel metal1 25898 2006 25898 2006 0 _0324_
rlabel metal1 9108 1734 9108 1734 0 _0325_
rlabel metal1 10534 3026 10534 3026 0 _0326_
rlabel metal1 12650 4080 12650 4080 0 _0327_
rlabel metal1 11914 1904 11914 1904 0 _0328_
rlabel metal1 16330 1904 16330 1904 0 _0329_
rlabel metal1 21528 10098 21528 10098 0 _0330_
rlabel metal2 19550 5916 19550 5916 0 _0331_
rlabel metal1 24794 4624 24794 4624 0 _0332_
rlabel metal1 21689 5134 21689 5134 0 _0333_
rlabel metal2 24242 6222 24242 6222 0 _0334_
rlabel metal1 23414 7378 23414 7378 0 _0335_
rlabel metal3 24702 9724 24702 9724 0 _0336_
rlabel metal2 23230 11900 23230 11900 0 _0337_
rlabel metal2 23598 10914 23598 10914 0 _0338_
rlabel metal1 23138 10166 23138 10166 0 _0339_
rlabel metal1 24150 13498 24150 13498 0 _0340_
rlabel metal2 21942 16796 21942 16796 0 _0341_
rlabel metal2 22310 18564 22310 18564 0 _0342_
rlabel metal1 22402 21658 22402 21658 0 _0343_
rlabel metal1 26450 18292 26450 18292 0 _0344_
rlabel metal1 22954 16422 22954 16422 0 _0345_
rlabel metal2 23414 20570 23414 20570 0 _0346_
rlabel metal2 23322 21318 23322 21318 0 _0347_
rlabel metal2 27554 16524 27554 16524 0 _0348_
rlabel metal1 28106 11866 28106 11866 0 _0349_
rlabel metal1 28152 15130 28152 15130 0 _0350_
rlabel metal1 25208 14382 25208 14382 0 _0351_
rlabel metal2 27186 13362 27186 13362 0 _0352_
rlabel metal1 23782 13158 23782 13158 0 _0353_
rlabel metal2 23598 13260 23598 13260 0 _0354_
rlabel metal1 27968 12818 27968 12818 0 _0355_
rlabel metal1 27186 12614 27186 12614 0 _0356_
rlabel metal1 24380 7854 24380 7854 0 _0357_
rlabel metal1 25714 10676 25714 10676 0 _0358_
rlabel metal1 24794 14416 24794 14416 0 _0359_
rlabel metal2 23322 15436 23322 15436 0 _0360_
rlabel metal1 21482 13940 21482 13940 0 _0361_
rlabel metal2 26358 11458 26358 11458 0 _0362_
rlabel metal1 18124 6426 18124 6426 0 _0363_
rlabel metal2 24702 5372 24702 5372 0 _0364_
rlabel metal2 20562 3468 20562 3468 0 _0365_
rlabel metal1 21620 3366 21620 3366 0 _0366_
rlabel metal2 22310 3094 22310 3094 0 _0367_
rlabel metal1 21114 3366 21114 3366 0 _0368_
rlabel metal1 19780 3366 19780 3366 0 _0369_
rlabel viali 21206 4116 21206 4116 0 _0370_
rlabel metal2 20286 6732 20286 6732 0 _0371_
rlabel metal1 20792 6970 20792 6970 0 _0372_
rlabel metal1 17388 6970 17388 6970 0 _0373_
rlabel metal1 8602 7888 8602 7888 0 _0374_
rlabel metal1 7866 6766 7866 6766 0 _0375_
rlabel via2 13754 13923 13754 13923 0 _0376_
rlabel metal1 6348 4590 6348 4590 0 _0377_
rlabel viali 9246 9675 9246 9675 0 _0378_
rlabel metal2 2806 30243 2806 30243 0 _0379_
rlabel via2 3450 25925 3450 25925 0 _0380_
rlabel metal1 2438 25908 2438 25908 0 _0381_
rlabel metal2 4278 27914 4278 27914 0 _0382_
rlabel metal1 1886 28084 1886 28084 0 _0383_
rlabel metal2 4186 26622 4186 26622 0 _0384_
rlabel metal2 1886 24038 1886 24038 0 _0385_
rlabel metal1 2208 26962 2208 26962 0 _0386_
rlabel metal1 2254 30124 2254 30124 0 _0387_
rlabel metal2 1978 20604 1978 20604 0 _0388_
rlabel metal2 6118 20060 6118 20060 0 _0389_
rlabel metal1 4324 13158 4324 13158 0 _0390_
rlabel metal2 1794 11917 1794 11917 0 _0391_
rlabel metal2 1242 8670 1242 8670 0 _0392_
rlabel metal2 12834 18071 12834 18071 0 _0393_
rlabel metal1 5842 18258 5842 18258 0 _0394_
rlabel metal1 6532 16218 6532 16218 0 _0395_
rlabel metal1 7406 16558 7406 16558 0 _0396_
rlabel metal2 7406 14450 7406 14450 0 _0397_
rlabel metal1 7406 12138 7406 12138 0 _0398_
rlabel metal1 7130 11866 7130 11866 0 _0399_
rlabel metal2 5658 11900 5658 11900 0 _0400_
rlabel metal2 5842 8432 5842 8432 0 _0401_
rlabel metal1 5934 3706 5934 3706 0 _0402_
rlabel metal2 13110 8602 13110 8602 0 _0403_
rlabel metal1 4416 4794 4416 4794 0 _0404_
rlabel metal1 5566 3536 5566 3536 0 _0405_
rlabel metal2 6578 5712 6578 5712 0 _0406_
rlabel metal2 18814 4573 18814 4573 0 _0407_
rlabel metal1 6900 14382 6900 14382 0 _0408_
rlabel metal1 6762 10234 6762 10234 0 _0409_
rlabel via2 14674 26197 14674 26197 0 _0410_
rlabel metal1 2024 29478 2024 29478 0 _0411_
rlabel metal1 6026 19856 6026 19856 0 _0412_
rlabel metal1 7958 24786 7958 24786 0 _0413_
rlabel metal1 5842 30158 5842 30158 0 _0414_
rlabel metal1 5244 27506 5244 27506 0 _0415_
rlabel metal4 17940 27336 17940 27336 0 _0416_
rlabel metal1 8464 25670 8464 25670 0 _0417_
rlabel metal1 2300 29546 2300 29546 0 _0418_
rlabel metal1 3404 22610 3404 22610 0 _0419_
rlabel metal1 6854 21930 6854 21930 0 _0420_
rlabel metal1 11086 19278 11086 19278 0 _0421_
rlabel metal2 20746 24497 20746 24497 0 _0422_
rlabel metal1 10994 24922 10994 24922 0 _0423_
rlabel metal2 2714 32096 2714 32096 0 _0424_
rlabel metal1 7130 21658 7130 21658 0 _0425_
rlabel via2 23230 26299 23230 26299 0 _0426_
rlabel metal1 8602 22032 8602 22032 0 _0427_
rlabel metal1 2208 22950 2208 22950 0 _0428_
rlabel metal2 8970 20332 8970 20332 0 _0429_
rlabel metal1 2898 22066 2898 22066 0 _0430_
rlabel via1 5198 17646 5198 17646 0 _0431_
rlabel metal1 5934 19414 5934 19414 0 _0432_
rlabel metal1 1748 20434 1748 20434 0 _0433_
rlabel via2 10810 19261 10810 19261 0 _0434_
rlabel metal1 2622 20264 2622 20264 0 _0435_
rlabel metal1 4002 12954 4002 12954 0 _0436_
rlabel metal2 10810 14654 10810 14654 0 _0437_
rlabel metal1 3450 20842 3450 20842 0 _0438_
rlabel metal2 6210 20468 6210 20468 0 _0439_
rlabel metal1 16008 13158 16008 13158 0 _0440_
rlabel via1 18170 10693 18170 10693 0 _0441_
rlabel metal1 7590 20230 7590 20230 0 _0442_
rlabel metal1 15042 19278 15042 19278 0 _0443_
rlabel via1 19000 17170 19000 17170 0 _0444_
rlabel metal1 13616 10778 13616 10778 0 _0445_
rlabel metal1 7176 18666 7176 18666 0 _0446_
rlabel metal1 7866 17578 7866 17578 0 _0447_
rlabel metal1 17664 9554 17664 9554 0 _0448_
rlabel metal1 20102 17272 20102 17272 0 _0449_
rlabel metal1 16468 8534 16468 8534 0 _0450_
rlabel metal1 21344 15062 21344 15062 0 _0451_
rlabel metal1 18684 21590 18684 21590 0 _0452_
rlabel metal1 15364 18734 15364 18734 0 _0453_
rlabel metal1 13248 21114 13248 21114 0 _0454_
rlabel metal1 19374 8806 19374 8806 0 _0455_
rlabel metal2 17342 19244 17342 19244 0 _0456_
rlabel metal1 20608 14994 20608 14994 0 _0457_
rlabel metal2 15870 19533 15870 19533 0 _0458_
rlabel metal2 13386 15980 13386 15980 0 _0459_
rlabel metal1 17848 20366 17848 20366 0 _0460_
rlabel metal1 13064 20570 13064 20570 0 _0461_
rlabel via1 18178 12886 18178 12886 0 _0462_
rlabel via1 16148 24786 16148 24786 0 _0463_
rlabel metal1 17480 21590 17480 21590 0 _0464_
rlabel metal1 14086 19414 14086 19414 0 _0465_
rlabel metal2 15962 25534 15962 25534 0 _0466_
rlabel metal1 13432 21046 13432 21046 0 _0467_
rlabel metal1 16008 28050 16008 28050 0 _0468_
rlabel metal2 15134 27982 15134 27982 0 _0469_
rlabel metal2 14858 26469 14858 26469 0 _0470_
rlabel metal1 15548 20026 15548 20026 0 _0471_
rlabel metal2 17894 20672 17894 20672 0 _0472_
rlabel viali 19368 20434 19368 20434 0 _0473_
rlabel metal1 17948 21590 17948 21590 0 _0474_
rlabel metal1 18216 16626 18216 16626 0 _0475_
rlabel via3 8533 20740 8533 20740 0 _0476_
rlabel metal1 9338 16660 9338 16660 0 _0477_
rlabel metal1 20010 11254 20010 11254 0 _0478_
rlabel metal2 18906 16694 18906 16694 0 _0479_
rlabel metal1 17664 19890 17664 19890 0 _0480_
rlabel metal1 13018 6868 13018 6868 0 _0481_
rlabel metal2 12650 21284 12650 21284 0 _0482_
rlabel metal1 10856 21318 10856 21318 0 _0483_
rlabel metal1 13570 14450 13570 14450 0 _0484_
rlabel metal1 15242 19414 15242 19414 0 _0485_
rlabel metal2 10718 24718 10718 24718 0 _0486_
rlabel metal1 10488 23086 10488 23086 0 _0487_
rlabel metal1 12052 24174 12052 24174 0 _0488_
rlabel metal1 15502 19822 15502 19822 0 _0489_
rlabel metal2 9614 14603 9614 14603 0 _0490_
rlabel metal1 11270 15504 11270 15504 0 _0491_
rlabel metal1 13708 8942 13708 8942 0 _0492_
rlabel metal1 13524 6766 13524 6766 0 _0493_
rlabel metal2 9890 7684 9890 7684 0 _0494_
rlabel via1 15602 8602 15602 8602 0 _0495_
rlabel metal1 14398 8534 14398 8534 0 _0496_
rlabel metal1 11822 10234 11822 10234 0 _0497_
rlabel metal1 16238 9894 16238 9894 0 _0498_
rlabel metal1 15318 6426 15318 6426 0 _0499_
rlabel metal1 16606 16558 16606 16558 0 _0500_
rlabel metal1 18032 16082 18032 16082 0 _0501_
rlabel metal1 16008 12818 16008 12818 0 _0502_
rlabel metal1 17342 6426 17342 6426 0 _0503_
rlabel metal1 16652 12614 16652 12614 0 _0504_
rlabel metal1 20148 15402 20148 15402 0 _0505_
rlabel metal1 20288 13906 20288 13906 0 _0506_
rlabel metal1 18170 19754 18170 19754 0 _0507_
rlabel metal1 18124 20026 18124 20026 0 _0508_
rlabel metal1 19826 13974 19826 13974 0 _0509_
rlabel metal1 22586 12818 22586 12818 0 _0510_
rlabel metal1 20010 13328 20010 13328 0 _0511_
rlabel metal1 20102 13158 20102 13158 0 _0512_
rlabel metal1 13386 10200 13386 10200 0 _0513_
rlabel metal2 19458 8024 19458 8024 0 _0514_
rlabel metal1 16192 7990 16192 7990 0 _0515_
rlabel metal1 9246 13872 9246 13872 0 _0516_
rlabel metal1 6762 13872 6762 13872 0 _0517_
rlabel metal1 10626 12614 10626 12614 0 _0518_
rlabel metal1 8740 9962 8740 9962 0 _0519_
rlabel metal1 7038 13974 7038 13974 0 _0520_
rlabel metal1 2990 8874 2990 8874 0 _0521_
rlabel metal1 15180 19210 15180 19210 0 _0522_
rlabel metal1 16146 19822 16146 19822 0 _0523_
rlabel metal2 15870 16592 15870 16592 0 _0524_
rlabel metal2 15594 17612 15594 17612 0 _0525_
rlabel metal1 17756 19958 17756 19958 0 _0526_
rlabel metal1 17572 20026 17572 20026 0 _0527_
rlabel metal1 17342 19822 17342 19822 0 _0528_
rlabel metal2 15778 17918 15778 17918 0 _0529_
rlabel metal3 16583 15844 16583 15844 0 _0530_
rlabel metal1 14720 19414 14720 19414 0 _0531_
rlabel metal1 17664 16082 17664 16082 0 _0532_
rlabel metal1 18262 15606 18262 15606 0 _0533_
rlabel metal1 16054 16116 16054 16116 0 _0534_
rlabel metal2 14536 13260 14536 13260 0 _0535_
rlabel metal1 17710 14348 17710 14348 0 _0536_
rlabel metal1 17802 14586 17802 14586 0 _0537_
rlabel metal1 16790 14586 16790 14586 0 _0538_
rlabel metal2 14950 15946 14950 15946 0 _0539_
rlabel metal1 13524 14586 13524 14586 0 _0540_
rlabel metal3 15732 13396 15732 13396 0 _0541_
rlabel metal1 16146 11254 16146 11254 0 _0542_
rlabel metal2 14214 14076 14214 14076 0 _0543_
rlabel metal1 14674 7514 14674 7514 0 _0544_
rlabel metal1 17020 8058 17020 8058 0 _0545_
rlabel metal1 15410 8058 15410 8058 0 _0546_
rlabel metal1 11822 9146 11822 9146 0 _0547_
rlabel metal2 12558 10200 12558 10200 0 _0548_
rlabel metal1 11776 14246 11776 14246 0 _0549_
rlabel metal2 11914 12682 11914 12682 0 _0550_
rlabel metal1 20424 15606 20424 15606 0 _0551_
rlabel metal1 15134 17782 15134 17782 0 _0552_
rlabel metal1 18446 17850 18446 17850 0 _0553_
rlabel metal1 15272 13906 15272 13906 0 _0554_
rlabel metal2 13846 13736 13846 13736 0 _0555_
rlabel metal1 8326 12784 8326 12784 0 _0556_
rlabel metal2 6624 12988 6624 12988 0 _0557_
rlabel metal1 14904 23834 14904 23834 0 _0558_
rlabel metal1 15824 23222 15824 23222 0 _0559_
rlabel metal1 14168 23290 14168 23290 0 _0560_
rlabel metal1 12742 10064 12742 10064 0 _0561_
rlabel metal2 13478 9282 13478 9282 0 _0562_
rlabel metal1 9982 9044 9982 9044 0 _0563_
rlabel metal1 15640 9146 15640 9146 0 _0564_
rlabel metal2 13018 9690 13018 9690 0 _0565_
rlabel metal1 18492 7242 18492 7242 0 _0566_
rlabel metal1 17986 7310 17986 7310 0 _0567_
rlabel metal2 14858 7208 14858 7208 0 _0568_
rlabel metal1 17158 7514 17158 7514 0 _0569_
rlabel metal1 15686 6868 15686 6868 0 _0570_
rlabel metal1 14076 5814 14076 5814 0 _0571_
rlabel metal2 12926 6324 12926 6324 0 _0572_
rlabel metal1 12696 6970 12696 6970 0 _0573_
rlabel metal2 13202 10387 13202 10387 0 _0574_
rlabel metal1 13018 16048 13018 16048 0 _0575_
rlabel metal2 12512 15878 12512 15878 0 _0576_
rlabel metal1 13478 18802 13478 18802 0 _0577_
rlabel metal1 15732 18938 15732 18938 0 _0578_
rlabel metal1 16468 21386 16468 21386 0 _0579_
rlabel metal1 16836 21454 16836 21454 0 _0580_
rlabel metal1 13294 17306 13294 17306 0 _0581_
rlabel metal1 14582 18700 14582 18700 0 _0582_
rlabel metal2 21850 15742 21850 15742 0 _0583_
rlabel metal1 21252 13430 21252 13430 0 _0584_
rlabel metal1 21160 16014 21160 16014 0 _0585_
rlabel metal1 20010 16218 20010 16218 0 _0586_
rlabel metal2 13662 18496 13662 18496 0 _0587_
rlabel metal1 8970 10234 8970 10234 0 _0588_
rlabel metal2 6670 8160 6670 8160 0 _0589_
rlabel metal2 6486 8092 6486 8092 0 _0590_
rlabel metal1 3956 9622 3956 9622 0 _0591_
rlabel via2 2162 18411 2162 18411 0 _0592_
rlabel metal1 16100 14790 16100 14790 0 _0593_
rlabel metal2 17250 12886 17250 12886 0 _0594_
rlabel metal1 16882 14994 16882 14994 0 _0595_
rlabel metal1 15410 14960 15410 14960 0 _0596_
rlabel metal2 13846 12886 13846 12886 0 _0597_
rlabel metal1 17434 12954 17434 12954 0 _0598_
rlabel metal1 14536 15606 14536 15606 0 _0599_
rlabel metal1 14766 14790 14766 14790 0 _0600_
rlabel metal1 17618 14042 17618 14042 0 _0601_
rlabel metal1 15594 14450 15594 14450 0 _0602_
rlabel metal1 17066 12342 17066 12342 0 _0603_
rlabel metal2 16146 14722 16146 14722 0 _0604_
rlabel metal1 15318 12818 15318 12818 0 _0605_
rlabel metal1 14536 12750 14536 12750 0 _0606_
rlabel metal1 15824 10778 15824 10778 0 _0607_
rlabel metal1 14904 12954 14904 12954 0 _0608_
rlabel via2 8970 11747 8970 11747 0 _0609_
rlabel metal2 13938 15147 13938 15147 0 _0610_
rlabel metal1 12972 14858 12972 14858 0 _0611_
rlabel metal1 13662 14994 13662 14994 0 _0612_
rlabel metal1 14030 13294 14030 13294 0 _0613_
rlabel metal1 15824 8602 15824 8602 0 _0614_
rlabel metal1 18492 14518 18492 14518 0 _0615_
rlabel metal1 18906 7990 18906 7990 0 _0616_
rlabel metal1 16008 13498 16008 13498 0 _0617_
rlabel metal2 17618 22338 17618 22338 0 _0618_
rlabel metal1 14720 22474 14720 22474 0 _0619_
rlabel metal1 13708 21862 13708 21862 0 _0620_
rlabel metal2 14398 13651 14398 13651 0 _0621_
rlabel metal2 12190 6919 12190 6919 0 _0622_
rlabel metal1 16698 11594 16698 11594 0 _0623_
rlabel metal1 14904 13226 14904 13226 0 _0624_
rlabel metal1 10074 11798 10074 11798 0 _0625_
rlabel metal1 6808 9146 6808 9146 0 _0626_
rlabel metal1 8924 15130 8924 15130 0 _0627_
rlabel metal1 8004 12614 8004 12614 0 _0628_
rlabel metal1 8234 11526 8234 11526 0 _0629_
rlabel metal1 7544 10710 7544 10710 0 _0630_
rlabel metal4 17204 5984 17204 5984 0 _0631_
rlabel metal1 20240 16014 20240 16014 0 _0632_
rlabel metal1 19596 15946 19596 15946 0 _0633_
rlabel metal2 20516 14076 20516 14076 0 _0634_
rlabel metal2 19366 17136 19366 17136 0 _0635_
rlabel metal1 16928 23834 16928 23834 0 _0636_
rlabel metal1 17204 24174 17204 24174 0 _0637_
rlabel metal2 17802 24480 17802 24480 0 _0638_
rlabel metal1 15410 18054 15410 18054 0 _0639_
rlabel metal3 19849 18020 19849 18020 0 _0640_
rlabel metal2 20654 14688 20654 14688 0 _0641_
rlabel metal1 19550 18734 19550 18734 0 _0642_
rlabel metal2 19458 18462 19458 18462 0 _0643_
rlabel metal1 10580 21658 10580 21658 0 _0644_
rlabel metal1 12604 22610 12604 22610 0 _0645_
rlabel metal2 12558 21216 12558 21216 0 _0646_
rlabel metal2 13340 21964 13340 21964 0 _0647_
rlabel metal1 13846 11764 13846 11764 0 _0648_
rlabel metal1 11408 6290 11408 6290 0 _0649_
rlabel metal2 14122 7888 14122 7888 0 _0650_
rlabel metal2 17250 8806 17250 8806 0 _0651_
rlabel metal1 17480 11118 17480 11118 0 _0652_
rlabel metal2 13662 8262 13662 8262 0 _0653_
rlabel metal1 14858 8602 14858 8602 0 _0654_
rlabel metal2 17526 8194 17526 8194 0 _0655_
rlabel metal2 22494 12665 22494 12665 0 _0656_
rlabel metal1 19826 9044 19826 9044 0 _0657_
rlabel metal2 22310 13532 22310 13532 0 _0658_
rlabel metal1 21390 12614 21390 12614 0 _0659_
rlabel via2 17342 11339 17342 11339 0 _0660_
rlabel metal1 7958 11628 7958 11628 0 _0661_
rlabel metal1 7820 10234 7820 10234 0 _0662_
rlabel metal1 9200 12682 9200 12682 0 _0663_
rlabel metal3 17204 8024 17204 8024 0 _0664_
rlabel metal4 2300 10064 2300 10064 0 _0665_
rlabel metal1 7728 8942 7728 8942 0 _0666_
rlabel metal2 7590 10030 7590 10030 0 _0667_
rlabel metal2 7038 7990 7038 7990 0 _0668_
rlabel metal1 7406 8976 7406 8976 0 _0669_
rlabel metal2 5750 7344 5750 7344 0 _0670_
rlabel metal2 1794 10353 1794 10353 0 _0671_
rlabel metal2 2346 9792 2346 9792 0 _0672_
rlabel metal1 5842 7888 5842 7888 0 _0673_
rlabel metal1 4416 8398 4416 8398 0 _0674_
rlabel metal1 3036 10098 3036 10098 0 _0675_
rlabel metal2 7682 6732 7682 6732 0 _0676_
rlabel metal2 5290 9724 5290 9724 0 _0677_
rlabel metal2 7406 7004 7406 7004 0 _0678_
rlabel metal1 3404 10030 3404 10030 0 _0679_
rlabel metal1 4002 9554 4002 9554 0 _0680_
rlabel metal1 2024 10710 2024 10710 0 _0681_
rlabel metal2 2162 11322 2162 11322 0 _0682_
rlabel metal1 19826 16762 19826 16762 0 _0683_
rlabel metal1 17848 17306 17848 17306 0 _0684_
rlabel metal2 15686 26316 15686 26316 0 _0685_
rlabel metal1 15962 24582 15962 24582 0 _0686_
rlabel metal2 19366 10540 19366 10540 0 _0687_
rlabel metal1 19826 12954 19826 12954 0 _0688_
rlabel metal1 15502 20468 15502 20468 0 _0689_
rlabel metal1 12006 23052 12006 23052 0 _0690_
rlabel metal1 14398 20502 14398 20502 0 _0691_
rlabel metal4 15548 16728 15548 16728 0 _0692_
rlabel metal2 9246 6596 9246 6596 0 _0693_
rlabel metal1 13294 6732 13294 6732 0 _0694_
rlabel metal2 19918 14484 19918 14484 0 _0695_
rlabel metal1 13478 11186 13478 11186 0 _0696_
rlabel metal1 13386 9452 13386 9452 0 _0697_
rlabel metal3 15686 14348 15686 14348 0 _0698_
rlabel metal1 13064 5746 13064 5746 0 _0699_
rlabel metal1 15962 5542 15962 5542 0 _0700_
rlabel metal1 14260 8806 14260 8806 0 _0701_
rlabel metal1 9430 13260 9430 13260 0 _0702_
rlabel metal1 9522 13498 9522 13498 0 _0703_
rlabel metal1 9200 15334 9200 15334 0 _0704_
rlabel metal2 1978 11458 1978 11458 0 _0705_
rlabel metal1 4830 9520 4830 9520 0 _0706_
rlabel via2 6670 5219 6670 5219 0 _0707_
rlabel metal1 4508 9554 4508 9554 0 _0708_
rlabel metal2 4186 8636 4186 8636 0 _0709_
rlabel metal1 4370 8942 4370 8942 0 _0710_
rlabel metal2 2714 10098 2714 10098 0 _0711_
rlabel metal1 1794 12138 1794 12138 0 _0712_
rlabel metal1 4416 12750 4416 12750 0 _0713_
rlabel metal1 4692 12818 4692 12818 0 _0714_
rlabel metal1 2438 8976 2438 8976 0 _0715_
rlabel metal1 1978 3094 1978 3094 0 _0716_
rlabel metal2 1610 6460 1610 6460 0 _0717_
rlabel via1 2714 12869 2714 12869 0 _0718_
rlabel metal1 4876 9146 4876 9146 0 _0719_
rlabel metal1 1978 13804 1978 13804 0 _0720_
rlabel metal1 5198 13906 5198 13906 0 _0721_
rlabel metal1 5244 15470 5244 15470 0 _0722_
rlabel metal2 7590 15351 7590 15351 0 _0723_
rlabel metal2 2254 16932 2254 16932 0 _0724_
rlabel metal2 2162 14433 2162 14433 0 _0725_
rlabel metal1 2622 12784 2622 12784 0 _0726_
rlabel metal1 2024 12954 2024 12954 0 _0727_
rlabel metal1 5198 16082 5198 16082 0 _0728_
rlabel metal1 1886 13736 1886 13736 0 _0729_
rlabel via2 5014 4811 5014 4811 0 _0730_
rlabel metal1 1978 13940 1978 13940 0 _0731_
rlabel metal1 2392 13906 2392 13906 0 _0732_
rlabel metal1 1794 16558 1794 16558 0 _0733_
rlabel metal2 2346 14518 2346 14518 0 _0734_
rlabel metal1 2208 17170 2208 17170 0 _0735_
rlabel metal2 2806 19618 2806 19618 0 _0736_
rlabel metal1 1380 8942 1380 8942 0 _0737_
rlabel metal1 6440 20026 6440 20026 0 _0738_
rlabel metal1 7133 19482 7133 19482 0 _0739_
rlabel metal1 3864 19958 3864 19958 0 _0740_
rlabel metal2 21298 23800 21298 23800 0 _0741_
rlabel metal1 3496 22202 3496 22202 0 _0742_
rlabel metal1 4370 22644 4370 22644 0 _0743_
rlabel metal1 2369 23834 2369 23834 0 _0744_
rlabel metal2 2162 22117 2162 22117 0 _0745_
rlabel metal1 3634 31790 3634 31790 0 _0746_
rlabel metal1 4278 21046 4278 21046 0 _0747_
rlabel metal2 2070 16082 2070 16082 0 _0748_
rlabel metal1 2254 14960 2254 14960 0 _0749_
rlabel metal1 2116 17578 2116 17578 0 _0750_
rlabel metal1 2070 18666 2070 18666 0 _0751_
rlabel metal1 2162 17680 2162 17680 0 _0752_
rlabel metal2 4002 18598 4002 18598 0 _0753_
rlabel metal2 5750 12070 5750 12070 0 _0754_
rlabel metal1 6118 19346 6118 19346 0 _0755_
rlabel metal1 4784 18938 4784 18938 0 _0756_
rlabel metal1 3729 19482 3729 19482 0 _0757_
rlabel metal2 7774 19159 7774 19159 0 _0758_
rlabel metal2 10258 25041 10258 25041 0 _0759_
rlabel metal1 2254 19380 2254 19380 0 _0760_
rlabel metal2 1794 20366 1794 20366 0 _0761_
rlabel via2 3082 21539 3082 21539 0 _0762_
rlabel metal2 9246 26010 9246 26010 0 _0763_
rlabel metal1 12052 14518 12052 14518 0 _0764_
rlabel metal1 5612 15674 5612 15674 0 _0765_
rlabel metal1 5612 16762 5612 16762 0 _0766_
rlabel via1 4536 18258 4536 18258 0 _0767_
rlabel metal1 4554 18054 4554 18054 0 _0768_
rlabel metal1 3064 20910 3064 20910 0 _0769_
rlabel metal1 2530 23732 2530 23732 0 _0770_
rlabel via2 1794 23749 1794 23749 0 _0771_
rlabel metal1 2208 22610 2208 22610 0 _0772_
rlabel metal1 6026 28390 6026 28390 0 _0773_
rlabel metal1 3818 14586 3818 14586 0 _0774_
rlabel metal1 5198 15878 5198 15878 0 _0775_
rlabel metal2 3266 16626 3266 16626 0 _0776_
rlabel metal1 4462 14416 4462 14416 0 _0777_
rlabel metal1 3496 14246 3496 14246 0 _0778_
rlabel via1 2880 18258 2880 18258 0 _0779_
rlabel metal1 1886 20944 1886 20944 0 _0780_
rlabel via1 1702 20910 1702 20910 0 _0781_
rlabel metal1 2438 21114 2438 21114 0 _0782_
rlabel metal2 4094 23426 4094 23426 0 _0783_
rlabel metal2 26082 27523 26082 27523 0 _0784_
rlabel metal1 1702 15674 1702 15674 0 _0785_
rlabel metal1 5244 15606 5244 15606 0 _0786_
rlabel metal1 3984 17170 3984 17170 0 _0787_
rlabel metal1 5152 17306 5152 17306 0 _0788_
rlabel metal1 5152 21658 5152 21658 0 _0789_
rlabel metal1 7912 22202 7912 22202 0 _0790_
rlabel metal1 4646 21998 4646 21998 0 _0791_
rlabel metal2 1794 17748 1794 17748 0 _0792_
rlabel metal1 3174 18802 3174 18802 0 _0793_
rlabel metal2 3082 17306 3082 17306 0 _0794_
rlabel metal1 1748 9146 1748 9146 0 _0795_
rlabel metal1 3312 18938 3312 18938 0 _0796_
rlabel metal1 4922 19210 4922 19210 0 _0797_
rlabel metal1 5290 22542 5290 22542 0 _0798_
rlabel metal1 5336 22746 5336 22746 0 _0799_
rlabel metal2 9706 24599 9706 24599 0 _0800_
rlabel metal1 6900 25738 6900 25738 0 _0801_
rlabel metal1 5382 23120 5382 23120 0 _0802_
rlabel metal1 4738 22950 4738 22950 0 _0803_
rlabel via2 5842 24803 5842 24803 0 _0804_
rlabel metal1 3174 19822 3174 19822 0 _0805_
rlabel metal1 4554 23494 4554 23494 0 _0806_
rlabel metal2 4002 20740 4002 20740 0 _0807_
rlabel metal1 5842 16116 5842 16116 0 _0808_
rlabel metal1 7636 13294 7636 13294 0 _0809_
rlabel metal2 9522 15232 9522 15232 0 _0810_
rlabel metal1 9062 12852 9062 12852 0 _0811_
rlabel metal1 6072 5678 6072 5678 0 _0812_
rlabel via2 5842 5083 5842 5083 0 _0813_
rlabel metal1 4324 5678 4324 5678 0 _0814_
rlabel metal2 18722 6035 18722 6035 0 _0815_
rlabel metal3 5359 19516 5359 19516 0 _0816_
rlabel metal2 22034 27506 22034 27506 0 _0817_
rlabel metal1 3772 17850 3772 17850 0 _0818_
rlabel metal2 4278 17578 4278 17578 0 _0819_
rlabel metal1 5796 18802 5796 18802 0 _0820_
rlabel metal2 4370 19822 4370 19822 0 _0821_
rlabel metal1 6532 21114 6532 21114 0 _0822_
rlabel metal1 10028 27098 10028 27098 0 _0823_
rlabel metal1 3220 31926 3220 31926 0 _0824_
rlabel metal2 21390 27489 21390 27489 0 _0825_
rlabel metal2 14582 25500 14582 25500 0 _0826_
rlabel metal1 8556 17102 8556 17102 0 _0827_
rlabel metal1 9844 21114 9844 21114 0 _0828_
rlabel metal1 9752 23834 9752 23834 0 _0829_
rlabel metal2 2346 32708 2346 32708 0 _0830_
rlabel metal1 3542 32232 3542 32232 0 _0831_
rlabel metal2 9154 23001 9154 23001 0 _0832_
rlabel metal1 11500 23834 11500 23834 0 _0833_
rlabel metal1 10258 25466 10258 25466 0 _0834_
rlabel metal3 17204 24616 17204 24616 0 _0835_
rlabel metal2 2438 11152 2438 11152 0 _0836_
rlabel metal1 11132 5678 11132 5678 0 _0837_
rlabel metal1 12742 19822 12742 19822 0 _0838_
rlabel metal1 1518 24786 1518 24786 0 _0839_
rlabel metal2 8602 6970 8602 6970 0 _0840_
rlabel metal1 15318 17544 15318 17544 0 _0841_
rlabel metal2 10626 8330 10626 8330 0 _0842_
rlabel metal1 5290 5202 5290 5202 0 _0843_
rlabel metal2 5106 4777 5106 4777 0 _0844_
rlabel metal1 5980 6630 5980 6630 0 _0845_
rlabel metal2 11178 11373 11178 11373 0 _0846_
rlabel metal1 7544 22746 7544 22746 0 _0847_
rlabel metal1 9154 22712 9154 22712 0 _0848_
rlabel metal1 11316 18258 11316 18258 0 _0849_
rlabel metal2 17158 17391 17158 17391 0 _0850_
rlabel metal1 17940 19346 17940 19346 0 _0851_
rlabel metal1 14812 17170 14812 17170 0 _0852_
rlabel metal2 16238 17612 16238 17612 0 _0853_
rlabel metal2 21206 19516 21206 19516 0 _0854_
rlabel metal1 23874 16422 23874 16422 0 _0855_
rlabel metal1 25024 16218 25024 16218 0 _0856_
rlabel metal2 22494 17340 22494 17340 0 _0857_
rlabel metal1 19826 18802 19826 18802 0 _0858_
rlabel metal1 18906 19278 18906 19278 0 _0859_
rlabel metal1 17756 20570 17756 20570 0 _0860_
rlabel metal2 15686 16490 15686 16490 0 _0861_
rlabel metal1 15732 14586 15732 14586 0 _0862_
rlabel metal1 19642 19822 19642 19822 0 _0863_
rlabel metal1 20332 20026 20332 20026 0 _0864_
rlabel metal1 21298 23732 21298 23732 0 _0865_
rlabel metal2 18906 23732 18906 23732 0 _0866_
rlabel metal1 20194 22746 20194 22746 0 _0867_
rlabel metal1 20562 24378 20562 24378 0 _0868_
rlabel metal1 20010 23290 20010 23290 0 _0869_
rlabel metal1 19044 24718 19044 24718 0 _0870_
rlabel metal1 17526 22746 17526 22746 0 _0871_
rlabel metal1 9200 19822 9200 19822 0 _0872_
rlabel metal1 13018 22066 13018 22066 0 _0873_
rlabel metal2 12374 24786 12374 24786 0 _0874_
rlabel metal1 16376 29274 16376 29274 0 _0875_
rlabel metal1 19320 27438 19320 27438 0 _0876_
rlabel metal1 18400 25806 18400 25806 0 _0877_
rlabel metal1 13432 23834 13432 23834 0 _0878_
rlabel metal1 9568 18394 9568 18394 0 _0879_
rlabel metal1 10580 13838 10580 13838 0 _0880_
rlabel metal1 11086 12954 11086 12954 0 _0881_
rlabel metal2 11822 11594 11822 11594 0 _0882_
rlabel metal1 14306 14586 14306 14586 0 _0883_
rlabel metal1 10718 9384 10718 9384 0 cal_lut\[100\]
rlabel metal1 13984 12954 13984 12954 0 cal_lut\[101\]
rlabel metal1 15180 11254 15180 11254 0 cal_lut\[102\]
rlabel metal1 19780 15402 19780 15402 0 cal_lut\[103\]
rlabel via1 19992 17170 19992 17170 0 cal_lut\[104\]
rlabel via2 19550 8483 19550 8483 0 cal_lut\[105\]
rlabel metal1 18722 8568 18722 8568 0 cal_lut\[106\]
rlabel metal2 20194 11560 20194 11560 0 cal_lut\[107\]
rlabel via2 19642 11067 19642 11067 0 cal_lut\[108\]
rlabel metal1 21298 11016 21298 11016 0 cal_lut\[109\]
rlabel metal1 14306 17136 14306 17136 0 cal_lut\[10\]
rlabel metal1 20700 13226 20700 13226 0 cal_lut\[110\]
rlabel via2 19918 7837 19918 7837 0 cal_lut\[111\]
rlabel metal1 18124 7854 18124 7854 0 cal_lut\[112\]
rlabel metal1 19734 6868 19734 6868 0 cal_lut\[113\]
rlabel metal1 19090 9622 19090 9622 0 cal_lut\[114\]
rlabel metal1 19872 10234 19872 10234 0 cal_lut\[115\]
rlabel metal2 20838 10438 20838 10438 0 cal_lut\[116\]
rlabel metal1 20148 9418 20148 9418 0 cal_lut\[117\]
rlabel metal1 18814 5678 18814 5678 0 cal_lut\[118\]
rlabel via3 17549 12444 17549 12444 0 cal_lut\[119\]
rlabel metal1 15732 18258 15732 18258 0 cal_lut\[11\]
rlabel metal1 13662 4148 13662 4148 0 cal_lut\[120\]
rlabel metal1 10672 1326 10672 1326 0 cal_lut\[121\]
rlabel metal2 9798 4012 9798 4012 0 cal_lut\[122\]
rlabel metal1 11822 4692 11822 4692 0 cal_lut\[123\]
rlabel metal1 14444 4590 14444 4590 0 cal_lut\[124\]
rlabel metal1 14490 6120 14490 6120 0 cal_lut\[125\]
rlabel metal1 12650 4624 12650 4624 0 cal_lut\[126\]
rlabel metal2 13570 3162 13570 3162 0 cal_lut\[127\]
rlabel metal1 15732 1326 15732 1326 0 cal_lut\[128\]
rlabel metal2 23506 1632 23506 1632 0 cal_lut\[129\]
rlabel metal1 21068 19346 21068 19346 0 cal_lut\[12\]
rlabel metal2 23414 2108 23414 2108 0 cal_lut\[130\]
rlabel metal1 17572 5814 17572 5814 0 cal_lut\[131\]
rlabel metal1 18170 4726 18170 4726 0 cal_lut\[132\]
rlabel metal1 22218 2584 22218 2584 0 cal_lut\[133\]
rlabel metal2 17710 4998 17710 4998 0 cal_lut\[134\]
rlabel metal2 20838 952 20838 952 0 cal_lut\[135\]
rlabel metal1 16100 1462 16100 1462 0 cal_lut\[136\]
rlabel metal1 16790 2618 16790 2618 0 cal_lut\[137\]
rlabel metal2 13110 5406 13110 5406 0 cal_lut\[138\]
rlabel metal2 4738 2142 4738 2142 0 cal_lut\[139\]
rlabel metal1 23736 16694 23736 16694 0 cal_lut\[13\]
rlabel metal1 3910 4216 3910 4216 0 cal_lut\[140\]
rlabel metal1 6900 2890 6900 2890 0 cal_lut\[141\]
rlabel metal2 7406 2210 7406 2210 0 cal_lut\[142\]
rlabel metal1 10764 2618 10764 2618 0 cal_lut\[143\]
rlabel metal1 14490 1802 14490 1802 0 cal_lut\[144\]
rlabel metal1 13846 3162 13846 3162 0 cal_lut\[145\]
rlabel metal2 15594 1190 15594 1190 0 cal_lut\[146\]
rlabel metal2 23414 952 23414 952 0 cal_lut\[147\]
rlabel metal1 25806 1190 25806 1190 0 cal_lut\[148\]
rlabel metal1 20608 5066 20608 5066 0 cal_lut\[149\]
rlabel metal1 23920 15946 23920 15946 0 cal_lut\[14\]
rlabel via2 21022 6171 21022 6171 0 cal_lut\[150\]
rlabel metal1 20424 12818 20424 12818 0 cal_lut\[151\]
rlabel metal1 21850 10166 21850 10166 0 cal_lut\[152\]
rlabel metal1 20470 14552 20470 14552 0 cal_lut\[153\]
rlabel metal1 21436 13498 21436 13498 0 cal_lut\[154\]
rlabel metal1 18170 12648 18170 12648 0 cal_lut\[155\]
rlabel metal1 17112 13430 17112 13430 0 cal_lut\[156\]
rlabel metal1 20056 17034 20056 17034 0 cal_lut\[157\]
rlabel metal2 22310 21199 22310 21199 0 cal_lut\[158\]
rlabel metal1 20470 17782 20470 17782 0 cal_lut\[159\]
rlabel metal2 22402 16592 22402 16592 0 cal_lut\[15\]
rlabel metal1 22862 16694 22862 16694 0 cal_lut\[160\]
rlabel metal1 22011 19346 22011 19346 0 cal_lut\[161\]
rlabel metal2 16238 19635 16238 19635 0 cal_lut\[162\]
rlabel metal1 25944 20774 25944 20774 0 cal_lut\[163\]
rlabel metal1 26680 15878 26680 15878 0 cal_lut\[164\]
rlabel metal2 25990 15096 25990 15096 0 cal_lut\[165\]
rlabel metal1 21873 15674 21873 15674 0 cal_lut\[166\]
rlabel metal2 22770 13362 22770 13362 0 cal_lut\[167\]
rlabel metal1 21114 15606 21114 15606 0 cal_lut\[168\]
rlabel metal1 26404 14790 26404 14790 0 cal_lut\[169\]
rlabel metal1 18722 18802 18722 18802 0 cal_lut\[16\]
rlabel metal1 25484 13498 25484 13498 0 cal_lut\[170\]
rlabel metal1 23368 12954 23368 12954 0 cal_lut\[171\]
rlabel metal1 20562 8908 20562 8908 0 cal_lut\[172\]
rlabel metal1 21482 13736 21482 13736 0 cal_lut\[173\]
rlabel metal2 20378 15810 20378 15810 0 cal_lut\[174\]
rlabel metal1 26174 16626 26174 16626 0 cal_lut\[175\]
rlabel metal1 20930 14926 20930 14926 0 cal_lut\[176\]
rlabel metal1 23322 5814 23322 5814 0 cal_lut\[177\]
rlabel metal1 25254 2278 25254 2278 0 cal_lut\[178\]
rlabel metal1 21206 3638 21206 3638 0 cal_lut\[179\]
rlabel viali 18261 19346 18261 19346 0 cal_lut\[17\]
rlabel metal2 17434 5712 17434 5712 0 cal_lut\[180\]
rlabel metal2 20654 4658 20654 4658 0 cal_lut\[181\]
rlabel via2 19826 3621 19826 3621 0 cal_lut\[182\]
rlabel metal2 20470 3927 20470 3927 0 cal_lut\[183\]
rlabel metal1 25852 2618 25852 2618 0 cal_lut\[184\]
rlabel metal3 16767 12716 16767 12716 0 cal_lut\[185\]
rlabel metal3 16537 13124 16537 13124 0 cal_lut\[186\]
rlabel metal2 12006 8415 12006 8415 0 cal_lut\[187\]
rlabel metal1 12972 5338 12972 5338 0 cal_lut\[188\]
rlabel metal1 10580 4794 10580 4794 0 cal_lut\[189\]
rlabel metal2 17526 20077 17526 20077 0 cal_lut\[18\]
rlabel metal1 7912 1190 7912 1190 0 cal_lut\[190\]
rlabel metal1 11500 12614 11500 12614 0 cal_lut\[191\]
rlabel metal1 14996 7174 14996 7174 0 cal_lut\[192\]
rlabel metal3 19067 22644 19067 22644 0 cal_lut\[19\]
rlabel metal2 8418 2329 8418 2329 0 cal_lut\[1\]
rlabel metal2 20102 14620 20102 14620 0 cal_lut\[20\]
rlabel metal1 19596 19958 19596 19958 0 cal_lut\[21\]
rlabel metal1 17687 18666 17687 18666 0 cal_lut\[22\]
rlabel via3 16445 17884 16445 17884 0 cal_lut\[23\]
rlabel metal1 18584 16218 18584 16218 0 cal_lut\[24\]
rlabel metal1 20056 24310 20056 24310 0 cal_lut\[25\]
rlabel metal3 19343 20604 19343 20604 0 cal_lut\[26\]
rlabel metal1 19642 24344 19642 24344 0 cal_lut\[27\]
rlabel metal1 17434 22610 17434 22610 0 cal_lut\[28\]
rlabel metal1 12696 21930 12696 21930 0 cal_lut\[29\]
rlabel metal2 10534 8160 10534 8160 0 cal_lut\[2\]
rlabel via3 14053 17884 14053 17884 0 cal_lut\[30\]
rlabel metal1 16192 29002 16192 29002 0 cal_lut\[31\]
rlabel metal2 22954 32402 22954 32402 0 cal_lut\[32\]
rlabel metal1 18952 25738 18952 25738 0 cal_lut\[33\]
rlabel metal2 15870 21869 15870 21869 0 cal_lut\[34\]
rlabel metal1 13478 18938 13478 18938 0 cal_lut\[35\]
rlabel metal2 12742 14960 12742 14960 0 cal_lut\[36\]
rlabel metal1 11638 13430 11638 13430 0 cal_lut\[37\]
rlabel metal2 12374 11390 12374 11390 0 cal_lut\[38\]
rlabel metal1 14260 14518 14260 14518 0 cal_lut\[39\]
rlabel metal1 9246 8330 9246 8330 0 cal_lut\[3\]
rlabel metal1 12650 17000 12650 17000 0 cal_lut\[40\]
rlabel metal2 12558 19873 12558 19873 0 cal_lut\[41\]
rlabel metal3 13501 17884 13501 17884 0 cal_lut\[42\]
rlabel metal2 13846 29274 13846 29274 0 cal_lut\[43\]
rlabel metal1 10074 32402 10074 32402 0 cal_lut\[44\]
rlabel metal1 11316 31654 11316 31654 0 cal_lut\[45\]
rlabel metal2 14812 29546 14812 29546 0 cal_lut\[46\]
rlabel metal1 13340 30022 13340 30022 0 cal_lut\[47\]
rlabel metal1 13846 25262 13846 25262 0 cal_lut\[48\]
rlabel metal1 10580 23018 10580 23018 0 cal_lut\[49\]
rlabel metal2 8234 4046 8234 4046 0 cal_lut\[4\]
rlabel metal1 10304 31926 10304 31926 0 cal_lut\[50\]
rlabel metal1 13340 22746 13340 22746 0 cal_lut\[51\]
rlabel metal2 15134 26860 15134 26860 0 cal_lut\[52\]
rlabel via3 13317 19244 13317 19244 0 cal_lut\[53\]
rlabel metal3 14697 19380 14697 19380 0 cal_lut\[54\]
rlabel metal1 14444 31654 14444 31654 0 cal_lut\[55\]
rlabel metal1 12604 32266 12604 32266 0 cal_lut\[56\]
rlabel metal1 14950 30056 14950 30056 0 cal_lut\[57\]
rlabel metal1 15134 32198 15134 32198 0 cal_lut\[58\]
rlabel metal1 15824 19958 15824 19958 0 cal_lut\[59\]
rlabel metal1 5980 1530 5980 1530 0 cal_lut\[5\]
rlabel metal1 19366 29104 19366 29104 0 cal_lut\[60\]
rlabel metal1 14720 28050 14720 28050 0 cal_lut\[61\]
rlabel metal2 22402 29342 22402 29342 0 cal_lut\[62\]
rlabel metal1 20056 32198 20056 32198 0 cal_lut\[63\]
rlabel metal1 21298 31178 21298 31178 0 cal_lut\[64\]
rlabel metal1 19780 25194 19780 25194 0 cal_lut\[65\]
rlabel metal1 17802 21114 17802 21114 0 cal_lut\[66\]
rlabel metal1 25530 21862 25530 21862 0 cal_lut\[67\]
rlabel metal2 20194 19159 20194 19159 0 cal_lut\[68\]
rlabel metal1 21804 22134 21804 22134 0 cal_lut\[69\]
rlabel metal1 8648 10642 8648 10642 0 cal_lut\[6\]
rlabel metal1 20056 23698 20056 23698 0 cal_lut\[70\]
rlabel metal2 20470 21471 20470 21471 0 cal_lut\[71\]
rlabel metal2 20930 20536 20930 20536 0 cal_lut\[72\]
rlabel via1 19624 20910 19624 20910 0 cal_lut\[73\]
rlabel metal2 21574 20672 21574 20672 0 cal_lut\[74\]
rlabel metal1 20792 20842 20792 20842 0 cal_lut\[75\]
rlabel metal1 19826 21454 19826 21454 0 cal_lut\[76\]
rlabel via1 20654 20315 20654 20315 0 cal_lut\[77\]
rlabel metal1 19734 21590 19734 21590 0 cal_lut\[78\]
rlabel metal2 21022 17833 21022 17833 0 cal_lut\[79\]
rlabel metal1 10350 23052 10350 23052 0 cal_lut\[7\]
rlabel metal2 19642 17527 19642 17527 0 cal_lut\[80\]
rlabel metal2 21574 16983 21574 16983 0 cal_lut\[81\]
rlabel metal1 19688 24650 19688 24650 0 cal_lut\[82\]
rlabel metal2 17710 25806 17710 25806 0 cal_lut\[83\]
rlabel metal1 18952 21386 18952 21386 0 cal_lut\[84\]
rlabel metal2 24978 28339 24978 28339 0 cal_lut\[85\]
rlabel metal1 17618 33626 17618 33626 0 cal_lut\[86\]
rlabel metal3 17733 31756 17733 31756 0 cal_lut\[87\]
rlabel metal1 16238 21964 16238 21964 0 cal_lut\[88\]
rlabel metal1 13892 22406 13892 22406 0 cal_lut\[89\]
rlabel metal1 10074 26350 10074 26350 0 cal_lut\[8\]
rlabel metal2 14122 20281 14122 20281 0 cal_lut\[90\]
rlabel metal2 8878 24752 8878 24752 0 cal_lut\[91\]
rlabel metal1 8326 24174 8326 24174 0 cal_lut\[92\]
rlabel metal2 10258 21699 10258 21699 0 cal_lut\[93\]
rlabel metal2 11730 20774 11730 20774 0 cal_lut\[94\]
rlabel metal1 11868 14790 11868 14790 0 cal_lut\[95\]
rlabel metal1 12880 13702 12880 13702 0 cal_lut\[96\]
rlabel metal1 12765 8602 12765 8602 0 cal_lut\[97\]
rlabel metal1 10764 9894 10764 9894 0 cal_lut\[98\]
rlabel metal1 9246 2074 9246 2074 0 cal_lut\[99\]
rlabel metal2 12926 24140 12926 24140 0 cal_lut\[9\]
rlabel metal2 2622 24752 2622 24752 0 clknet_0__0380_
rlabel metal2 2622 15436 2622 15436 0 clknet_0_io_in[0]
rlabel metal2 1610 30906 1610 30906 0 clknet_0_net57
rlabel metal2 15686 29325 15686 29325 0 clknet_0_temp1.dcdel_capnode_notouch_
rlabel metal1 4738 30158 4738 30158 0 clknet_0_temp1.i_precharge_n
rlabel metal1 3036 23154 3036 23154 0 clknet_1_0__leaf__0380_
rlabel metal2 1610 1904 1610 1904 0 clknet_1_0__leaf_io_in[0]
rlabel via2 4094 26843 4094 26843 0 clknet_1_0__leaf_net57
rlabel metal1 14352 32402 14352 32402 0 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_
rlabel metal2 2622 30566 2622 30566 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal1 4830 26452 4830 26452 0 clknet_1_1__leaf__0380_
rlabel metal1 1610 22576 1610 22576 0 clknet_1_1__leaf_io_in[0]
rlabel metal4 17204 29444 17204 29444 0 clknet_1_1__leaf_net57
rlabel metal1 19136 28730 19136 28730 0 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_
rlabel metal2 15870 29291 15870 29291 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal1 2254 20434 2254 20434 0 ctr\[0\]
rlabel metal2 13202 9809 13202 9809 0 ctr\[10\]
rlabel via3 3749 16660 3749 16660 0 ctr\[11\]
rlabel metal1 4416 1190 4416 1190 0 ctr\[12\]
rlabel metal1 1058 11730 1058 11730 0 ctr\[1\]
rlabel metal1 690 11866 690 11866 0 ctr\[2\]
rlabel metal1 5980 18598 5980 18598 0 ctr\[3\]
rlabel metal1 5612 24922 5612 24922 0 ctr\[4\]
rlabel metal1 6532 16150 6532 16150 0 ctr\[5\]
rlabel via2 6670 20995 6670 20995 0 ctr\[6\]
rlabel metal2 2714 8755 2714 8755 0 ctr\[7\]
rlabel metal2 2530 4743 2530 4743 0 ctr\[8\]
rlabel metal1 7544 12750 7544 12750 0 ctr\[9\]
rlabel metal1 7314 21590 7314 21590 0 dbg3\[0\]
rlabel metal2 7268 23732 7268 23732 0 dbg3\[1\]
rlabel metal1 7268 19346 7268 19346 0 dbg3\[2\]
rlabel metal2 6808 22508 6808 22508 0 dbg3\[3\]
rlabel metal1 7774 19346 7774 19346 0 dbg3\[4\]
rlabel metal1 3266 24038 3266 24038 0 dbg3\[5\]
rlabel metal2 2070 13872 2070 13872 0 dec1.i_ones
rlabel metal2 2898 13719 2898 13719 0 io_in[0]
rlabel metal3 406 3740 406 3740 0 io_in[1]
rlabel metal3 406 5780 406 5780 0 io_in[2]
rlabel via2 15778 9333 15778 9333 0 io_in[3]
rlabel metal3 406 9860 406 9860 0 io_in[4]
rlabel metal4 5612 7888 5612 7888 0 io_in[5]
rlabel metal3 406 13940 406 13940 0 io_in[6]
rlabel metal3 406 15980 406 15980 0 io_in[7]
rlabel metal3 452 18020 452 18020 0 io_out[0]
rlabel metal3 406 20060 406 20060 0 io_out[1]
rlabel metal3 406 22100 406 22100 0 io_out[2]
rlabel metal1 4416 23766 4416 23766 0 io_out[3]
rlabel metal1 4048 22066 4048 22066 0 io_out[4]
rlabel metal3 406 28220 406 28220 0 io_out[5]
rlabel metal3 1119 30260 1119 30260 0 io_out[6]
rlabel metal3 1878 32300 1878 32300 0 io_out[7]
rlabel metal1 12880 9622 12880 9622 0 net1
rlabel metal1 12650 28560 12650 28560 0 net10
rlabel metal1 15456 27438 15456 27438 0 net11
rlabel metal2 8510 32504 8510 32504 0 net12
rlabel metal1 6072 31314 6072 31314 0 net13
rlabel metal1 4646 1938 4646 1938 0 net14
rlabel metal1 9890 2414 9890 2414 0 net15
rlabel metal1 13800 5134 13800 5134 0 net16
rlabel metal1 6716 1326 6716 1326 0 net17
rlabel metal1 20148 2414 20148 2414 0 net18
rlabel metal2 19458 6528 19458 6528 0 net19
rlabel metal2 16422 18785 16422 18785 0 net2
rlabel metal1 22632 2482 22632 2482 0 net20
rlabel metal1 24518 2414 24518 2414 0 net21
rlabel metal2 21758 7174 21758 7174 0 net22
rlabel metal2 26450 6256 26450 6256 0 net23
rlabel metal2 26450 12784 26450 12784 0 net24
rlabel metal1 23920 12818 23920 12818 0 net25
rlabel metal1 19274 14790 19274 14790 0 net26
rlabel metal2 12650 25024 12650 25024 0 net27
rlabel metal1 10442 29614 10442 29614 0 net28
rlabel metal1 26910 19890 26910 19890 0 net29
rlabel metal2 16146 8925 16146 8925 0 net3
rlabel metal1 26404 22066 26404 22066 0 net30
rlabel metal1 23276 17510 23276 17510 0 net31
rlabel metal1 19412 28934 19412 28934 0 net32
rlabel metal2 19458 32062 19458 32062 0 net33
rlabel metal1 16882 27948 16882 27948 0 net34
rlabel metal1 21804 25806 21804 25806 0 net35
rlabel metal1 21804 31246 21804 31246 0 net36
rlabel metal1 22586 25228 22586 25228 0 net37
rlabel metal3 18147 21964 18147 21964 0 net38
rlabel metal1 27324 31246 27324 31246 0 net39
rlabel metal1 6624 9622 6624 9622 0 net4
rlabel metal2 14490 32912 14490 32912 0 net40
rlabel metal1 24012 32742 24012 32742 0 net41
rlabel metal2 23506 29614 23506 29614 0 net42
rlabel metal1 24518 32334 24518 32334 0 net43
rlabel metal1 28014 32266 28014 32266 0 net44
rlabel metal1 24012 32470 24012 32470 0 net45
rlabel metal1 24794 30736 24794 30736 0 net46
rlabel metal2 22862 29206 22862 29206 0 net47
rlabel metal1 27370 26928 27370 26928 0 net48
rlabel metal1 26496 30906 26496 30906 0 net49
rlabel metal1 5336 3978 5336 3978 0 net5
rlabel metal1 24104 28662 24104 28662 0 net50
rlabel metal1 26726 32402 26726 32402 0 net51
rlabel metal1 24610 28050 24610 28050 0 net52
rlabel metal1 26910 31926 26910 31926 0 net53
rlabel metal1 23092 28730 23092 28730 0 net54
rlabel metal1 18400 27506 18400 27506 0 net55
rlabel metal1 10534 26826 10534 26826 0 net56
rlabel via2 2530 31331 2530 31331 0 net57
rlabel via2 2162 30277 2162 30277 0 net58
rlabel via2 2438 29597 2438 29597 0 net59
rlabel metal1 3220 5882 3220 5882 0 net6
rlabel metal2 2898 32028 2898 32028 0 net60
rlabel metal1 2622 15436 2622 15436 0 net7
rlabel metal1 7682 29240 7682 29240 0 net8
rlabel metal1 6716 30702 6716 30702 0 net9
rlabel metal1 8004 25874 8004 25874 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 14674 29240 14674 29240 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal4 7636 24072 7636 24072 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel via2 9154 26435 9154 26435 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 5290 27693 5290 27693 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 3358 32232 3358 32232 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal2 16790 33218 16790 33218 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal2 27370 32538 27370 32538 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal1 9154 27880 9154 27880 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 6624 32334 6624 32334 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal1 7452 32334 7452 32334 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal1 10764 32266 10764 32266 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 16514 33048 16514 33048 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal2 14398 28526 14398 28526 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal3 17388 30872 17388 30872 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal2 13662 20247 13662 20247 0 temp1.dac.vdac_single.en_pupd
rlabel metal2 5198 32402 5198 32402 0 temp1.dac_vout_notouch_
rlabel metal1 15042 31790 15042 31790 0 temp1.dcdel_capnode_notouch_
rlabel metal2 14766 26401 14766 26401 0 temp1.i_precharge_n
rlabel metal2 3174 28288 3174 28288 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>
