* PEX produced on Sun Apr 23 11:24:37 AM CEST 2023 using /foss/tools/iic-osic/iic-pex.sh with m=1 and s=1
* NGSPICE file created from hpretl_tt03_temperature_sensor_golden.ext - technology: sky130A

.subckt hpretl_tt03_temperature_sensor io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_in[0] vccd1 vssd1
X0 a_18041_32143# a_17507_32149# a_17946_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1 a_11960_29967# a_11711_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2 vccd1 a_23903_26922# _1342_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3 a_27859_29098# _1451_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4 vssd1 a_21051_24746# _1887_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5 a_14223_1679# a_13441_1685# a_14139_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 vssd1 a_28015_5755# a_27973_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7 _1234_.A1 a_2807_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_19973_32149# a_19807_32149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 vccd1 a_25455_27613# a_25623_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 vccd1 a_24087_20394# _1525_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13 a_13311_25615# a_12447_25621# a_13054_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15 a_9037_9661# a_8767_9295# a_8947_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 a_6186_21041# _1327_.A1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X18 a_27379_24349# a_26597_23983# a_27295_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 vccd1 _1860_.CLK a_9595_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X21 vccd1 _1899_.Q a_11558_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 vccd1 _1448_.A a_12815_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 a_18427_15279# _1723_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 vssd1 a_18475_30676# _1842_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X25 _1840_.Q a_17527_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 _0952_.A2 a_26267_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1683_27791# _1767_.B _1767_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X29 vccd1 _1696_.B a_23115_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X31 a_17826_5263# _1150_.A2 a_17736_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X32 a_24278_21237# a_24110_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X33 a_24087_20394# _1525_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X34 _1191_.X a_19899_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X35 a_17385_21807# _1893_.Q a_17313_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X36 a_18459_13131# _1110_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X37 _1424_.A_N a_11711_15831# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X38 vccd1 a_17895_29941# a_17811_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X39 _0952_.A2 a_26267_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 vccd1 _1344_.B a_5271_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X43 vccd1 a_25842_24501# a_25769_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X44 vccd1 _1075_.C a_18243_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X45 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X46 vccd1 _0930_.A a_1673_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X47 a_17217_1679# _1624_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X48 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X49 vccd1 _0918_.A a_10593_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X50 vssd1 _0974_.B1 a_18940_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X51 a_16531_24349# a_15667_23983# a_16274_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X52 a_11269_16600# _1762_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X53 vccd1 a_14103_10383# _1110_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X54 a_26352_4399# a_25953_4399# a_26226_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X56 vssd1 _1126_.Y a_4447_6581# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X58 vccd1 a_2471_22869# _1771_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X59 vssd1 a_20039_5162# _1929_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X61 vccd1 a_7479_24527# _1242_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X63 a_2932_18517# _1325_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X64 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X65 vccd1 _1301_.A1 a_2778_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X67 vssd1 _1226_.A2 a_4253_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X68 vssd1 _1877_.Q a_21089_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X69 a_6682_24233# _0911_.A a_6600_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X70 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8215_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X71 vssd1 a_15243_3855# a_15411_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X72 a_26777_7663# a_25787_7663# a_26651_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X73 vssd1 _1761_.X a_3514_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 a_25214_3855# a_24775_3861# a_25129_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X76 vccd1 _0987_.Y a_11877_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X77 vccd1 a_19954_31029# a_19881_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X78 vssd1 _0906_.X a_7479_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X79 a_16083_14954# _1401_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X80 vccd1 temp1.capload\[5\].cap.A temp1.capload\[5\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X81 a_11023_5162# _1646_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X82 vccd1 a_25566_21919# a_25493_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X83 vccd1 _1102_.B a_19619_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X84 a_21235_7338# _1597_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X85 a_27337_3311# _1674_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X87 vssd1 a_9000_14967# _1298_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X88 vccd1 _1140_.C a_11711_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X91 a_23098_27613# a_22659_27247# a_23013_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X92 a_2626_12879# _1222_.B1 a_2331_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X94 a_7101_3561# _1317_.X _1800_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X97 a_19693_18377# a_18703_18005# a_19567_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X99 a_4324_31849# a_4075_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X100 a_21633_26159# _1838_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X101 a_4697_7497# a_3707_7125# a_4571_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X102 a_21108_7663# a_20709_7663# a_20982_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X103 vccd1 a_3635_24501# _2006_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X104 a_7667_22901# _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 vssd1 _1304_.B _1300_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 a_23837_21269# a_23671_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 vccd1 _1298_.A1 a_1769_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X109 a_5081_19087# _1325_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X110 vssd1 a_3635_24501# _2006_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X112 _1760_.X a_2309_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X113 vccd1 a_22806_20149# a_22733_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X114 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X116 vccd1 _1841_.CLK a_14931_32149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X117 vssd1 a_17895_29941# a_17853_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X118 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.LO a_17139_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X119 vssd1 a_10167_7093# a_10125_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X122 a_23266_11039# a_23098_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X123 a_2658_24095# a_2490_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X124 _1762_.A a_7755_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X125 a_6553_17705# _1325_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X126 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X127 vssd1 _1139_.C a_11865_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 _1029_.B1 a_14747_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X129 a_14467_28879# a_14287_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X130 a_22454_1501# a_22181_1135# a_22369_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X131 a_15189_29423# a_15023_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X132 a_17853_2057# a_16863_1685# a_17727_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X133 vccd1 a_12502_4917# a_12429_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X134 _1547_.A a_11476_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X135 a_26225_6409# a_25235_6037# a_26099_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X136 a_26183_13647# a_25401_13653# a_26099_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_9460_25847# _1332_.Y a_9602_25654# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X138 vccd1 a_4519_9991# _1172_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X139 vssd1 _1179_.C1 a_18519_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X140 a_10034_2589# a_9761_2223# a_9949_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X141 a_25030_9117# a_24757_8751# a_24945_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X142 a_23155_18909# a_22291_18543# a_22898_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
R0 temp1.capload\[10\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X143 a_20617_27791# a_20083_27797# a_20522_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X145 a_22963_1679# a_22181_1685# a_22879_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 vccd1 a_4497_7637# _1170_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X148 a_3983_28585# _1764_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X149 a_13932_21641# a_13533_21269# a_13806_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X150 vccd1 _1999_.CLK a_13275_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X151 vssd1 _1184_.A2 a_19325_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X152 a_22238_14735# _1032_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X153 a_19605_5487# a_19439_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X154 vccd1 _1010_.A a_19439_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X155 vccd1 a_18114_32117# a_18041_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X157 a_21089_18365# a_20819_17999# a_20999_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X158 vccd1 _1850_.CLK a_8307_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X159 vssd1 a_21115_11445# a_21073_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X160 vccd1 a_3083_24251# a_2999_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X161 vccd1 a_25283_14356# _1707_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X162 _1150_.B2 a_23047_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X165 a_12429_4943# a_11895_4949# a_12334_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X166 vssd1 input3.X a_5404_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 vccd1 _0958_.B a_20267_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X168 vssd1 a_26026_18655# a_25984_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X169 vssd1 a_16175_1898# _1957_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X170 a_26597_23983# a_26431_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X171 a_9949_22351# _1817_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X172 vssd1 clkbuf_0_net57.X a_2686_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X173 vccd1 _1242_.B1 a_5061_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X174 vssd1 _1075_.C a_18121_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X175 a_10839_20884# _1443_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X176 vssd1 _0932_.A a_5455_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X177 vssd1 a_23266_21919# a_23224_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X178 vccd1 a_9779_19087# _1860_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 a_12689_6721# _1065_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X181 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X182 vssd1 _0922_.Y a_8480_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X183 _0983_.X a_10147_26409# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X184 vccd1 _0964_.A a_12907_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X186 vssd1 _1154_.A1 a_23757_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X189 _1095_.C1 a_17967_12672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X190 vssd1 _1855_.CLK a_10699_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X191 a_6326_25071# _1242_.A2 a_6236_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X192 a_2382_3829# a_2214_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X194 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X195 vssd1 a_27663_21085# a_27831_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X196 _1234_.A2 a_5455_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X198 a_18409_2773# a_18243_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X200 vccd1 a_13054_25589# a_12981_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X201 _1406_.A a_18836_23555# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X202 a_15151_16733# a_14453_16367# a_14894_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X203 vssd1 _1448_.A a_12815_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X204 a_25401_12565# a_25235_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X205 a_17217_27791# _1899_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X206 vccd1 _1133_.C a_17415_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X208 vccd1 _1459_.A a_18151_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X209 a_11711_14848# _1905_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X211 _1744_.X a_19803_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X212 vssd1 a_12743_8181# a_12701_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X213 vccd1 _1156_.Y a_7834_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X214 vssd1 _0966_.A2 a_15277_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X215 a_2603_21807# _0925_.Y a_2781_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X216 vccd1 a_21235_31274# _1487_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X217 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X219 vccd1 _1924_.CLK a_26983_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X220 a_27847_10205# a_26983_9839# a_27590_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X222 a_12189_24825# _1287_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X224 vccd1 _2003_.Q a_7571_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X226 a_8822_2741# a_8654_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X227 a_3401_12925# _0917_.A a_3329_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X228 vccd1 a_17381_14337# _1034_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X229 a_19395_5162# _1667_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X233 a_24945_6575# _1605_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X234 vccd1 a_21695_19796# _1393_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X235 a_9301_7125# a_9135_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X236 a_27422_26525# a_26983_26159# a_27337_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X238 a_2873_18319# _1280_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X239 vssd1 a_26394_4511# a_26352_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X240 vssd1 _1059_.B a_17456_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X241 _1810_.A2 a_6600_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X242 vccd1 _1353_.A a_25869_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X243 a_17577_13103# _1528_.A a_17139_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X244 _1075_.C a_10938_16341# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X245 a_15207_14557# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X246 vssd1 _1821_.Q a_15616_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 vccd1 a_17359_31965# a_17527_31867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X248 vssd1 _1156_.D _1156_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X249 a_11889_6351# _1145_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X250 vccd1 _1080_.B a_18550_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X252 a_5888_31055# a_5639_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X253 a_6824_13647# _1012_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X254 vssd1 a_27215_4074# _1367_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X255 a_24294_25615# a_23855_25621# a_24209_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X256 a_4150_21263# _1310_.Y a_3759_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X258 a_25340_4233# a_24941_3861# a_25214_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X261 vccd1 _1874_.Q a_17170_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X262 a_27337_19631# _1967_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X263 vccd1 _1139_.C a_11711_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X264 a_2547_13469# a_1683_13103# a_2290_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X265 vccd1 _1850_.CLK a_12171_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X266 a_4035_30485# _1329_.X a_4262_30833# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X267 _1338_.A a_1827_32117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 a_12425_2223# a_11435_2223# a_12299_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X269 a_15795_32143# a_14931_32149# a_15538_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X270 vssd1 a_2103_31573# _1329_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 a_14287_28879# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X272 a_16192_27791# a_15943_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X273 _1394_.A a_23323_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X274 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_4324_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X275 a_2686_10383# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X276 a_21407_23261# a_20543_22895# a_21150_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X277 a_14802_7093# a_14634_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X278 a_2382_3829# a_2214_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X279 vccd1 a_22587_31867# a_22503_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X281 _1289_.A2 _1249_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X282 vssd1 _1719_.B a_22285_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X284 vssd1 a_2807_7093# a_2765_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X285 vccd1 a_13035_10383# a_13203_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X286 a_27755_11293# a_27057_10927# a_27498_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X287 a_14993_25071# _1897_.Q a_14921_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X289 vssd1 a_25455_1501# a_25623_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X291 a_13275_4765# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X292 a_4587_24501# _1261_.A1 a_4814_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X293 a_19497_18689# _1137_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X294 vccd1 _1489_.A_N a_19899_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X295 a_27479_16733# a_26781_16367# a_27222_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X296 vssd1 a_21150_7775# a_21108_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X298 a_15465_32143# a_14931_32149# a_15370_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X300 a_21143_23658# _1406_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X301 a_27054_16733# a_26615_16367# a_26969_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X302 a_6843_16911# _0930_.Y a_6588_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X303 a_21077_23261# a_20543_22895# a_20982_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X304 vssd1 _2006_.Q a_12337_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X306 _0909_.A _1255_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X307 a_6548_14191# _1332_.Y a_6245_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X308 a_13599_29588# _1469_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X309 vssd1 a_24703_21237# a_24661_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X310 vssd1 _1459_.A a_23671_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X311 a_8822_2741# a_8654_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X312 a_24639_7828# _1717_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X313 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_3063_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X314 a_3551_27791# a_2769_27797# a_3467_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 vccd1 a_22622_25589# a_22549_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X316 _1021_.X a_17691_22464# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X317 vssd1 a_7479_24527# _1242_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X318 vssd1 _1159_.X a_4800_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X319 a_11934_9295# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X320 a_11759_29098# _1429_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X321 a_27422_10205# a_27149_9839# a_27337_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X322 a_2054_32143# a_2005_32375# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X323 vccd1 a_10811_8181# a_10727_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X324 vssd1 _1764_.Y _2004_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X325 _1691_.A a_22195_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X327 a_14461_9661# _1127_.A a_14379_9408# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X328 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X329 _0981_.B _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X330 a_15883_13131# _0935_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X331 a_21725_30511# _1487_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X333 vccd1 _1841_.CLK a_14931_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X334 a_22898_18655# a_22730_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X336 vssd1 a_22063_29098# _1873_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X337 a_13261_27791# a_13084_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X339 a_24941_3861# a_24775_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X340 vssd1 _1074_.C a_13429_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X341 vccd1 a_16185_14337# _1104_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X342 _1243_.Y _1243_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X346 vccd1 _1850_.CLK a_14287_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X347 a_26225_5321# a_25235_4949# a_26099_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X349 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X350 a_20709_2223# a_20543_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X351 a_22825_2223# a_22659_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X352 a_20858_14735# _1113_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X353 vssd1 io_in[2] a_1591_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X354 a_10931_2986# _1611_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X355 vssd1 _0998_.B2 a_17604_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X356 a_4789_18319# _1267_.A1 a_4351_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X357 vccd1 _1690_.A_N a_20911_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X358 vccd1 a_21327_13866# _1986_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X359 vccd1 input3.X a_5486_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X360 _2005_.Q a_2991_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X362 _1476_.B a_18171_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X363 vccd1 a_6797_19605# _1325_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X364 a_27149_19631# a_26983_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X365 vssd1 a_19107_2767# a_19275_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X366 _1165_.A a_6467_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X367 vssd1 a_3083_24251# a_3041_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X368 a_2122_13469# a_1849_13103# a_2037_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X369 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X370 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X372 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X373 a_25198_24095# a_25030_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X376 _1685_.A_N a_21187_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X377 a_21327_13866# _1725_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X379 a_5565_22649# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X380 a_12226_16341# a_12079_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X382 a_2505_16911# _1230_.A4 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X383 a_16185_14337# _1099_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X384 _1434_.X a_9912_13763# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X385 a_22285_10749# a_22015_10383# a_22195_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X386 _1186_.X a_11987_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X387 _1414_.A a_19619_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X388 vccd1 _1855_.CLK a_12723_29973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X389 _1188_.B a_5015_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X391 a_1932_31055# a_1683_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X392 vccd1 _1775_.C1 a_1775_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X393 a_25674_22351# a_25235_22357# a_25589_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X394 vssd1 a_9195_17973# _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 a_25750_26271# a_25582_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X397 _1772_.A0 _2008_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X398 a_21123_4765# a_20341_4399# a_21039_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X399 a_10506_30511# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X400 vssd1 _0987_.Y a_14092_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X402 vccd1 a_19952_12533# _1184_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X403 a_22339_19796# _1689_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X404 vccd1 _1809_.B a_5448_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X407 a_23098_27613# a_22825_27247# a_23013_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X408 vssd1 a_26007_26525# a_26175_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X409 a_27149_9839# a_26983_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X410 a_5455_27791# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X411 vccd1 a_25198_8863# a_25125_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X412 vssd1 a_25623_5755# a_25581_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X414 vssd1 a_26267_12533# a_26225_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X415 vccd1 a_25467_28010# _1856_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X416 vccd1 a_28015_27515# a_27931_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X417 a_17029_12559# _1830_.Q a_16945_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X418 _1353_.Y _1353_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X419 a_13035_10383# a_12171_10389# a_12778_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X420 a_25769_16911# a_25235_16917# a_25674_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X421 a_22454_1679# a_22015_1685# a_22369_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X422 vccd1 a_20591_7338# _1996_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X423 vccd1 fanout24.A a_23671_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X427 a_23818_23413# a_23650_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X428 a_26781_14557# a_26247_14191# a_26686_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X429 vccd1 _1639_.X a_4351_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X430 vssd1 _1006_.X a_19991_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X431 vccd1 _1150_.B2 a_20263_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X432 vssd1 a_12539_7663# _1577_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X433 a_20315_25236# _1416_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X435 a_2485_29423# _1760_.B a_2413_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X437 vccd1 a_16911_32362# _1540_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X438 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_10876_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X439 a_25467_28010# _1453_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X440 vssd1 a_14335_25834# _1431_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X442 vssd1 _1850_.CLK a_11711_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X443 _0925_.A2 _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X444 _0984_.B1 a_10731_17483# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X445 vssd1 _1073_.A2 a_16473_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X446 vccd1 _0958_.A a_10791_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X447 vssd1 a_17647_23658# _1839_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X448 _1286_.A1 a_2623_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X449 vccd1 a_24535_11471# a_24703_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X450 _1453_.X a_10419_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X451 a_18607_26525# a_18427_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X453 vccd1 _1821_.Q a_15698_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X454 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X456 _1438_.X a_12259_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X457 _1874_.Q a_23047_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X458 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_16192_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X460 a_13485_17483# _0961_.A a_13399_17483# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X461 a_27330_28701# a_26891_28335# a_27245_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X462 _1270_.A _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X463 vccd1 _1033_.A1 a_17812_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X464 vccd1 a_9183_12180# _1571_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X466 a_23650_23439# a_23377_23445# a_23565_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X467 vssd1 a_20131_21972# _1889_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X468 a_2609_19881# _1311_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X469 a_21181_17277# a_20911_16911# a_21091_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X470 a_23351_7828# _1602_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X471 vssd1 a_24535_11471# a_24703_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X474 a_14894_16479# a_14726_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X475 _1874_.Q a_23047_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 a_17647_23658# _1418_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X478 vccd1 _1572_.B a_14467_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X480 a_15696_21263# _0965_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X481 a_19310_17973# a_19142_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X484 a_24021_25621# a_23855_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X485 vccd1 a_26927_25437# a_27095_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X486 a_17221_18793# _1826_.Q a_17139_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X487 a_25455_17821# a_24757_17455# a_25198_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X488 _0935_.X a_8307_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X490 a_9574_7119# a_9135_7125# a_9489_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X491 a_20437_28879# _1870_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X492 vccd1 a_24639_12180# _1978_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X493 vssd1 _1464_.B a_9865_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X494 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X495 vssd1 _1768_.A _1769_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X496 _1073_.A2 a_17171_16395# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X497 a_13495_2767# a_12631_2773# a_13238_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X498 vssd1 _1985_.CLK a_26799_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X499 vssd1 a_25743_1898# _1952_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X500 vccd1 a_15538_32117# a_15465_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X501 _1006_.B2 a_25623_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X502 vssd1 _1242_.A1 a_5416_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X503 a_2290_7775# a_2122_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X504 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X505 a_5908_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X506 vssd1 a_20690_28853# a_20648_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X507 vssd1 _1885_.Q a_20584_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 a_13386_9001# _1060_.C1 a_13306_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X510 vssd1 a_14563_21807# _0958_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X511 a_21048_16367# _1113_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X512 a_12938_6825# _1068_.D1 a_12689_6721# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X513 a_4101_8779# _1177_.B a_4015_8779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X515 vssd1 _1020_.A2 a_20245_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X516 a_15483_23552# _1867_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X517 a_11797_4399# a_11527_4765# a_11707_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X518 _1563_.A a_7980_9411# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X519 a_13245_19453# _1863_.Q a_13173_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X520 a_17231_19200# _1881_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X521 a_9602_15606# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X522 a_18383_3476# _1631_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X523 vccd1 _1532_.A a_5731_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X524 vccd1 a_26175_29691# a_26091_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X525 vssd1 _1325_.A2 a_7743_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X526 a_7510_24233# _1537_.B a_7428_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X527 a_6454_23145# _1282_.A2 a_6151_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X528 a_14553_6575# _0939_.A a_14471_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X529 a_17677_28879# _1469_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X531 a_20353_4221# a_20083_3855# a_20263_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X532 vssd1 _1075_.X a_15265_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X535 a_11264_31599# a_10865_31599# a_11138_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X536 _1127_.X a_20267_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X537 vccd1 _1313_.X a_6559_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X538 vssd1 a_13238_2741# a_13196_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X539 a_7159_20884# _1557_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X542 vccd1 a_8447_10004# _1563_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X543 _1198_.B2 a_13183_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X544 a_19605_31599# a_19439_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X545 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X546 a_2398_25437# a_2125_25071# a_2313_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X549 a_9503_16911# _1269_.A1 a_9921_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X550 _1130_.D1 a_19807_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X551 vssd1 _0921_.A _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X552 vccd1 a_20303_5853# a_20471_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X553 a_25030_2589# a_24591_2223# a_24945_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X554 a_27146_2589# a_26707_2223# a_27061_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X555 vccd1 a_22622_1247# a_22549_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X556 _1782_.X a_1816_11587# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X557 a_9429_15033# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X558 a_24661_21641# a_23671_21269# a_24535_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X559 a_24113_14741# a_23947_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X560 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X561 a_16232_23983# a_15833_23983# a_16106_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X564 a_14226_26819# _1484_.B a_14144_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X565 a_14833_18115# _1138_.X a_14737_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X566 vccd1 a_10202_2335# a_10129_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X567 a_8447_10004# _1563_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X568 _1314_.X a_6559_15936# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X569 a_12042_2335# a_11874_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X573 vccd1 _0958_.B a_15483_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X574 vssd1 _0994_.B2 a_15477_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X575 a_14852_30511# a_14453_30511# a_14726_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X576 vssd1 a_1823_19796# _1777_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X577 _1060_.C1 a_9595_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X578 vccd1 _1032_.C a_17231_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X579 vccd1 _0935_.X a_13551_8215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X580 _1186_.C1 a_10331_23145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X582 a_22729_5487# a_21739_5487# a_22603_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X583 a_18367_25099# _0958_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X584 a_18869_18005# a_18703_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X585 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X586 a_26007_3677# a_25309_3311# a_25750_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X587 a_21721_31599# a_21555_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X588 vssd1 a_20947_27791# a_21115_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X589 a_1849_13103# a_1683_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 a_11693_17821# a_11527_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X591 _1766_.A0 _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 vssd1 _1045_.C1 a_11953_11073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X593 vccd1 _1394_.A a_16616_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X595 a_17485_26159# a_16495_26159# a_17359_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X596 a_24535_11471# a_23671_11477# a_24278_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X597 a_19878_31965# a_19439_31599# a_19793_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X599 a_10129_2589# a_9595_2223# a_10034_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X600 vssd1 a_22879_1501# a_23047_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X601 a_25125_9117# a_24591_8751# a_25030_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X602 vccd1 _1873_.CLK a_21371_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X603 a_6607_30186# _1555_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X604 a_9865_31599# a_9595_31965# a_9775_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X605 a_10094_4943# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X606 a_5911_16617# _1265_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X607 vssd1 a_17541_15307# _1024_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X608 a_25539_2589# a_24757_2223# a_25455_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X609 a_27655_2589# a_26873_2223# a_27571_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 a_8209_15529# _1273_.A1 _1790_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X611 a_5048_14165# _1218_.B a_5271_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X612 vccd1 _1907_.CLK a_9779_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X613 vssd1 _1855_.Q a_10509_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X614 vccd1 _1133_.C a_17415_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X615 vccd1 _0964_.A a_17231_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X616 a_9786_20719# _1282_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X617 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X618 vssd1 a_17047_17455# _1405_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X619 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.A a_14370_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X620 a_12276_14025# a_11877_13653# a_12150_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X622 vssd1 _1074_.C a_11497_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X623 a_23757_29423# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X624 a_10777_27247# _1555_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X625 a_15514_21263# _1077_.D1 a_15265_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X626 a_10570_19743# a_10402_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X627 _1173_.X a_5547_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X628 _1477_.A a_12535_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X630 a_6923_16617# _1780_.B1 a_6705_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X631 _1686_.A a_23759_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X633 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12532_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X634 vccd1 _1032_.C a_21279_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X636 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A _0913_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X637 vccd1 a_26854_14303# a_26781_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X638 a_6099_27247# _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X639 a_25842_26677# a_25674_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X640 a_24393_19087# _1826_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X641 _1572_.B a_15319_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X642 vssd1 a_10827_19997# a_10995_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X643 vssd1 a_6607_30186# _1555_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X644 _1755_.A a_6831_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X646 a_21994_31965# a_21555_31599# a_21909_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X648 a_11240_16367# a_10791_16367# a_10938_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X649 a_22580_2057# a_22181_1685# a_22454_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X650 vccd1 a_8356_20407# _1233_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X651 a_24209_1679# _1628_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X652 a_16797_15307# _1021_.A a_16711_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X653 vccd1 a_13599_1300# _1947_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X654 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X655 vssd1 a_26819_7931# a_26777_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X656 a_22856_28169# a_22457_27797# a_22730_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X657 vccd1 a_25899_11195# a_25815_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X658 a_26417_25071# _1882_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X659 a_27054_16733# a_26781_16367# a_26969_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X660 a_6835_7439# _1086_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X661 vssd1 _0983_.A2 a_14920_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X662 vssd1 _1113_.C a_17385_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X663 a_4441_27247# _1764_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X666 a_12249_15279# _1433_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X667 a_17710_14441# _1031_.X a_17630_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X668 vssd1 _1043_.B a_9360_3971# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 a_3593_28169# a_2603_27797# a_3467_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X670 _1582_.A a_18560_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X671 a_16301_22057# _1530_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X672 a_27807_14735# a_27627_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X673 a_18560_8323# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X674 _1545_.A a_14467_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X675 _1141_.C a_10667_16885# a_10279_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X676 _1744_.A_N a_18151_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X677 vssd1 a_12321_22325# _1142_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X678 a_21545_18543# _0958_.A a_21463_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X679 a_15381_6575# _0939_.A a_15299_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X680 vssd1 a_27038_24095# a_26996_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X682 _1171_.Y _1165_.A a_7657_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X684 a_7993_11989# _1082_.X a_8280_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X685 a_1674_28879# clkbuf_0_temp1.i_precharge_n.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X686 _1819_.Q a_14491_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X687 vssd1 a_18151_6031# _1744_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X689 vssd1 _1249_.A2 a_2132_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X690 a_4036_14165# _1279_.A1 a_4256_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X691 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_6736_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X692 vccd1 _1316_.X a_8392_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X693 a_27443_11471# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X694 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X695 a_3329_13647# _1246_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X696 _1819_.Q a_14491_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X697 a_27801_31849# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE _1347_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X698 vccd1 a_13643_3855# _1941_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X700 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X703 vccd1 _1775_.A2 a_6682_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X704 vssd1 a_1643_21237# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X705 a_9700_7497# a_9301_7125# a_9574_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X706 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X707 a_11371_3677# a_10589_3311# a_11287_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X708 vssd1 _1191_.X a_13183_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X709 a_9460_15431# _1764_.A a_9602_15606# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X710 a_26141_4399# _1959_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 a_24110_11471# a_23837_11477# a_24025_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X712 vssd1 _1353_.Y a_8158_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X713 a_10379_25398# _1305_.B a_9920_25223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X714 a_13599_13866# _1755_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X715 a_10509_29245# a_10239_28879# a_10419_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X717 a_3681_13647# _1246_.A2 a_3553_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X718 a_15151_10205# a_14287_9839# a_14894_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X719 vssd1 a_8723_4074# _1567_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X720 a_20437_27791# _1875_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X721 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X722 vssd1 fanout37.A a_16863_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X723 vccd1 _1092_.B a_8947_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X724 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X725 vccd1 _1109_.B a_13455_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X726 _1269_.A1 a_6927_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X727 a_22549_1679# a_22015_1685# a_22454_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X728 vccd1 _0921_.B _0930_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X729 vssd1 a_2915_24349# a_3083_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X730 vssd1 a_23323_24251# a_23281_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X731 a_3225_20719# _1269_.A1 a_2787_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X732 vssd1 _1154_.C1 a_22073_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X734 a_13437_25993# a_12447_25621# a_13311_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X735 vssd1 a_10287_2986# _1659_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X736 _1051_.A1 a_8051_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X737 a_20395_30877# a_19531_30511# a_20138_30623# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X738 vccd1 a_8548_23413# _1329_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X739 vccd1 _0973_.B a_21827_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X740 a_6611_29111# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X741 vccd1 _0964_.A a_13643_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X742 _1709_.X a_22563_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X743 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X745 vccd1 _1006_.B2 a_27347_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X747 a_24845_2057# a_23855_1685# a_24719_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X748 a_25156_2223# a_24757_2223# a_25030_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X749 a_27272_2223# a_26873_2223# a_27146_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X750 _1221_.A _1123_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X751 a_26229_25071# a_26063_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X752 a_3247_13967# _1246_.B2 _1247_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.105625 ps=0.975 w=0.65 l=0.15
X753 a_23105_22351# _1828_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X757 vssd1 _1090_.C a_12325_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X758 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_1683_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X759 a_27847_27613# a_27149_27247# a_27590_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X760 a_23005_27081# a_22015_26709# a_22879_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X761 vccd1 a_20303_31965# a_20471_31867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X763 a_20065_30877# a_19531_30511# a_19970_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X764 _1257_.X a_3087_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X766 vccd1 a_6073_25045# _1344_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X767 a_4847_25437# a_3983_25071# a_4590_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X768 a_2009_21583# _1308_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X770 a_17541_15307# _0964_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X772 _1976_.Q a_25439_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X773 a_16514_14441# _1097_.X a_16434_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X774 a_10227_11471# _1198_.A2 _1122_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X775 a_1945_1135# _1808_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X776 vssd1 a_26007_10205# a_26175_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X777 vssd1 a_27831_22075# a_27789_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X778 vssd1 a_11287_3677# a_11455_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X779 _1611_.X a_9360_3971# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X780 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X782 a_11865_7663# _1148_.B a_11793_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X783 vccd1 _1010_.A a_12171_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X784 vssd1 _0985_.A a_15575_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 _1693_.A a_23667_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X786 temp1.capload\[13\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X787 a_15971_29789# a_15189_29423# a_15887_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X788 a_3217_14191# _1249_.A2 a_3145_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X789 a_17930_28853# a_17762_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X790 vccd1 _0930_.B _1326_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X791 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X792 a_20709_7663# a_20543_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X793 _1010_.A a_13551_8215# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X794 a_14379_9408# _1030_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X795 a_2198_9269# a_2030_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X796 a_17630_25321# _1537_.B a_17548_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X797 vccd1 a_27847_5853# a_28015_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X798 vccd1 _1876_.CLK a_23855_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X800 vssd1 a_22063_8426# _1916_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X802 a_14407_24527# a_13625_24533# a_14323_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X803 a_23013_27247# _1893_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X804 a_27627_14735# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X805 a_9186_13255# _1187_.X a_9323_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X806 vccd1 temp1.capload\[0\].cap.A temp1.capload\[0\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X808 _1886_.Q a_27923_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X809 vssd1 a_8971_1653# a_8929_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X810 vssd1 a_16911_32362# _1540_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X811 a_8785_15974# _0956_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X812 a_10765_19407# _0921_.A a_10515_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X813 vccd1 _1286_.A1 a_7657_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X814 a_22322_12559# _1153_.X a_22073_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X816 a_26735_4765# a_25953_4399# a_26651_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X817 vccd1 _0963_.B a_16863_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X818 vssd1 a_25842_20149# a_25800_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X819 vccd1 _1841_.CLK a_17139_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X820 a_27364_15279# a_26965_15279# a_27238_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X821 a_17366_6351# _0998_.A2 a_17276_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X822 vssd1 _1849_.CLK a_20543_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X823 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X824 _1684_.A a_22747_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X825 a_25030_17821# a_24757_17455# a_24945_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X826 _1193_.X a_16127_16617# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X827 a_16749_2223# a_15759_2223# a_16623_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X828 vccd1 a_20046_1247# a_19973_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X829 _1660_.X a_12351_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X830 vssd1 _1896_.CLK a_19807_32149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X831 vssd1 _1823_.CLK a_23211_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X833 vssd1 a_20303_5853# a_20471_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X834 a_25455_6941# a_24757_6575# a_25198_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X835 vssd1 a_2382_4511# a_2340_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X836 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X837 a_5710_2589# a_5271_2223# a_5625_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X838 vccd1 _1127_.A a_15483_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X839 _1680_.A a_22563_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X840 a_2490_24349# a_2217_23983# a_2405_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X841 _1887_.CLK a_23395_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X842 vssd1 _1768_.A _0951_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X843 vssd1 _1116_.X a_14287_13353# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X844 vccd1 _1127_.A a_18427_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X845 vccd1 a_25623_24251# a_25539_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X846 a_3410_2767# a_3137_2773# a_3325_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X847 a_25401_26709# a_25235_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X848 a_6703_26133# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X849 vccd1 a_26099_13647# a_26267_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X850 a_16290_4399# a_16113_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X851 _1226_.A1 a_1775_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X852 vssd1 a_17359_26525# a_17527_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X854 a_4590_1653# a_4422_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X855 a_19789_28335# a_19623_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X856 a_10677_22895# _1859_.Q a_10331_23145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X858 vccd1 a_18151_19631# _1032_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X859 vccd1 _0956_.C a_7479_17277# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X860 a_23289_3855# _1991_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X861 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X862 vssd1 _1818_.Q a_8945_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X864 vssd1 a_12467_2491# a_12425_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X865 a_7189_3855# _1365_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X866 vssd1 a_26099_13647# a_26267_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X867 vssd1 a_17647_2388# _1944_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X868 fanout24.A a_22935_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X869 clkbuf_0_net57.A temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X870 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X871 vccd1 _1887_.CLK a_26983_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X872 a_10769_2057# a_9779_1685# a_10643_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X873 vccd1 a_10167_5755# a_10083_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X874 vssd1 _0916_.A a_3401_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X875 a_12295_20747# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X876 vssd1 _1874_.Q a_17088_26819# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X878 a_10034_29789# a_9761_29423# a_9949_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X880 vssd1 _2006_.Q a_12299_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X881 a_7383_29967# a_7203_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X882 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X883 vccd1 _1828_.Q a_16986_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X884 vccd1 _1590_.A_N a_17139_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X885 a_4422_25437# a_4149_25071# a_4337_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X887 a_23013_10927# _1716_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X888 a_2695_17999# _1281_.B1 a_2873_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
D0 vssd1 _1652_.X sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X889 a_27253_5263# _1159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X890 _1147_.C1 a_16863_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X891 a_18581_15279# _1723_.B a_18509_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X894 a_4495_11989# _1301_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X895 a_25589_12559# _1965_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X896 a_12609_23983# _1451_.B a_12171_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X897 vccd1 a_1644_18517# _1300_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X898 a_10133_1679# _1616_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X899 a_14549_7119# _1759_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X900 a_12318_29535# a_12150_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X901 vccd1 a_9742_31029# a_9669_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X902 vssd1 _1762_.Y _2003_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X903 a_1757_9301# a_1591_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X905 vccd1 a_13663_2741# a_13579_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X906 a_4897_15823# _1277_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X907 a_20303_29789# a_19605_29423# a_20046_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X908 vccd1 a_24243_16885# a_24159_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X909 vccd1 a_1829_16341# _1311_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X910 vssd1 fanout24.A a_22659_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X911 vssd1 a_13875_23658# _1840_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X912 a_23377_23445# a_23211_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X913 vccd1 _1900_.Q a_9223_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X914 a_25355_17999# a_24573_18005# a_25271_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X915 a_12337_24233# _1902_.Q a_12253_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X916 vssd1 _1039_.B a_7704_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X917 vccd1 _2023_.CLK a_1683_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X919 a_21733_12015# a_21463_12381# a_21643_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X920 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_6559_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X921 a_19793_29423# _1471_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X923 a_2129_4943# _2021_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X925 vssd1 _0903_.C _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X926 temp1.capload\[5\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X927 a_23021_15279# a_22751_15645# a_22931_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X928 a_4847_1679# a_4149_1685# a_4590_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X929 vssd1 _1007_.A1 a_20905_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X930 vccd1 _1329_.S a_7006_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X931 vccd1 _1474_.B a_13455_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X932 a_19878_31965# a_19605_31599# a_19793_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X933 a_5541_3311# a_5349_3616# _2021_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X934 vccd1 _1165_.A _1210_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X935 vssd1 _1020_.A2 a_18957_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X936 a_22438_29535# a_22270_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X937 vccd1 _1880_.CLK a_23947_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X938 vccd1 a_8286_27247# a_8392_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X939 _1650_.X a_4531_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X940 a_27421_17455# a_26431_17455# a_27295_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X941 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X942 vssd1 _1298_.A1 a_6743_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.12675 ps=1.04 w=0.65 l=0.15
X943 a_9580_22057# _0921_.B a_9496_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X944 vccd1 _1985_.CLK a_24591_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X945 vssd1 a_22695_29789# a_22863_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X946 a_26225_23817# a_25235_23445# a_26099_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X947 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X948 vccd1 a_22081_13621# _1006_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X949 vccd1 _1133_.C a_17539_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X950 a_14726_16733# a_14453_16367# a_14641_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X951 _1490_.A a_18607_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X952 _1294_.X a_5203_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X953 vssd1 a_7561_22941# a_7667_22901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X954 a_10129_22351# a_9595_22357# a_10034_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X955 vccd1 a_20138_30623# a_20065_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X956 a_18003_29789# a_17305_29423# a_17746_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X957 _1090_.C a_9282_16341# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X958 _1277_.A _1217_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X959 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_7606_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X960 a_22015_16911# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X961 _1184_.B1 a_17999_16395# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X962 vssd1 a_25198_2335# a_25156_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X963 a_10344_20495# a_9963_20175# _1232_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X964 a_2214_3677# a_1775_3311# a_2129_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X965 vssd1 a_27314_2335# a_27272_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X966 vssd1 a_2639_7119# a_2807_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X967 vssd1 _1133_.C a_14809_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X969 _0930_.A a_6559_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X970 a_24757_31599# a_24591_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X971 a_22580_25993# a_22181_25621# a_22454_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X972 _1583_.X a_18607_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X973 a_1657_10901# _1263_.A a_1910_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X974 a_18129_29423# a_17139_29423# a_18003_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X975 vssd1 _1884_.Q a_21412_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X976 a_4590_25183# a_4422_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X977 a_21994_31965# a_21721_31599# a_21909_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X978 vssd1 _1150_.B2 a_18064_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X979 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_5888_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X980 vssd1 _1760_.X a_27167_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X982 a_19480_15529# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X984 vccd1 _1374_.A_N a_15299_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X985 a_14073_19453# _1900_.Q a_14001_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X986 vssd1 _2006_.Q a_11141_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X987 a_10594_14735# _1762_.A a_10397_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X988 a_26099_13647# a_25235_13653# a_25842_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X989 a_6747_13967# _1766_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X991 a_23197_29967# _1843_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X992 a_21787_8916# _1590_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X993 a_16382_25071# a_16205_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X994 _1366_.X a_4760_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X995 _1242_.B1 a_7479_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X997 a_1766_26159# clkbuf_1_1__f__0380_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X998 vssd1 _0963_.B a_16245_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X999 a_2698_23217# a_2649_23047# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X1000 _1230_.B1 _1249_.A2 a_5241_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X1001 vccd1 _1764_.A a_3983_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1003 a_25340_16367# a_24941_16367# a_25214_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1005 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1006 a_6135_2589# a_5271_2223# a_5878_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1007 _1049_.C1 a_14287_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1009 a_25030_27613# a_24591_27247# a_24945_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1010 vccd1 _2009_.CLK a_2603_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1011 a_7649_15279# a_7472_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1012 vssd1 a_15503_2741# a_15461_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1013 _1441_.A a_14467_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1014 a_9879_12675# a_9687_12919# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1015 _1250_.B2 _1311_.B1 a_5187_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1016 vssd1 a_2198_9269# a_2156_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1017 _1486_.X a_13455_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1018 a_24757_15279# a_24591_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1019 a_17319_5853# a_17139_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1021 vccd1 _1056_.X a_12973_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1022 _1051_.A1 a_8051_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1025 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1026 vccd1 a_3467_27791# a_3635_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1028 a_18957_17231# _1967_.Q a_18519_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1032 a_5836_2223# a_5437_2223# a_5710_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1033 vssd1 _1113_.C a_19961_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1034 a_1814_11177# _1170_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X1036 vccd1 _1873_.CLK a_21831_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1037 _1884_.Q a_26267_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1039 a_15017_10499# _0999_.X a_14921_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1040 a_3210_27765# a_3042_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1041 vssd1 _1999_.CLK a_12631_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1042 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_10968_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1044 a_7641_1135# a_6651_1135# a_7515_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1045 a_2405_27247# _2003_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1046 vssd1 _1763_.A2 a_2601_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1047 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1048 a_12460_15279# a_12061_15279# a_12334_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1049 _1574_.X a_19480_15529# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1051 vccd1 _1985_.CLK a_25235_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1052 vccd1 _1054_.C a_18151_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1053 a_7883_4765# a_7185_4399# a_7626_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1054 a_18371_31055# a_17673_31061# a_18114_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1055 _1884_.Q a_26267_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1056 a_21491_8029# a_20709_7663# a_21407_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1057 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1058 a_17221_13353# _1070_.A2 a_17305_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1060 vssd1 _1883_.Q a_20216_22467# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1061 vssd1 _1068_.A1 a_14328_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1062 vccd1 _1374_.A_N a_6835_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1065 vssd1 _1022_.X a_17013_19777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X1066 _1633_.X a_17319_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1067 vccd1 a_2327_5487# _1532_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1068 vccd1 a_23047_2741# a_22963_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1069 vccd1 _0963_.B a_14287_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1070 a_2405_9839# a_2228_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1072 a_6747_13967# _1175_.B2 a_6610_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X1073 vssd1 a_2290_13215# a_2248_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1074 a_16945_10749# _1110_.A a_16863_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1075 a_4059_15431# _0930_.B a_4209_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1076 _1459_.A a_12815_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1077 a_27517_5853# a_26983_5487# a_27422_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1078 vssd1 _1083_.A a_4760_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1079 vssd1 _1896_.CLK a_19439_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1081 vccd1 a_20487_28701# a_20655_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1082 a_17845_8573# _1040_.B a_17773_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1084 a_2455_8207# a_1757_8213# a_2198_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1085 a_26873_8751# a_26707_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1086 a_24757_8751# a_24591_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1087 _0909_.A _1234_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1088 temp1.capload\[2\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1089 vssd1 a_27847_5853# a_28015_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 _1840_.Q a_17527_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1092 a_17359_31965# a_16661_31599# a_17102_31711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1093 a_15616_18115# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1094 _1158_.X a_9879_12675# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X1095 vccd1 _1775_.A2 a_8213_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1099 a_2309_29789# _1775_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X1101 vccd1 a_20601_15797# _1082_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1102 vssd1 _1807_.Y a_5357_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X1103 vssd1 _1196_.C a_14287_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1104 a_27379_17821# a_26597_17455# a_27295_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1105 vccd1 a_21235_25834# _1513_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1106 vccd1 a_2195_12533# _1223_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1107 a_8855_8207# a_8675_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1109 a_6457_12265# _1314_.X _1793_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1110 vssd1 _1317_.X a_5573_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1111 _1621_.X a_14283_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1112 vccd1 a_4739_7093# a_4655_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1114 a_12978_27791# a_12801_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1115 vssd1 a_24243_23413# a_24201_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1116 vccd1 a_6835_18543# _1768_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1117 a_15917_5461# _0997_.X a_16074_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1118 vccd1 fanout24.A a_22659_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1120 vssd1 _1041_.A1 a_20997_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1121 vssd1 _1823_.CLK a_22291_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1122 vssd1 a_23627_6740# _1593_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1123 a_10160_28169# a_9761_27797# a_10034_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1124 a_10007_20719# _1304_.B a_9644_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1125 a_25221_10927# _1680_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1127 vccd1 _0965_.A2 a_18785_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1129 a_12873_14337# _1035_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X1130 a_17029_29973# a_16863_29973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1132 a_10413_23145# _1817_.Q a_10331_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1133 vccd1 _1255_.A1 a_8027_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1134 vccd1 _0930_.B a_6588_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1135 a_9735_9514# _1759_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1136 _1126_.Y _1125_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X1137 a_6363_10927# _1304_.B _1797_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1138 a_10218_29967# a_9779_29973# a_10133_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1139 _1822_.Q a_23231_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1140 vccd1 _1195_.A2 a_16986_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1141 vccd1 _1207_.B1_N _1226_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1142 vccd1 temp1.capload\[4\].cap.A temp1.capload\[4\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1143 vssd1 a_11455_27515# a_11413_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1144 vssd1 _1838_.Q a_16904_22467# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1145 a_2129_3855# _1796_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1146 a_20349_10927# _0952_.A1 a_20267_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1148 vssd1 a_23903_26922# _1342_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1149 a_25581_23983# a_24591_23983# a_25455_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1150 io_out[5] a_3759_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1151 vccd1 _1110_.A a_18519_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1152 _1822_.Q a_23231_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1154 vssd1 clkbuf_1_1__f__0380_.A a_1766_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1156 vccd1 _1723_.A_N a_27167_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1157 a_14637_2773# a_14471_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1158 vccd1 _1902_.Q a_7510_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1160 a_23266_2335# a_23098_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1161 a_17861_1135# _1956_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1162 vssd1 a_22771_5755# a_22729_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1163 _1140_.X a_10791_23552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1164 a_16097_10749# _1102_.B a_16025_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1165 vssd1 _1775_.C1 _2004_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1166 vssd1 a_9644_20871# _1335_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 a_2340_3311# a_1941_3311# a_2214_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1168 a_18078_9295# _1110_.X a_17998_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1169 a_23266_21919# a_23098_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1170 a_4533_18793# _1232_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1171 vssd1 _1234_.A1 _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1173 a_23742_4399# a_23565_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1174 a_20046_29535# a_19878_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1175 vccd1 _1841_.Q a_15939_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1176 a_5547_7913# _1210_.B a_5629_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1177 a_3467_27791# a_2603_27797# a_3210_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1178 a_21150_2335# a_20982_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1179 a_2639_4943# a_1775_4949# a_2382_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1180 a_13805_11471# _1156_.C a_13999_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1181 vccd1 _0963_.B a_11159_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1182 a_23837_10389# a_23671_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1185 a_13257_31061# a_13091_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1186 a_26183_24527# a_25401_24533# a_26099_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1189 vssd1 a_2639_6031# a_2807_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 a_21718_26525# a_21279_26159# a_21633_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1192 a_24113_28885# a_23947_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1193 vccd1 _0909_.A a_3801_28981# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1194 vccd1 _1863_.Q a_14226_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1195 vssd1 a_25566_8181# a_25524_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1197 a_25582_29789# a_25309_29423# a_25497_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1198 a_19793_26159# _1542_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1199 vssd1 a_27295_17821# a_27463_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 a_9775_31965# a_9595_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1201 a_4293_15529# _1289_.A2 a_4209_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1202 vssd1 clkbuf_0_net57.A a_2594_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1204 vccd1 _1849_.CLK a_16127_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1205 a_3137_27791# a_2603_27797# a_3042_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1206 a_18560_7913# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1207 a_4036_14165# _1325_.A2 a_4428_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1208 _1265_.A2 _1250_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1209 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1210 a_2566_25183# a_2398_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1211 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1213 a_17746_29535# a_17578_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1214 vssd1 fanout20.X a_22015_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1215 vccd1 _1532_.A a_12815_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1216 _1030_.B a_14307_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1217 vccd1 _1153_.A a_19439_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1218 a_7749_9839# _1156_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1219 vssd1 a_5015_25339# a_4973_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1220 a_21042_16617# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1221 vssd1 a_11023_7338# _1649_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1222 a_19970_30877# a_19697_30511# a_19885_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1223 a_16904_25731# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1224 vssd1 a_14231_21263# a_14399_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1225 a_22825_4949# a_22659_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1226 vccd1 temp1.capload\[11\].cap.A temp1.capload\[11\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1227 vccd1 fanout33.A a_14931_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1228 a_15607_12043# _0958_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1229 vccd1 a_25455_5853# a_25623_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1230 a_10506_30511# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1231 a_13948_14735# _0987_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1232 a_11023_5162# _1646_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1233 _1119_.A1 a_22771_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1234 a_2036_32509# a_2005_32375# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X1235 vccd1 a_17470_27765# a_17397_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1236 a_18512_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1237 a_15538_31029# a_15370_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1240 a_22195_4765# a_22015_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1241 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1242 a_25401_23445# a_25235_23445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1243 vccd1 a_11693_17821# _1113_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1244 vssd1 a_5878_2335# a_5836_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1246 a_8855_22351# a_8675_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1248 vssd1 a_13479_25589# a_13437_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1250 a_2103_31573# _1329_.A0 a_2312_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X1251 a_4805_4175# _1801_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1252 vccd1 _1982_.CLK a_23246_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1253 vssd1 _1054_.C a_18151_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1254 a_17811_1679# a_17029_1685# a_17727_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1255 _1109_.B a_16791_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1256 a_20387_26525# a_19605_26159# a_20303_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1257 vccd1 _2004_.Q a_10791_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1258 vssd1 _1188_.B a_4621_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1262 a_23147_20175# a_22365_20181# a_23063_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1263 vccd1 a_6559_9295# _0930_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1265 vccd1 a_6927_17999# _1764_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1266 vssd1 a_4341_6621# a_4447_6581# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1267 a_15370_31055# a_15097_31061# a_15285_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1268 vssd1 a_9871_24527# _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1269 vssd1 a_24087_20394# _1525_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1270 vccd1 a_3945_4917# _2020_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1272 _1222_.A1 a_5303_9633# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1274 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1275 a_2639_3855# a_1941_3861# a_2382_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1276 vssd1 _1113_.C a_18949_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1277 _1670_.A a_22195_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1278 a_7656_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1280 _1217_.A2 a_1775_12265# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1281 a_17967_4765# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1282 _1103_.D1 a_15943_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1283 vccd1 _1721_.B a_22379_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1284 a_15151_30877# a_14287_30511# a_14894_30623# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1285 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11888_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1286 vssd1 _0921_.B _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 a_24087_20394# _1525_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1288 vssd1 _1194_.B2 a_12625_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1289 a_8177_12533# _1052_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1290 a_9574_7119# a_9301_7125# a_9489_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1291 a_13330_29941# a_13162_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1292 vssd1 _1083_.A a_9176_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1293 _1137_.X a_18519_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1294 _1187_.X a_15299_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X1295 vccd1 a_22879_31055# a_23047_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1296 vssd1 _1019_.B a_17409_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1297 vssd1 a_4259_13103# _1780_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1298 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1300 a_12778_10357# a_12610_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1301 vssd1 a_22879_31055# a_23047_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1302 a_1735_29941# _1775_.C1 a_2291_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1303 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1304 vccd1 _1353_.A a_27801_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1305 a_11711_21263# _0984_.B1 a_11793_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1306 vccd1 a_19487_2388# _1993_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1307 _1041_.A1 a_26267_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1308 _1773_.Y _1773_.B a_1775_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1309 a_13162_29967# a_12889_29973# a_13077_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1310 a_16014_3677# a_15575_3311# a_15929_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1311 vccd1 a_22935_10383# fanout24.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1312 _1769_.B1 _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1314 a_25455_21085# a_24591_20719# a_25198_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1315 a_7258_1247# a_7090_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1316 vssd1 _1968_.Q a_22285_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1317 a_2030_6941# a_1757_6575# a_1945_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1318 a_8109_14796# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1320 vssd1 _1924_.CLK a_22659_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1321 _1833_.Q a_23047_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1322 a_19310_17973# a_19142_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1323 a_23903_1300# _1736_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1324 a_9786_21046# _1282_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1325 a_14231_21263# a_13367_21269# a_13974_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1326 vssd1 a_7571_20175# _0956_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1327 vssd1 _2023_.CLK a_1775_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1328 a_12113_20495# a_11711_20175# a_12027_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X1329 a_12500_15797# _1070_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X1330 vccd1 a_22155_23658# _1691_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1331 a_14733_4943# _1749_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1332 vssd1 _0987_.Y a_10596_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1333 _1086_.Y _1086_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1334 vssd1 a_20303_26525# a_20471_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1335 vssd1 _1053_.A a_13183_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1336 vccd1 a_17841_17601# _1049_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1337 a_24945_7119# _1599_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1338 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1339 a_4547_30833# _1353_.A a_4035_30485# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X1340 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_10506_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1341 vccd1 a_16863_23439# fanout33.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1342 a_27422_19997# a_26983_19631# a_27337_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1343 _1833_.Q a_23047_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1344 vccd1 a_4035_20693# _1268_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X1345 vccd1 a_11907_20175# a_12027_20495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1346 vccd1 _1079_.B a_21643_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1348 vccd1 a_12299_2589# a_12467_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1350 vccd1 _1033_.A2 a_20065_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X1351 a_2455_1501# a_1757_1135# a_2198_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1352 vssd1 a_22879_1679# a_23047_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1354 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1356 vssd1 _1170_.A3 a_3217_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1357 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9135_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1358 vssd1 a_21831_25071# _1876_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1359 vccd1 _1690_.A_N a_22843_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1360 a_23211_16733# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1363 a_24639_23060# _1517_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1364 a_19142_17999# a_18869_18005# a_19057_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1365 _1147_.X a_17139_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1366 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_6736_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1367 a_7479_28585# _1273_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1368 _1056_.D1 a_13367_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1370 vssd1 _1440_.B a_14557_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1371 vccd1 _1442_.A a_9442_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1372 a_9921_16911# _1269_.A1 a_9503_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1373 vssd1 _0921_.B a_7481_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1374 a_2686_15823# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1375 a_7295_6031# _1173_.X a_7295_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X1376 a_15795_31055# a_15097_31061# a_15538_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1377 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1379 _1313_.A a_2623_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1380 a_10212_32143# a_9963_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1382 _1738_.X a_20539_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1383 vssd1 a_12042_25183# a_12000_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1385 vssd1 _1219_.A2 a_2850_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
X1386 vccd1 _1153_.A a_19439_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1387 vccd1 _1263_.A a_3063_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1388 a_14373_32463# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 vccd1 _0918_.A a_6651_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1391 a_17444_19881# _1021_.X a_17342_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1392 _1311_.B1 a_4899_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1393 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1394 a_12528_10927# _1572_.B a_11953_11073# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X1396 vssd1 _1038_.A1 a_9681_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1397 vssd1 a_25455_24349# a_25623_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1398 a_27061_2223# _1731_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1399 vssd1 a_16791_2491# a_16749_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1400 vssd1 _1306_.A2 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1402 vccd1 _1489_.A_N a_18427_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1404 a_20701_14709# _0952_.A1 a_20954_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1405 vccd1 a_7993_11989# _1086_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X1406 vccd1 a_23443_31764# _1475_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1407 vccd1 a_6303_2491# a_6219_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1409 vccd1 a_26819_7931# a_26735_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1410 a_12318_11445# a_12150_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1412 vssd1 a_25283_14356# _1707_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1415 vssd1 _1277_.B a_3217_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1417 vccd1 _2004_.Q a_11527_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1418 a_19789_28335# a_19623_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1419 a_27337_12015# _1978_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1421 vccd1 _1217_.A3 a_4709_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1422 a_5878_2335# a_5710_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1423 a_4069_5737# _1801_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1424 vssd1 a_19487_21972# _1828_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1425 a_22285_21629# a_22015_21263# a_22195_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1426 a_24757_2223# a_24591_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1427 a_26873_2223# a_26707_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1428 vccd1 _1941_.CLK a_16863_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1429 vccd1 a_2623_8181# _1242_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1430 a_11685_9813# _0991_.X a_11842_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1431 vssd1 _1887_.CLK a_26983_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1432 a_21787_8916# _1590_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1434 _1442_.A a_15319_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1435 a_5503_4074# io_in[5] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1436 a_9999_5853# a_9301_5487# a_9742_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1437 a_10948_28585# a_10699_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1438 a_23607_9117# a_22825_8751# a_23523_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1439 a_10459_29789# a_9761_29423# a_10202_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1440 a_5871_1898# _1368_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1441 vssd1 a_25198_31711# a_25156_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1442 vccd1 a_20471_29691# a_20387_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1443 a_17132_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1444 vssd1 _0951_.B a_19593_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1445 _1464_.X a_9775_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1446 vssd1 _1112_.A1 a_21089_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1447 a_10034_29789# a_9595_29423# a_9949_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1448 a_10593_22057# _0921_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1449 a_19487_21972# _1395_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1450 _0983_.B1 a_13399_17483# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1451 _1722_.A a_22379_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1453 vssd1 a_26267_23413# a_26225_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1454 vssd1 a_24087_13866# _1967_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1455 _2005_.Q a_2991_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1456 vccd1 _1877_.Q a_20999_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1457 vssd1 fanout21.X a_24591_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1458 _1072_.X a_11711_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1459 a_4441_27247# _1242_.A1 _2004_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1460 a_6651_23439# _0921_.Y _0922_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1461 a_24535_11471# a_23837_11477# a_24278_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1463 vssd1 a_11731_31867# a_11689_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1464 a_6743_27791# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1465 a_25566_21919# a_25398_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1466 a_27238_22173# a_26965_21807# a_27153_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1467 a_20079_19087# a_19899_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1468 vssd1 a_16439_3677# a_16607_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1469 a_14557_14191# a_14287_14557# a_14467_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1470 a_7993_11989# _1084_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X1471 vssd1 _1353_.B a_12482_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1472 a_23523_27613# a_22825_27247# a_23266_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1473 a_24087_13866# _1686_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1475 a_15097_32149# a_14931_32149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1476 a_1674_28879# clkbuf_0_temp1.i_precharge_n.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1478 _1564_.X a_7843_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1480 a_15115_14851# _1104_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1481 a_5356_13109# a_5169_13149# a_5269_13367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1482 vssd1 _1041_.C1 a_15725_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X1484 vssd1 a_16699_24251# a_16657_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1485 vccd1 a_23671_15279# _1690_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1486 _1775_.A2 a_2327_20183# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1487 vssd1 a_21695_19796# _1393_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1488 vssd1 _1177_.C a_3181_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1489 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1490 _1793_.Y a_8109_14796# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X1491 vssd1 _0930_.A a_9879_12675# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1492 a_4896_3855# _1800_.A2 _2019_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1494 vccd1 _1780_.B1 a_4613_3916# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X1496 vssd1 a_21235_31274# _1487_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1497 a_12061_15279# a_11895_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1498 _1868_.Q a_15963_32117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1499 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1501 a_11877_11477# a_11711_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1502 a_2639_28701# a_1941_28335# a_2382_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1503 vccd1 a_26007_26525# a_26175_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1504 a_2658_24095# a_2490_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1505 vssd1 a_1735_29941# _1775_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X1506 vssd1 _1075_.C a_18581_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1507 a_25582_3677# a_25143_3311# a_25497_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1508 vccd1 _1153_.A a_18243_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1509 a_24757_7125# a_24591_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1510 a_2214_28701# a_1775_28335# a_2129_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1511 a_20267_10927# _0973_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1513 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1514 a_25674_6031# a_25401_6037# a_25589_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1515 _1459_.A a_12815_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1516 _1868_.Q a_15963_32117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1518 a_25455_28701# a_24757_28335# a_25198_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1520 a_20930_15823# _1081_.C1 a_20850_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1522 vssd1 a_25455_5853# a_25623_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1524 a_9644_20871# _1304_.B a_9786_21046# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1525 a_13349_20175# _0913_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1526 _1119_.A1 a_22771_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 vssd1 a_20138_30623# a_20096_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1528 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A _1274_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1529 _0988_.X a_14319_7691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1530 vssd1 _2023_.CLK a_1591_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1531 a_16140_3311# a_15741_3311# a_16014_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1532 vccd1 _1590_.A_N a_9503_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1534 vccd1 a_2715_7931# _1261_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1535 _1127_.A a_14839_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1536 vccd1 temp1.capload\[1\].cap.A temp1.capload\[1\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 vccd1 _1976_.Q a_22931_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1538 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_12440_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1539 vssd1 a_20499_23658# _1835_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1541 a_8548_23413# a_8399_23492# a_8998_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1542 _1269_.A1 a_6927_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1543 a_9674_17705# _1762_.A a_9477_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1544 a_10791_13469# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1546 a_23818_16885# a_23650_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1547 a_22181_24533# a_22015_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1548 a_14335_2388# _1619_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1549 vssd1 _0913_.Y a_3435_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1555 a_24278_10357# a_24110_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1556 vccd1 a_3635_27765# _2004_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1557 _1238_.X a_7667_22901# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1560 a_9945_1685# a_9779_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1562 _1153_.A a_18059_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1563 _2003_.D _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1564 a_22603_6941# a_21905_6575# a_22346_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1566 _1410_.A a_19388_22467# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1567 a_4526_22057# _1308_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1568 a_21361_14191# _1153_.A a_21279_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1569 a_10428_5263# _0988_.X a_9937_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X1570 _1304_.B a_2807_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1571 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1572 vssd1 a_12035_2986# _1934_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1573 vccd1 _1008_.A a_15089_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1574 vssd1 a_1591_15279# _0929_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 vssd1 _1086_.A a_6467_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1579 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_10212_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1580 a_25455_31965# a_24591_31599# a_25198_31711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1581 vccd1 a_8447_20884# _1433_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1582 a_10094_4943# _1140_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X1583 a_23650_16911# a_23377_16917# a_23565_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1584 vssd1 _0989_.B2 a_9773_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1585 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1586 a_17428_18377# a_17029_18005# a_17302_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1588 _1329_.S a_8548_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1590 vccd1 a_2807_4917# a_2723_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1592 a_22856_23983# a_22457_23983# a_22730_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1593 vccd1 _1842_.Q a_18239_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1596 _1067_.B a_8143_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1597 _0974_.B1 a_20267_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1599 vssd1 _0921_.A a_9963_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
X1600 a_2455_2589# a_1591_2223# a_2198_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1601 a_10515_6575# _0988_.X a_10693_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1602 a_16064_11471# _1179_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1603 a_14726_10205# a_14287_9839# a_14641_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1604 vssd1 _1897_.Q a_13408_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1605 _0989_.B2 a_9247_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1606 a_13629_1679# _1659_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1607 vssd1 _1183_.A2 a_22653_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1608 a_21886_26271# a_21718_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1609 _1116_.C1 a_13643_22464# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1610 a_8447_20884# _1433_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1611 vccd1 a_3983_17455# _0921_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1612 a_14453_30511# a_14287_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1613 a_2962_14735# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1614 a_24757_15279# a_24591_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1615 a_20303_31965# a_19605_31599# a_20046_31711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1617 a_25581_8751# a_24591_8751# a_25455_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1618 a_25589_20175# _1970_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1619 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1620 a_10202_27765# a_10034_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1621 vccd1 _0963_.B a_12907_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1622 a_8756_16189# a_8307_15823# a_8454_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1623 vccd1 a_7896_11079# _1162_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1624 vssd1 _1132_.C a_14073_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1625 a_7975_2589# a_7277_2223# a_7718_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1626 vccd1 a_2198_6687# a_2125_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1627 vssd1 _1071_.B1 a_13183_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1628 a_15633_19061# _1020_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X1629 vccd1 a_25271_17999# a_25439_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1630 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1631 vccd1 _1308_.B a_1779_22453# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1633 a_8701_25953# _0911_.A a_8615_25953# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1634 a_21077_8029# a_20543_7663# a_20982_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1636 a_8624_17027# _1313_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1638 _1789_.A1 _1261_.A1 a_5909_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1639 vccd1 _1055_.C a_14563_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1640 a_2966_19131# _0930_.Y a_2965_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X1642 vccd1 a_4036_14165# _1281_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1644 a_9032_11471# _1104_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X1645 a_15887_29789# a_15023_29423# a_15630_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1646 vccd1 a_10883_21271# _1132_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1647 a_22745_32463# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1648 a_10034_27791# a_9761_27797# a_9949_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1649 a_27517_26525# a_26983_26159# a_27422_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1650 vssd1 a_25198_7093# a_25156_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1651 a_5639_10089# _1218_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X1652 a_25313_8207# _1578_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1653 a_2957_27791# _2004_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1654 a_24389_15829# a_24223_15829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1655 vccd1 _1816_.CLK a_2143_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1656 a_17317_4399# a_17047_4765# a_17227_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1657 vccd1 _1880_.CLK a_25143_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1658 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1659 _1527_.A a_19480_17705# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X1662 vccd1 _1862_.Q a_15054_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1663 vssd1 _1905_.Q a_10188_14441# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1665 a_25401_6037# a_25235_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1666 temp1.capload\[0\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1667 a_8998_23439# _0921_.A a_8914_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1669 a_19807_10496# _1129_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1670 a_25953_4399# a_25787_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1671 a_20341_4399# a_20175_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1672 a_20175_12879# _1183_.A2 a_20081_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1673 vssd1 _1342_.B a_4719_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1674 vssd1 _1117_.B a_10417_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1675 a_20690_11445# a_20522_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1676 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1677 a_15557_29789# a_15023_29423# a_15462_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1678 temp1.capload\[3\].cap.Y temp1.capload\[3\].cap_48.LO a_27253_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1679 a_19973_16911# _1914_.Q a_19889_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1680 a_24757_1135# a_24591_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1682 a_27590_9951# a_27422_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1683 vssd1 a_24278_10357# a_24236_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1684 vssd1 a_5047_21237# _1294_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1685 vssd1 a_8177_21781# _1294_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1686 _1502_.A a_20079_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1687 a_12659_11471# a_11877_11477# a_12575_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1689 a_22339_19796# _1689_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1690 vssd1 _1860_.CLK a_11711_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1691 _0909_.X a_3801_28981# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X1692 a_18597_3855# _1935_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1693 vccd1 a_19439_9839# _0952_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1694 a_10452_10089# _1011_.B1 a_10350_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1695 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8307_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1696 vccd1 a_24823_28010# _1902_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1697 a_9323_13103# _1198_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1698 _1007_.X a_19991_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1701 _1436_.X a_10971_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1702 _1313_.A a_2623_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1703 vccd1 _1896_.CLK a_19531_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1704 a_2129_3311# _1798_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1705 vccd1 a_24719_1679# a_24887_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1706 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1707 _0951_.B _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1708 vssd1 _1255_.A1 _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1709 vssd1 _1873_.CLK a_25235_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1710 _1642_.X a_14328_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1711 a_23266_3423# a_23098_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1712 vssd1 _1907_.CLK a_14195_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1713 vssd1 a_19275_3829# a_19233_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1715 vssd1 _0993_.X a_14725_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1716 vssd1 _1234_.A2 a_9123_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X1717 a_15163_2388# _1642_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1718 vssd1 _1459_.A a_15207_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1719 _1032_.C a_18151_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1720 a_12447_17024# _1442_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1721 vccd1 fanout20.X a_22659_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1723 a_24535_10383# a_23837_10389# a_24278_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1724 vssd1 _1764_.B _1764_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1725 vssd1 _1187_.A a_15299_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1726 _1967_.Q a_28015_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1727 vccd1 _1037_.B a_18147_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1728 a_26387_9514# _1677_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1729 vccd1 _1083_.A a_9258_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1730 a_20671_32143# a_19807_32149# a_20414_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1731 vccd1 a_9742_7093# a_9669_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1733 a_23351_25236# _1412_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1734 vccd1 _2006_.Q a_11858_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X1735 a_15097_31061# a_14931_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1736 a_17088_26819# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1738 _1823_.CLK a_22659_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1739 vssd1 _1231_.B1 a_1855_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X1741 a_12384_11177# _1045_.B1 a_12282_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X1743 vssd1 _1775_.C1 _2003_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1744 _1135_.B a_26175_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1745 vssd1 a_9183_12180# _1571_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1746 a_26812_14191# a_26413_14191# a_26686_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1747 a_25708_3311# a_25309_3311# a_25582_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1748 _1914_.Q a_25623_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1749 vccd1 a_11023_16042# _1817_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1751 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1752 a_22195_16911# a_22015_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1753 a_2408_25615# _1762_.Y a_2153_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1754 a_21150_23007# a_20982_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1755 _1616_.A a_9683_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1756 a_26502_25437# a_26063_25071# a_26417_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1757 vssd1 a_12743_11445# a_12701_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1758 a_1857_12015# _1219_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1759 _1471_.A a_14144_26819# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1760 vssd1 _1325_.A2 a_7100_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1761 a_24945_27247# _1835_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1762 a_26295_18218# _1693_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1763 vssd1 a_12631_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1764 a_22779_29789# a_21997_29423# a_22695_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1765 a_18187_28879# a_17489_28885# a_17930_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1766 a_20341_32143# a_19807_32149# a_20246_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1767 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1768 vssd1 a_24639_12180# _1978_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1770 a_5455_20541# _1242_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1771 a_9489_4399# _1753_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1772 a_4338_11177# _1226_.A2 a_4035_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X1773 temp1.capload\[12\].cap.Y temp1.capload\[12\].cap.A a_22101_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1774 a_18371_1501# a_17673_1135# a_18114_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1775 a_9268_24233# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1776 a_24761_2767# _1992_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1777 vssd1 _1121_.A1 a_5588_6825# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1779 a_8484_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1782 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1783 a_15078_2741# a_14910_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1784 a_21192_15055# _1024_.A2 a_20701_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X1786 vccd1 io_in[0] a_2962_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1787 _0909_.A _0903_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1788 vccd1 a_26267_26677# a_26183_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1790 a_8031_13353# _1050_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1791 vssd1 a_25439_2741# a_25397_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1793 vssd1 a_27831_15547# a_27789_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1794 a_18383_3476# _1631_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1795 a_25030_6941# a_24591_6575# a_24945_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1796 a_26007_29789# a_25309_29423# a_25750_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1799 _1108_.A1 a_13571_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1800 a_2455_9295# a_1591_9301# a_2198_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1801 vccd1 a_27647_16635# a_27563_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1802 a_27195_14557# a_26413_14191# a_27111_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1803 vccd1 a_12689_6721# _1069_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1804 a_25106_9269# a_24938_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1805 a_9496_22057# _0921_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1806 a_25823_8207# a_25125_8213# a_25566_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1807 a_2125_6941# a_1591_6575# a_2030_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1808 vssd1 _1896_.CLK a_19439_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1809 vssd1 _1863_.Q a_14144_26819# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1812 a_22195_3855# a_22015_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1813 _1108_.A1 a_13571_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1814 a_20131_27412# _1427_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1815 a_6469_20719# _1286_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1816 a_20337_31433# a_19347_31061# a_20211_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1817 vssd1 _0951_.B a_16097_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1818 a_4345_23145# _1329_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1819 a_1887_13647# _1246_.A2 a_1791_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X1820 _1762_.Y _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1821 vccd1 _1123_.X _1165_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X1822 _1175_.Y _1012_.Y a_7939_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1823 _1183_.A2 a_28015_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1825 a_4804_28111# _1344_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1826 vccd1 fanout33.A a_21279_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1828 vssd1 _1199_.X a_13009_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X1829 a_14852_9839# a_14453_9839# a_14726_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1830 vssd1 a_25639_3855# a_25807_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1831 a_23197_29967# _1843_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1833 _1218_.B a_2715_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1834 vssd1 fanout28.A a_2235_2775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1836 vccd1 _1246_.B2 _1216_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1837 a_4351_17999# _1267_.B1 a_4529_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1839 vssd1 _2005_.Q a_11895_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1840 a_6997_10383# _1086_.Y a_6743_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1841 a_10597_12265# _1015_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1843 a_1766_26159# clkbuf_1_1__f__0380_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1844 _1313_.X a_5455_20541# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X1848 a_10397_14735# _1762_.A a_10594_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1849 a_24554_28853# a_24386_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1850 _1373_.A a_7015_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1851 a_27517_19997# a_26983_19631# a_27422_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1852 a_12981_25615# a_12447_25621# a_12886_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1853 vssd1 _1764_.A _0981_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 a_17397_1679# a_16863_1685# a_17302_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1855 a_24639_23060# _1517_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1856 io_out[2] a_1643_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1857 a_17812_14441# _1033_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X1858 vssd1 a_2715_7931# _1261_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1859 a_18409_3861# a_18243_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1861 _1144_.B a_4003_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1862 vssd1 a_10386_29941# a_10344_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1863 vccd1 _1816_.CLK a_5271_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1864 a_18785_27791# _1842_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1865 a_15078_2741# a_14910_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1866 a_2505_8751# _1222_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1867 _1272_.A2 a_2787_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1868 a_1941_3311# a_1775_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1869 a_19693_2057# a_18703_1685# a_19567_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1870 a_24386_28879# a_24113_28885# a_24301_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1871 vccd1 _1973_.Q a_22238_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X1872 a_27215_31274# _1464_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1873 a_27425_28701# a_26891_28335# a_27330_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1874 _1769_.B1 _1764_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1875 a_22093_5487# _1923_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1876 a_5354_28335# clkbuf_0_temp1.i_precharge_n.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1877 a_4422_1679# a_3983_1685# a_4337_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1878 vccd1 _1074_.C a_16863_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1879 a_12171_3855# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1880 vssd1 a_10931_2986# _1612_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1881 a_16397_6575# a_16127_6941# a_16307_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1882 vssd1 clkbuf_1_1__f__0380_.A a_2686_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1883 a_25030_28701# a_24757_28335# a_24945_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1884 vssd1 _1140_.C a_14533_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1885 _1760_.A_N a_2807_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1886 vccd1 _1133_.C a_20267_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1887 a_23205_26159# _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1888 a_5061_23439# _2009_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1889 vccd1 _1311_.A2 a_1781_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1890 a_20046_31711# a_19878_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1891 vccd1 _1314_.X a_9167_14219# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1892 a_24803_1679# a_24021_1685# a_24719_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1893 vssd1 a_6644_5263# _1226_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 _2003_.D _0913_.A1 a_2601_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1896 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1897 vccd1 _1140_.C a_10791_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1898 vccd1 a_23742_4399# a_23848_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1901 a_10317_19631# _1557_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1902 a_17588_19631# _1828_.Q a_17013_19777# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X1904 a_24665_9301# a_24499_9301# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1905 vccd1 a_3761_9269# _1208_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1906 a_25455_21085# a_24757_20719# a_25198_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1907 _1027_.X a_17139_17024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1908 vssd1 _1092_.B a_9037_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1909 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1910 vssd1 _1322_.A a_5271_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1912 vccd1 a_26099_24527# a_26267_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1913 a_22563_8029# a_22383_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1914 a_27314_8863# a_27146_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1915 a_25198_8863# a_25030_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1916 vssd1 a_7619_2986# _1955_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1917 vssd1 a_13599_1300# _1947_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1918 a_27295_13469# a_26597_13103# a_27038_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1919 _1829_.Q a_21575_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1920 a_10594_14735# a_10814_14709# _0951_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1921 vccd1 a_23799_3855# a_23967_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1922 vssd1 a_26099_24527# a_26267_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1923 vccd1 a_7699_3855# a_7867_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1924 vccd1 a_7625_26677# _1261_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1925 a_16473_16367# _1889_.Q a_16127_16617# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1926 a_24573_2773# a_24407_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1927 a_13487_12559# a_12705_12565# a_13403_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1928 a_1925_23759# _1272_.A2 a_1841_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1929 a_20216_22467# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1930 vccd1 a_8307_5487# _1907_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1931 vccd1 fanout33.A a_18830_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1933 a_11776_28585# a_11527_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1934 vccd1 a_22235_30877# a_22403_30779# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1935 a_23013_21807# _1889_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1936 a_6610_13879# _1012_.Y a_6747_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1937 a_17301_12879# _1890_.Q a_16863_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
R1 vccd1 temp1.capload\[0\].cap_39.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1938 vccd1 a_20414_32117# a_20341_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1939 a_13449_16367# _1021_.A a_13367_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1941 a_25589_23439# _1888_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1942 vssd1 a_25750_3423# a_25708_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1944 a_26225_17289# a_25235_16917# a_26099_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1946 vccd1 _1544_.A_N a_14287_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1948 vccd1 _1824_.Q a_23483_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1949 vccd1 a_25842_6005# a_25769_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1950 vssd1 a_20131_30186# _1869_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1951 a_24209_25615# _1837_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1952 a_6245_14165# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1953 vccd1 a_10643_1679# a_10811_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1955 vccd1 fanout37.A a_15886_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1957 vccd1 _1639_.X a_17415_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1958 vccd1 a_15059_7119# a_15227_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1960 vccd1 a_17359_26525# a_17527_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1961 vccd1 _1639_.X a_12355_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1962 _1801_.Y _1801_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1963 vssd1 _1882_.CLK a_22659_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1965 a_28135_12778# _1713_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1966 vssd1 _1073_.A2 a_17577_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1969 vssd1 a_25807_16635# a_25765_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1970 a_20065_13647# _1877_.Q a_19981_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1971 vccd1 a_18355_28853# a_18271_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1972 vccd1 a_25731_11293# a_25899_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1973 vccd1 a_25623_17723# a_25539_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1974 vssd1 _1305_.B _1306_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1975 a_26785_6575# _1676_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1976 vccd1 a_27847_27613# a_28015_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1977 a_1965_14735# _1277_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1978 vccd1 a_22603_5853# a_22771_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1979 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_10791_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1980 vssd1 _1180_.X a_15667_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1981 _1768_.A a_6835_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1982 _1284_.B1 a_1591_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1983 vccd1 a_21407_2589# a_21575_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1984 a_25156_6575# a_24757_6575# a_25030_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1988 a_1865_22711# a_1673_22453# a_1779_22453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1991 a_5087_29967# _1242_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1993 a_10129_19631# a_9963_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1994 a_19980_16143# _1390_.B a_19405_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X1995 _1645_.A a_14651_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1996 vccd1 fanout24.A a_25143_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1997 a_10727_1679# a_9945_1685# a_10643_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1998 vssd1 _0918_.A _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1999 vssd1 a_17895_17973# a_17853_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2000 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2001 _1809_.B a_6223_3339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2002 a_7458_4765# a_7019_4399# a_7373_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2004 vccd1 _1325_.B1 a_5455_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2005 vssd1 _1024_.X _1034_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2007 a_9574_4765# a_9135_4399# a_9489_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2008 a_10988_27247# a_10589_27247# a_10862_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2010 vssd1 a_12927_15547# a_12885_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2011 vccd1 a_28015_12283# a_27931_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2012 vccd1 a_10627_29691# a_10543_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2013 vccd1 a_2623_2491# a_2539_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2014 vssd1 a_25106_9269# a_25064_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2015 vccd1 _1321_.C a_6223_3339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2016 vccd1 _0939_.A a_11711_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2017 vssd1 a_14894_9951# a_14852_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2018 a_12276_29423# a_11877_29423# a_12150_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2019 vssd1 _1346_.A a_7790_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2020 vccd1 _1054_.C a_15851_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2022 vssd1 _1764_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2023 _0958_.A a_13551_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2024 vccd1 _1855_.Q a_10419_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2025 a_4606_1501# a_4167_1135# a_4521_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2026 vssd1 clkbuf_0_net57.A a_2594_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2027 _1408_.A a_18560_23145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2028 vssd1 a_15163_4564# _1622_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2029 vccd1 a_23450_29941# a_23377_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2030 a_2198_2335# a_2030_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2031 _1723_.X a_22195_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2032 _1189_.C1 a_8859_6144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2033 a_6731_9839# _1122_.A1 _1221_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2034 a_26099_24527# a_25235_24533# a_25842_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2035 vccd1 a_22063_5162# _1960_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2037 a_2030_8207# a_1591_8213# a_1945_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2038 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2039 a_15277_16367# a_14287_16367# a_15151_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2040 vccd1 a_7366_15279# a_7472_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2041 a_18607_11293# a_18427_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2042 vssd1 _1164_.A2 a_7573_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X2043 vccd1 a_15335_2767# a_15503_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2045 a_4209_15529# _1278_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X2046 vccd1 a_27498_28447# a_27425_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2047 a_12478_22057# _1422_.B a_12396_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2048 a_1641_13879# _1246_.B2 a_1791_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X2052 vssd1 _0921_.B _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2053 a_16986_20291# _1405_.B a_16904_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2054 a_22622_1247# a_22454_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2055 a_12575_8207# a_11877_8213# a_12318_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2056 vccd1 fanout20.X a_23855_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2057 vssd1 _1139_.C a_10209_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2058 _1489_.A_N a_12815_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2059 vccd1 _1152_.B a_18642_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2060 a_22545_31599# a_21555_31599# a_22419_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2061 vssd1 a_25842_24501# a_25800_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2062 a_14818_3855# a_14545_3861# a_14733_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2063 a_5911_19881# _1781_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2064 vccd1 _1021_.A a_13919_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2065 a_12189_18150# _0956_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X2066 a_20249_11477# a_20083_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2067 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_18512_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2068 vccd1 a_20046_5599# a_19973_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2069 a_2129_28335# _1775_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2070 vccd1 _0952_.A2 a_20858_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2071 a_4548_2057# a_4149_1685# a_4422_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2072 a_26387_1898# _1650_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2073 vssd1 _1234_.A2 a_4789_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2076 a_27859_29098# _1451_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2077 _1768_.A a_6835_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2078 vccd1 _1532_.A a_12539_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2080 _1553_.A a_7428_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2081 vccd1 _1034_.Y a_8395_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2082 a_4548_25071# a_4149_25071# a_4422_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2083 a_3185_20495# _1328_.S a_3087_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X2084 vssd1 _1101_.X a_15081_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2085 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2086 a_14651_1501# a_14471_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2087 vccd1 _1685_.A_N a_20727_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
R2 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2088 a_9079_2767# a_8215_2773# a_8822_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2089 a_12061_15279# a_11895_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2090 a_23450_29941# a_23282_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2091 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2092 a_23883_3855# a_23101_3861# a_23799_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2093 a_7783_3855# a_7001_3861# a_7699_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2094 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11776_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2095 vccd1 _1887_.CLK a_25235_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2096 a_26099_12559# a_25401_12565# a_25842_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2097 vssd1 a_25198_15391# a_25156_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2098 vssd1 a_25823_22173# a_25991_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2099 vccd1 a_26175_3579# a_26091_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2100 vccd1 _1853_.Q a_6923_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2101 vccd1 _1974_.Q a_27623_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2102 a_20062_28701# a_19623_28335# a_19977_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2104 vccd1 a_5015_1653# a_4931_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2107 a_27713_4399# _1170_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2108 a_10951_22057# a_10423_21807# _0925_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2109 a_14144_17027# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2110 vssd1 _1125_.X a_5496_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2111 a_16945_21629# _1053_.A a_16863_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2112 vssd1 a_24243_16885# a_24201_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2114 _1305_.B a_6559_24640# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2115 vssd1 _1023_.B a_19480_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2116 _1308_.B a_9871_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2119 a_2220_14735# _1247_.B1 a_1965_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2120 vccd1 _1924_.CLK a_24591_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2121 a_25198_7093# a_25030_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2122 a_1769_23145# _0922_.Y _0925_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2123 a_24938_9295# a_24499_9301# a_24853_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2125 a_15538_25589# a_15370_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2127 a_12759_4943# a_11895_4949# a_12502_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2128 a_1829_16341# _1230_.A4 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2129 vssd1 _1819_.Q a_12073_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2130 a_2490_27613# a_2051_27247# a_2405_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2132 _1864_.Q a_20471_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2133 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2134 a_2750_1653# a_2582_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2135 a_10239_28879# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2136 vccd1 _1532_.A a_4627_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2139 vccd1 a_18003_29789# a_18171_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2140 a_16911_1300# _1640_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2141 a_24294_1679# a_23855_1685# a_24209_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2142 a_13288_30345# a_12889_29973# a_13162_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2143 a_9326_23222# _0913_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2144 a_14001_19453# _1021_.A a_13919_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2146 a_2313_25071# _1767_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2147 _1629_.X a_17180_2883# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2148 a_16300_7663# _1041_.A1 a_15725_7809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X2150 vssd1 _1924_.CLK a_24591_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2151 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2152 a_15370_25615# a_15097_25621# a_15285_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2154 vccd1 a_11023_5652# _1356_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2155 a_22120_31599# a_21721_31599# a_21994_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2156 a_25842_4917# a_25674_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2158 vccd1 _1882_.CLK a_22659_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2160 a_2686_10383# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2162 a_10953_19631# a_9963_19631# a_10827_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2163 vssd1 _1846_.Q a_9912_13763# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2164 a_18969_6031# _1321_.C _1807_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2166 vccd1 _1476_.B a_12535_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2167 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_10506_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2169 vssd1 a_15457_6005# _1008_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X2170 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2171 vssd1 _1217_.A3 a_4351_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2172 a_25106_9269# a_24938_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2173 _1371_.A a_8440_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2174 a_25474_11039# a_25306_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2175 vssd1 a_25198_6687# a_25156_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2176 vssd1 a_23691_11195# a_23649_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2177 vccd1 a_2623_9269# a_2539_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2179 vccd1 a_22879_25615# a_23047_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2180 a_15575_19881# _0984_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2181 a_27337_3311# _1674_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2182 vccd1 a_26451_18811# a_26367_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2183 _1469_.A a_14972_26819# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2185 _0956_.C a_7571_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2186 a_21433_14191# _1975_.Q a_21361_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2187 a_14283_6031# a_14103_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2188 a_27337_26159# _1887_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2189 a_9301_5487# a_9135_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2191 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2193 a_21042_16617# _1823_.Q a_20885_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2194 a_9700_4399# a_9301_4399# a_9574_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2195 a_7584_4399# a_7185_4399# a_7458_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2196 a_17041_11177# _1155_.C a_16945_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2197 vssd1 a_22879_25615# a_23047_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2198 a_9761_22357# a_9595_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2199 vssd1 _1325_.B1 a_5455_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2201 a_25723_16733# a_24941_16367# a_25639_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2202 a_8947_9295# a_8767_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2204 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2205 a_2686_15823# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2206 a_14986_4917# a_14818_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2207 a_8447_7828# _1750_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2208 a_22825_27791# a_22291_27797# a_22730_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2209 a_23837_21269# a_23671_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2210 a_15369_4233# a_14379_3861# a_15243_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2211 temp1.capload\[14\].cap.Y temp1.capload\[14\].cap_44.LO a_27897_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2212 a_7019_12265# _1086_.B _1086_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2213 a_25455_15645# a_24591_15279# a_25198_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2214 _1270_.A _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2215 a_4732_1135# a_4333_1135# a_4606_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2216 vccd1 a_24151_8181# a_24067_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2217 vccd1 a_11299_12180# _1847_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2218 vccd1 a_9644_23671# _1336_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2220 a_12691_16367# _0956_.C a_12600_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X2221 a_15741_3311# a_15575_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2222 a_5536_11791# _1794_.Y a_5233_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2223 vssd1 _1841_.CLK a_14931_32149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2224 a_2156_8585# a_1757_8213# a_2030_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2225 a_16198_2589# a_15759_2223# a_16113_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2226 a_22799_7338# _1587_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2228 _1287_.A _1242_.B1 a_6559_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2229 a_18427_11293# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2230 _1893_.Q a_23691_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2231 a_12073_18543# a_11803_18909# a_11983_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2232 a_19480_25321# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2234 vccd1 _1924_.CLK a_25235_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2235 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2236 a_24757_1135# a_24591_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2237 a_10218_29967# a_9945_29973# a_10133_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2238 a_21235_25834# _1513_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2239 vssd1 _1862_.Q a_14972_26819# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2241 a_13130_5737# _1194_.B2 a_12973_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2242 _1092_.B a_10167_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2243 vccd1 _1374_.A_N a_10423_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2244 vssd1 _1816_.CLK a_3983_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2245 _1226_.A2 _1207_.B1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2246 a_25842_4917# a_25674_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2247 _1672_.A a_20999_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2248 vssd1 a_25842_6005# a_25800_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2249 vssd1 _1182_.B a_20308_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2250 a_4351_12879# _1217_.A2 a_4601_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2251 a_2009_21263# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2252 a_16219_17455# _1833_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2253 vccd1 a_25455_13469# a_25623_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2254 vssd1 a_20782_4511# a_20740_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2255 vccd1 _1489_.A_N a_18519_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2256 vssd1 a_22603_5853# a_22771_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2257 _1279_.A1 _1158_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X2259 a_13257_20495# _0913_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 vccd1 _1145_.A1 a_8579_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2262 a_12061_19087# _0956_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X2264 _1397_.A a_16904_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2265 a_17630_7119# _1064_.D1 a_17381_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X2266 vccd1 a_12042_2335# a_11969_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2267 vssd1 _1904_.Q a_8117_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2268 vssd1 a_4059_15431# _1278_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X2269 _1463_.A a_7383_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2270 a_19878_26525# a_19439_26159# a_19793_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2271 vccd1 _1053_.A a_15299_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2272 vccd1 _1269_.A1 a_8454_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X2273 vccd1 a_4404_18517# _1327_.A2_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2274 a_4709_13647# _1217_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2275 a_13599_2388# _1625_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2276 vssd1 a_12189_24825# a_12123_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2277 a_1945_2223# _1793_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2278 _1063_.B a_19735_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2280 vccd1 a_27295_17821# a_27463_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2282 a_19567_17999# a_18869_18005# a_19310_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2283 a_22707_9514# _1601_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2284 a_16707_2589# a_15925_2223# a_16623_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2285 vccd1 a_27755_11293# a_27923_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2287 vssd1 _1217_.B1 a_5048_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2288 a_4842_5737# _1782_.A a_4760_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2289 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2290 a_9644_20871# _1334_.A1 a_9786_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2291 _1189_.B2 a_12743_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2293 vccd1 _1273_.A1 a_5817_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X2295 _1602_.X a_20676_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2296 a_9459_14774# _1122_.A1 a_9000_14967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2297 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2298 _1725_.X a_23299_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2299 a_18751_24148# _1408_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2301 a_2030_1501# a_1591_1135# a_1945_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2302 vccd1 _0918_.A a_10423_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2305 a_1757_8213# a_1591_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2306 vccd1 _1816_.CLK a_2971_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2307 a_16945_11177# _1154_.X a_16863_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2309 vssd1 a_20379_31029# a_20337_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2310 a_23757_9839# a_23487_10205# a_23667_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2311 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A a_7932_25935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2312 vssd1 _1056_.C1 a_14345_24129# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2313 a_25401_12565# a_25235_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2314 _1496_.A a_19480_25321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2315 _1175_.Y _1175_.B2 a_7939_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2317 vccd1 _2006_.Q a_12061_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X2318 _1764_.A a_6927_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2319 vccd1 a_4859_5162# _1365_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2321 vssd1 clkbuf_0_temp1.i_precharge_n.X a_5354_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2322 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2323 a_12171_23983# _0984_.B1 a_12349_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2324 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2325 a_17180_2883# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2326 a_12575_1501# a_11877_1135# a_12318_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2327 vssd1 _0951_.B a_15453_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2328 a_16025_10749# _1010_.A a_15943_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2329 a_9184_23047# _1306_.A2 a_9326_23222# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2331 a_20046_1247# a_19878_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2333 _1690_.A_N a_23671_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2335 vssd1 _1972_.Q a_23113_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2337 vssd1 a_8102_30511# a_8208_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2338 vccd1 a_2807_7093# _1273_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2339 vccd1 a_27590_27359# a_27517_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2340 a_23759_13469# a_23579_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2341 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2342 a_12610_10383# a_12337_10389# a_12525_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2343 vssd1 a_22622_25589# a_22580_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2344 a_20046_1247# a_19878_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2345 a_24420_2057# a_24021_1685# a_24294_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2346 vccd1 _0939_.A a_15299_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2347 a_23374_3855# a_22935_3861# a_23289_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2348 vccd1 _0952_.A1 a_20267_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2349 vccd1 a_27675_29588# _1860_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2350 a_7274_3855# a_6835_3861# a_7189_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2352 a_24554_28853# a_24386_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2353 a_20081_12879# _0958_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X2355 a_17946_1501# a_17673_1135# a_17861_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2356 _1857_.Q a_13755_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2357 a_12604_28585# a_12355_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2358 a_8117_19631# a_7847_19997# a_8027_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2359 a_25014_17973# a_24846_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2361 vssd1 fanout33.A a_21279_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2362 vssd1 _1775_.C1 _2007_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2363 vccd1 _1255_.A1 a_7101_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2364 a_25497_3311# _1990_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2365 a_26513_28879# _1344_.B _1344_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2366 vssd1 a_9135_3311# _1607_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2367 a_17139_6941# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2368 vssd1 _1850_.CLK a_12171_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2369 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2370 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2371 temp1.capload\[1\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2372 a_27337_19631# _1967_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2373 vssd1 _1795_.X a_5536_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2374 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2375 a_9477_17705# _1762_.A a_9674_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2376 vssd1 _1824_.Q a_21192_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2377 a_11848_9839# _1139_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2378 a_23075_11690# _1680_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2379 vccd1 _1876_.CLK a_22015_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2381 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2382 vccd1 a_22898_27765# a_22825_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2383 _1183_.A2 a_28015_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2384 a_16074_5737# _1195_.B2 a_15917_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2385 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2386 a_3069_18793# _1300_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2387 a_13448_14191# _1038_.A1 a_12873_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X2388 vccd1 a_15243_4943# a_15411_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2389 a_22963_31055# a_22181_31061# a_22879_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2390 a_25125_27613# a_24591_27247# a_25030_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2392 vssd1 a_2309_29789# _1760_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X2393 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2395 vccd1 a_25455_7119# a_25623_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2396 vssd1 _1217_.B1 _1277_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X2397 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9963_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2398 vccd1 a_15963_31029# a_15879_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2399 _0997_.X a_15883_13131# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2400 a_14369_8207# _0991_.X a_14453_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2401 vssd1 a_7626_4511# a_7584_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2402 a_25842_26677# a_25674_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2403 vssd1 a_23323_18811# a_23281_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2404 _1628_.A a_15432_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2405 vccd1 _1261_.X a_9135_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2406 vccd1 _1217_.A2 a_5177_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2407 vccd1 _0981_.B a_15299_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2408 _1841_.CLK a_14287_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2409 a_27245_28335# _1886_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2410 _0929_.A a_1591_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2411 vssd1 a_17381_14337# _1034_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X2414 vssd1 _0922_.Y a_3225_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2415 a_11759_29098# _1429_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2416 a_20701_14709# _1024_.A2 a_20858_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2417 vccd1 _1171_.Y a_7295_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9595_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2419 vssd1 _2005_.Q a_6927_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2421 a_2686_26703# clkbuf_0_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2422 vssd1 a_4774_1247# a_4732_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2423 vccd1 _2023_.CLK a_1591_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2424 a_24021_1685# a_23855_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2425 vssd1 a_15630_29535# a_15588_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2427 vssd1 _1140_.C a_9841_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2428 vccd1 _1119_.A1 a_16064_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X2429 _1246_.B2 _1221_.A a_1677_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2430 a_24389_1679# a_23855_1685# a_24294_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2432 a_25674_26703# a_25401_26709# a_25589_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2433 a_13408_24233# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2434 a_23239_24349# a_22457_23983# a_23155_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2435 a_25842_22325# a_25674_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2436 a_16324_2223# a_15925_2223# a_16198_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2437 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2438 _0921_.B a_3983_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2439 a_23113_20719# a_22843_21085# a_23023_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2440 _1175_.B2 _1198_.A2 a_10597_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2441 vssd1 _1855_.CLK a_14287_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2442 vccd1 a_20303_26525# a_20471_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2443 vccd1 a_27463_13371# a_27379_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2444 vccd1 _1074_.C a_15207_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2445 a_16208_11791# _1119_.A1 a_15633_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X2446 a_26777_4399# a_25787_4399# a_26651_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2447 a_23266_4917# a_23098_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2450 vssd1 a_26267_16885# a_26225_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2451 vssd1 _1841_.CLK a_14931_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2452 a_10589_27247# a_10423_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2454 a_14641_9839# _1571_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2455 vccd1 _1544_.A_N a_10331_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2456 vccd1 a_13755_29941# a_13671_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2457 vssd1 fanout28.A a_15115_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2459 _1280_.Y _1234_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X2460 a_24604_19465# a_24205_19093# a_24478_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2461 a_9674_17705# a_9894_17429# _0981_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2462 vccd1 _0998_.B2 a_19619_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2463 vccd1 a_14986_3829# a_14913_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2465 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_11527_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2466 a_27590_26271# a_27422_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2467 a_24573_18005# a_24407_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2469 a_5909_16143# _1313_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 _1191_.B1 a_19103_13985# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2471 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2472 _1507_.A a_19664_23555# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2473 vccd1 _1723_.A_N a_23119_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2475 a_16573_4399# a_16396_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2478 vssd1 _1448_.A a_11711_15831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2479 vssd1 _1038_.X _1050_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2480 vssd1 _1159_.X a_5893_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2481 _2003_.Q a_3083_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2482 a_22821_29423# a_21831_29423# a_22695_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2484 vssd1 _1313_.A a_2327_20183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2485 vssd1 _1053_.A a_15299_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2486 vccd1 _1344_.Y a_9135_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2487 vssd1 _2007_.Q a_8307_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2488 a_6084_15529# _1289_.B1 a_5829_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2490 vssd1 _0973_.B a_21917_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2491 a_19701_31055# _1473_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2492 a_22155_23658# _1691_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2493 vccd1 a_23523_3677# a_23691_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2494 vssd1 _1839_.Q a_12396_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2495 vccd1 a_9247_2741# a_9163_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2496 a_10188_14441# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2497 vccd1 _1153_.A a_19807_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2498 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11796_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2499 a_22178_6941# a_21739_6575# a_22093_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2500 a_18682_2767# a_18409_2773# a_18597_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2503 vccd1 _1489_.A_N a_19439_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2505 vccd1 a_19735_17973# a_19651_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2507 a_19889_16911# _0953_.C1 a_19807_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2508 a_14139_1679# a_13275_1685# a_13882_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2509 a_12349_12015# a_12079_12381# a_12259_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2510 a_20775_30186# _1485_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2511 a_22622_24501# a_22454_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2512 _1108_.C1 a_11711_14848# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2513 a_2156_1135# a_1757_1135# a_2030_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2514 vccd1 a_16267_27412# _1542_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2515 a_7755_22351# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2517 a_27422_12381# a_26983_12015# a_27337_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2518 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2519 _1542_.A a_13408_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2520 a_20267_9295# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2521 _0952_.A1 a_19439_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2522 vssd1 a_10202_27765# a_10160_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2523 vssd1 fanout24.A a_24499_9301# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2524 vccd1 _1108_.A1 a_11834_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2525 a_1929_10749# _1177_.Y a_1857_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2526 vssd1 _1198_.A2 a_9323_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X2527 a_2129_7119# _1791_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2528 vccd1 fanout21.X a_25143_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2529 _1329_.X a_2103_31573# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2530 vccd1 _0909_.A _1308_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2532 vccd1 a_10202_22325# a_10129_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2533 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_6559_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2534 a_16267_27412# _1542_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2535 vssd1 _0922_.Y a_2029_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2536 a_22553_20175# _1822_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2537 _1442_.A a_15319_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2538 a_22879_1501# a_22015_1135# a_22622_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2539 a_19793_31599# _1540_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2540 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2541 a_1673_20969# _1270_.A a_1591_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2542 vssd1 fanout24.A a_23671_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2543 a_12321_22325# _1142_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X2544 vssd1 a_3983_19631# _0918_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2545 vccd1 _0961_.A a_12447_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2546 vccd1 a_12927_4917# a_12843_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2547 _1092_.B a_10167_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2549 temp1.inv2_2.Y temp1.inv2_2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2550 a_6600_7913# _1809_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2551 a_27590_5599# a_27422_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2552 vccd1 _0958_.A a_11895_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2553 vssd1 _1231_.B1 _1250_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2555 a_27295_6941# a_26597_6575# a_27038_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2556 vssd1 a_19439_9839# _0952_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2557 a_21051_22570# _1404_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2558 a_10459_2589# a_9595_2223# a_10202_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2559 a_25455_9117# a_24591_8751# a_25198_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2560 a_20815_10205# a_20635_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2562 vssd1 _1823_.CLK a_26983_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2564 a_27571_9117# a_26707_8751# a_27314_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2565 a_7550_2589# a_7111_2223# a_7465_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2566 vssd1 _1448_.A a_7571_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2567 _1242_.A1 a_2623_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2568 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12604_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2569 a_3324_18793# _1300_.B1 a_3069_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2570 _1640_.X a_17595_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2571 vccd1 _1489_.A_N a_22015_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2573 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8484_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2574 vccd1 a_2807_6005# _1255_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2575 _1440_.B a_17159_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2576 a_8546_1653# a_8378_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2577 _1168_.X a_6867_8545# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2578 a_16863_10496# _1089_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2579 vccd1 a_17527_31867# a_17443_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2580 a_23500_4233# a_23101_3861# a_23374_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2581 a_25129_3855# _1745_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2582 a_21813_26525# a_21279_26159# a_21718_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2584 a_7400_4233# a_7001_3861# a_7274_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2585 a_17773_21629# _0961_.A a_17691_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2586 _1558_.X a_10188_14441# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2589 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R3 vssd1 temp1.capload\[9\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2590 vssd1 a_19487_2388# _1993_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2591 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_12631_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2595 a_12065_8207# _1561_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2596 a_19057_14735# _1399_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2597 vccd1 a_25198_27359# a_25125_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2598 vssd1 _0984_.A2 a_12609_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2600 a_15391_8320# _1109_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2602 a_15531_15444# _1398_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2604 a_6645_10089# _1123_.X _1221_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2605 vssd1 _1869_.Q a_16904_25731# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2606 a_24278_21237# a_24110_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2607 a_16991_9117# a_16293_8751# a_16734_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2608 a_15097_25621# a_14931_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2611 a_23903_1300# _1736_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2612 a_25014_2741# a_24846_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2613 vssd1 a_7515_1501# a_7683_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2614 a_5169_10749# _1304_.B a_5087_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2617 a_19878_26525# a_19605_26159# a_19793_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2618 _1119_.C1 a_11803_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2619 vccd1 _0923_.Y a_7050_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2620 a_19617_20719# _1883_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2621 a_17139_18793# _1024_.A2 a_17221_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2622 vccd1 _1231_.B1 a_4173_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2623 vccd1 _1034_.Y a_8031_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2624 vccd1 _1329_.S a_6914_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X2625 a_1937_22711# _1242_.B1 a_1865_22711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X2626 vccd1 _0994_.B2 a_15387_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2628 a_23903_24746# _1507_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2629 a_22457_23983# a_22291_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2630 _1433_.A a_10188_18115# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2631 a_26226_8029# a_25953_7663# a_26141_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2632 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4804_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2633 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE a_8951_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2634 _1242_.A2 a_7111_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2635 vccd1 a_2915_24349# a_3083_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2636 a_23818_23413# a_23650_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2637 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2638 a_15614_6031# _0963_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2639 vssd1 a_22751_22895# _1882_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2642 a_17762_28879# a_17489_28885# a_17677_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2643 vccd1 _1424_.A_N a_18243_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2644 vssd1 a_2823_25437# a_2991_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2645 _1254_.A2 a_2143_17705# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2646 a_5629_7913# _1172_.X a_5547_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2647 a_14533_9661# _1030_.B a_14461_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2649 a_14913_3855# a_14379_3861# a_14818_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2650 vssd1 _1140_.C a_9013_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2651 a_5265_21263# _1261_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2653 a_3210_24501# a_3042_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2654 vssd1 a_23155_27791# a_23323_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2655 a_12529_17277# _0961_.A a_12447_17024# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2656 a_2290_13215# a_2122_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2657 a_8803_1679# a_8105_1685# a_8546_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2658 vccd1 a_25842_20149# a_25769_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2659 a_21533_7663# a_20543_7663# a_21407_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2660 a_13012_25993# a_12613_25621# a_12886_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2661 vssd1 _1816_.CLK a_8215_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2662 vssd1 a_16366_2335# a_16324_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2663 a_11707_4765# a_11527_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2664 vccd1 _1317_.X a_5487_5281# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2665 a_13304_14441# _0984_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X2666 vccd1 _1830_.Q a_15387_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2667 a_2696_11177# _1207_.B1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2668 a_2029_20719# _1768_.A a_1591_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2669 vssd1 a_26203_10602# _1728_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2671 a_7001_3861# a_6835_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2672 vccd1 _1141_.C a_17139_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2673 a_23469_3855# a_22935_3861# a_23374_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2674 vccd1 _2023_.CLK a_1591_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2675 a_7369_3855# a_6835_3861# a_7274_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2676 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12532_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2677 _1706_.X a_22931_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2678 vccd1 _1071_.B1 a_13551_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2679 a_19233_3145# a_18243_2773# a_19107_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2680 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2682 vssd1 _1985_.Q a_23389_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2683 a_23849_13103# a_23579_13469# a_23759_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2684 a_21031_28879# a_20249_28885# a_20947_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2685 a_26965_21807# a_26799_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2686 _0981_.B _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2687 a_11885_6575# _1010_.A a_11803_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2689 _1531_.A a_19619_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2690 a_23266_4917# a_23098_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2691 a_27314_8863# a_27146_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2692 vssd1 _1282_.A2 a_6369_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X2693 vccd1 a_12575_13647# a_12743_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2694 a_25765_4233# a_24775_3861# a_25639_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2695 a_1644_18517# _1231_.B1 a_2036_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2697 a_16945_12559# _0999_.C1 a_16863_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2699 a_27498_28447# a_27330_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2700 vssd1 clkbuf_1_1__f__0380_.A a_2686_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2701 _1617_.X a_11707_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2703 vssd1 _1068_.C1 a_12689_6721# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2705 vccd1 a_3983_19631# _0918_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2706 vssd1 a_12575_13647# a_12743_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2707 a_20407_24746# _1414_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2709 _1223_.A2 a_12927_13103# a_13165_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X2710 a_15477_2045# a_15207_1679# a_15387_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2711 _1065_.X a_15299_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2714 vssd1 _1924_.CLK a_24591_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2715 a_6375_6941# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2716 a_5183_21583# _1282_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X2717 a_25589_6031# _1591_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2718 _1252_.A a_5361_11191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2719 _0989_.A2 a_3175_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2720 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2721 vssd1 a_24278_21237# a_24236_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2722 a_22304_6575# a_21905_6575# a_22178_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2723 vccd1 _1823_.CLK a_22199_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2726 a_24639_4564# _1670_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2727 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_5639_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2728 vccd1 a_2639_28701# a_2807_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2729 vssd1 _1775_.A2 _0923_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2730 vssd1 a_6283_4399# _1999_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2731 _1474_.A_N a_8215_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X2733 vccd1 a_24703_10357# a_24619_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2734 vssd1 _1040_.B a_21273_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2735 vssd1 a_2198_1247# a_2156_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2736 vccd1 a_19107_3855# a_19275_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2737 vssd1 a_28015_26427# a_27973_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2738 a_25309_9839# a_25143_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2739 a_20429_29423# a_19439_29423# a_20303_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2740 _1190_.B1 a_21127_12897# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2741 a_10589_3311# a_10423_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2742 vssd1 fanout33.A a_18830_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2743 a_4250_8207# _1205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X2744 vccd1 a_26651_8029# a_26819_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2746 vssd1 _1102_.B a_19709_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2748 vccd1 _1074_.C a_11343_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2749 a_9591_11293# a_9411_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2750 vccd1 _1170_.A2 a_1814_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2751 a_13551_11471# _1143_.X a_13805_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2752 a_24535_21263# a_23837_21269# a_24278_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2753 a_9772_27247# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2754 vssd1 a_21407_23261# a_21575_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2755 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2756 a_15840_21583# _1844_.Q a_15265_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X2757 vssd1 a_14103_10383# _1110_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2758 vssd1 a_2971_16367# _0921_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2759 a_11313_14191# _1846_.Q a_11241_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2760 a_5455_27791# _1242_.B1 _0913_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X2761 _1450_.A a_6923_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2762 _2006_.Q a_3635_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2763 vccd1 a_23615_22351# a_23783_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2764 vccd1 _1293_.A1 a_8395_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2765 a_2129_6031# _2019_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2766 a_25539_6941# a_24757_6575# a_25455_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2767 vccd1 a_21143_8916# _1605_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2769 a_1828_19061# _1270_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X2770 a_3299_22325# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X2771 a_26413_14191# a_26247_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2773 vccd1 a_21886_26271# a_21813_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2774 _0958_.B a_14563_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2775 _1061_.X a_18795_7232# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2776 vccd1 _1038_.A1 a_9591_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2777 a_18751_24148# _1408_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2778 a_7676_2223# a_7277_2223# a_7550_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2779 io_out[4] a_4220_21959# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2781 a_25363_9295# a_24499_9301# a_25106_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2782 a_9945_29973# a_9779_29973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2783 _1894_.Q a_25623_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2785 vccd1 a_11023_26922# _1858_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2786 vssd1 a_23615_22351# a_23783_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2787 a_25581_1135# a_24591_1135# a_25455_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2789 a_12752_22351# _1142_.B1 a_12650_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2790 a_13530_31055# a_13091_31061# a_13445_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2791 vccd1 a_10627_27765# a_10543_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2792 a_22645_27791# _1876_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2795 a_23389_14191# a_23119_14557# a_23299_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2796 a_19991_13103# _1191_.B1 a_20169_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2797 a_19605_1135# a_19439_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2798 a_24386_28879# a_23947_28885# a_24301_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2799 a_6923_16617# _1788_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2800 a_2214_4943# a_1941_4949# a_2129_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2802 a_17359_26525# a_16661_26159# a_17102_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2803 a_10386_8181# a_10218_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2804 vccd1 a_17139_9839# _1293_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2805 _1652_.X a_3748_3971# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2806 a_9945_6037# a_9779_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2807 vssd1 _1050_.C _1050_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2808 _1416_.A a_18423_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2809 vssd1 a_9742_5599# a_9700_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2810 vssd1 _1139_.C a_9749_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2811 vccd1 a_12815_9295# _1459_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2812 vccd1 _1869_.Q a_16986_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2814 vssd1 _1841_.CLK a_17323_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2815 a_11371_27613# a_10589_27247# a_11287_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2816 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2817 a_14335_2388# _1619_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2818 a_5687_4564# _1756_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2820 _1142_.D1 a_11895_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2821 vccd1 _1133_.C a_19471_16395# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2822 a_3578_2741# a_3410_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2824 _1222_.B1 a_2644_11587# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X2825 vccd1 a_9889_25913# a_9919_25654# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2826 a_12575_13647# a_11711_13653# a_12318_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2827 a_26183_6031# a_25401_6037# a_26099_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2828 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2829 _1914_.Q a_25623_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2831 vccd1 _1226_.A1 a_3065_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2832 vssd1 _1189_.C1 a_10515_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2833 _1401_.A a_15387_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X2834 a_25769_13647# a_25235_13653# a_25674_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2835 vccd1 _0961_.A a_11067_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2836 a_19619_19997# a_19439_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2837 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2838 a_22806_20149# a_22638_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2840 vccd1 a_7803_20884# _1852_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
R4 vssd1 temp1.capload\[2\].cap_47.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2841 vccd1 _1030_.B a_12351_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2843 a_3095_9867# _1177_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2845 a_1674_30511# clkbuf_0_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2847 a_15335_2767# a_14637_2773# a_15078_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2848 vssd1 a_8447_10004# _1563_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2849 vssd1 fanout37.A a_23395_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2850 a_12245_13647# a_11711_13653# a_12150_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2851 vssd1 a_2623_8181# _1242_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2852 _1897_.Q a_20471_31867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2854 _1140_.C a_7442_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X2856 vccd1 _1639_.X a_7019_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2857 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2858 vccd1 _1860_.CLK a_11711_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2859 vccd1 _1195_.A2 a_16074_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2860 _1033_.A2 a_18551_11809# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2861 vccd1 _1924_.CLK a_21739_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2862 a_3467_27791# a_2769_27797# a_3210_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2863 vssd1 a_10423_21807# _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2864 a_16661_31599# a_16495_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2865 _1074_.C _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2866 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2867 _1112_.D1 a_19439_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X2868 a_23098_3677# a_22825_3311# a_23013_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2869 a_7373_4399# _1816_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2870 a_4127_22869# _1337_.S a_4558_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X2871 _1046_.B a_28015_12283# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2872 vccd1 a_23523_4943# a_23691_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2873 _1826_.Q a_25071_19061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2875 vssd1 a_10423_23983# _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2877 a_18114_32117# a_17946_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2878 _1081_.B1 a_21463_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2879 a_19310_14709# a_19142_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2880 vccd1 _1242_.B1 a_5639_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2881 vccd1 a_6559_9295# _0930_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2883 a_14776_15529# _1095_.B1 a_14674_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X2884 a_9949_22351# _1817_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2885 vccd1 a_21150_2335# a_21077_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2886 _1681_.X a_21643_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2887 a_18497_31433# a_17507_31061# a_18371_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2890 vccd1 _1873_.CLK a_26891_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2891 a_7619_26324# _1373_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2892 a_23615_22351# a_22751_22357# a_23358_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2893 vccd1 a_2623_2491# _1286_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2894 vssd1 a_11023_16042# _1817_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2895 vccd1 fanout33.A a_19439_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2896 a_18072_1135# a_17673_1135# a_17946_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2898 a_26965_21807# a_26799_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2899 vccd1 _1459_.A a_22015_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X2900 a_3578_2741# a_3410_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2901 a_21031_27791# a_20249_27797# a_20947_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2902 a_11067_15529# _0987_.B _0987_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2903 vssd1 _0998_.A2 a_17685_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2904 a_18785_28111# _1872_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2907 a_27011_25437# a_26229_25071# a_26927_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2908 _0921_.A a_2971_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2910 vssd1 _1013_.X a_9779_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2911 a_7728_31055# a_7479_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2912 a_8113_25117# _0911_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2913 a_16934_31965# a_16495_31599# a_16849_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2916 vssd1 a_22346_6687# a_22304_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2917 vccd1 _0963_.B a_16035_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2918 vssd1 _2006_.Q a_6835_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2919 a_25589_16911# _1527_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2920 a_12500_15797# _1820_.Q a_12720_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2921 a_23285_22351# a_22751_22357# a_23190_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2922 vccd1 a_18850_2741# a_18777_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2923 a_21051_22570# _1404_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2924 a_5996_19631# _0909_.B a_5693_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2925 _1325_.B1 a_5269_13367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2926 vccd1 a_14307_1653# a_14223_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2927 a_27839_11293# a_27057_10927# a_27755_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2928 vccd1 a_7442_17429# _1140_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.135 ps=1.27 w=1 l=0.15
X2929 vccd1 a_14323_24527# a_14491_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2930 _1773_.B a_4035_23957# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2931 _1020_.A2 a_19471_16395# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2932 vssd1 a_22622_26677# a_22580_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2933 vccd1 _0985_.X a_9309_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2934 _1592_.X a_18560_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2935 _1443_.A a_9360_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2936 a_17811_17999# a_17029_18005# a_17727_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2938 a_3979_9295# _1175_.Y a_3761_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2939 vssd1 _0987_.Y a_12528_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X2940 vssd1 a_14323_24527# a_14491_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2941 _1780_.B1 a_4259_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2942 a_21039_4765# a_20175_4399# a_20782_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2943 a_21138_16367# _1985_.Q a_21048_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X2944 _1008_.X a_14839_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X2945 a_9411_11293# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2946 _1896_.Q a_20839_32117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2947 vssd1 _1768_.A a_9135_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2948 a_15163_2388# _1642_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2949 a_6099_27247# _2009_.CLK _0909_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2951 a_15453_6575# _1065_.B a_15381_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2952 vssd1 a_12743_29691# a_12701_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2953 _1896_.Q a_20839_32117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2954 a_12153_23145# _1853_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2955 _0925_.A2 a_10423_21807# a_10951_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2956 a_22879_26703# a_22181_26709# a_22622_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2957 a_12042_25183# a_11874_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2958 vssd1 _0958_.B a_17845_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X2959 vccd1 _1438_.B a_12259_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2960 a_13091_19200# _1863_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2961 vccd1 a_10627_2491# a_10543_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2962 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2963 vccd1 a_25623_9019# a_25539_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2964 a_17673_32149# a_17507_32149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2965 vssd1 a_7718_2335# a_7676_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2966 a_22454_26703# a_22015_26709# a_22369_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2967 a_10402_19997# a_9963_19631# a_10317_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2968 a_5541_3311# _1321_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2969 a_24846_2767# a_24573_2773# a_24761_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2970 a_23351_25236# _1412_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2971 vccd1 a_22659_17455# _1823_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2972 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2973 vccd1 a_26007_29789# a_26175_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2974 vccd1 a_24462_25589# a_24389_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2975 a_15255_23060# _1545_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2976 a_24761_17999# _1976_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2977 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2978 a_7967_4765# a_7185_4399# a_7883_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2980 a_10202_2335# a_10034_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2981 vccd1 a_24979_28853# a_24895_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2982 a_12150_8207# a_11711_8213# a_12065_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2983 _1841_.Q a_18539_32117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2984 vccd1 a_2807_28603# a_2723_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2985 a_2686_10383# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X2986 vccd1 _0939_.A a_14287_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2987 vssd1 _1835_.Q a_20261_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2990 a_26387_9514# _1677_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2991 vccd1 a_25623_28603# a_25539_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2992 a_20499_23658# _1410_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2994 a_7199_1679# a_7019_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2996 _1841_.Q a_18539_32117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2997 a_3111_5652# io_in[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2998 vccd1 _1337_.S a_2339_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X2999 vccd1 _1882_.CLK a_26063_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3000 temp1.capload\[5\].cap.Y temp1.capload\[5\].cap.A a_26057_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3002 a_6929_22057# _0921_.Y a_6847_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3003 a_22081_14709# _1293_.A1 a_22334_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3004 a_21279_3677# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3005 vccd1 fanout24.A a_24039_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3006 vccd1 _1832_.Q a_18918_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X3007 vssd1 a_10386_8181# a_10344_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3008 vccd1 _1353_.A a_26513_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3009 a_23377_23445# a_23211_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3010 vccd1 _0981_.B a_13091_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3011 vssd1 _1826_.Q a_18560_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3012 vccd1 _1723_.A_N a_23119_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3013 a_25198_31711# a_25030_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3016 vssd1 _1976_.Q a_23021_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3017 vccd1 a_12318_13621# a_12245_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3019 a_8654_29967# a_8477_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3020 _1095_.B1 a_11711_12672# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3022 vccd1 a_26394_7775# a_26321_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3024 _1901_.Q a_13479_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3025 a_10349_25045# _1274_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3026 a_4262_24305# a_4213_24135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X3027 vssd1 a_26819_4667# a_26777_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3028 a_23523_4943# a_22659_4949# a_23266_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3029 a_23649_8751# a_22659_8751# a_23523_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3030 a_27038_24095# a_26870_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3032 a_10589_27247# a_10423_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3034 a_27149_5487# a_26983_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3036 a_25907_22173# a_25125_21807# a_25823_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3039 a_18601_21629# _1132_.A a_18519_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3041 a_27847_5853# a_26983_5487# a_27590_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3042 vssd1 _1403_.B a_19709_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3043 a_20131_27412# _1427_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3044 _1830_.CLK a_15115_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3045 vccd1 _1982_.CLK a_22015_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3046 _1598_.X a_19112_9411# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3047 vssd1 _1353_.Y a_7479_28887# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3048 _1901_.Q a_13479_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3049 a_23005_2057# a_22015_1685# a_22879_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3050 a_20223_8426# _1582_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3051 a_23005_24905# a_22015_24533# a_22879_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3052 a_25198_1247# a_25030_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3053 a_20905_9839# a_20635_10205# a_20815_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3054 vccd1 _1860_.CLK a_9595_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3056 a_21545_15279# _0939_.A a_21463_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3058 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3059 vccd1 _1744_.A_N a_20083_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3060 a_27897_27023# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3061 vssd1 _1849_.CLK a_13643_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3062 a_2214_7119# a_1775_7125# a_2129_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3064 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3065 a_9949_29423# _1903_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3066 vssd1 _0921_.B a_10423_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3067 a_17489_28885# a_17323_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3068 a_7002_4943# _1202_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3070 vssd1 _1999_.CLK a_13275_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3071 a_15381_20291# _1186_.X a_15299_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X3072 vssd1 _1139_.C a_11865_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3073 _1440_.B a_17159_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3074 vssd1 _1190_.B1 a_22648_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X3075 a_22178_5853# a_21905_5487# a_22093_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3076 vccd1 a_20471_31867# a_20387_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3078 a_25309_16733# a_24775_16367# a_25214_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3079 _1170_.A3 a_4447_6581# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X3081 vssd1 _0965_.A2 a_18140_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X3082 a_2861_17999# _1281_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3083 vssd1 _1970_.Q a_22193_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3084 a_26965_15279# a_26799_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3086 vssd1 a_24719_1679# a_24887_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3087 vccd1 fanout24.A a_26707_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3088 vssd1 _1436_.B a_12268_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X3089 vssd1 a_21575_7931# a_21533_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3092 vssd1 a_23047_1653# a_23005_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3094 a_27153_21807# _1878_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3095 a_16113_2223# _1947_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3096 vssd1 a_18114_1247# a_18072_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3097 vccd1 a_2382_28447# a_2309_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3098 vccd1 _1801_.B a_4896_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X3099 a_20138_30623# a_19970_30877# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3100 vccd1 a_11760_24759# _1352_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3102 vccd1 a_23358_22325# a_23285_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3103 a_19142_1679# a_18869_1685# a_19057_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3104 _1177_.Y _1175_.Y a_3873_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3105 a_15285_25615# _1900_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3106 a_1683_27791# _1775_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3108 _1132_.X a_14839_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3109 vccd1 _0958_.A a_7009_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3110 a_10227_11471# _1121_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3111 a_19928_18793# _1184_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X3112 vssd1 _1316_.A a_6870_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3113 a_5031_1501# a_4167_1135# a_4774_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3114 a_1765_9001# _1232_.Y _1300_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3115 vccd1 _1474_.A_N a_14563_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3116 vssd1 _1259_.X a_2706_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X3117 vccd1 a_26267_12533# a_26183_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3118 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3119 a_4149_25071# a_3983_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3120 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_7925_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3122 a_9000_14967# _1122_.A1 a_9142_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3123 vssd1 _1924_.CLK a_24959_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3124 a_14405_7691# _0935_.X a_14319_7691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3125 vccd1 _1058_.B a_6555_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3126 a_8454_15797# _1764_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3127 a_18455_32143# a_17673_32149# a_18371_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3128 _1973_.Q a_25623_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3129 a_1791_13967# _1246_.B1 a_1641_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X3130 a_26870_13469# a_26597_13103# a_26785_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3131 vccd1 _1147_.X a_17113_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3132 a_20648_29257# a_20249_28885# a_20522_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3133 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3134 _1061_.B a_27739_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3135 vccd1 _1982_.CLK a_23303_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3136 _1177_.C _1173_.X a_7742_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X3137 a_27295_17821# a_26597_17455# a_27038_17567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3138 vssd1 _1075_.C a_18085_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
R5 vssd1 temp1.capload\[3\].cap_48.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3140 a_26927_25437# a_26229_25071# a_26670_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3141 a_12429_15645# a_11895_15279# a_12334_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3142 a_6559_4943# _1208_.A1 a_6644_5263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3143 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3144 a_21633_26159# _1838_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3146 a_15925_2223# a_15759_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3147 vccd1 _1985_.CLK a_26983_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3149 a_26099_23439# a_25401_23445# a_25842_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3150 _1977_.Q a_27463_13371# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3151 vccd1 a_8143_2491# a_8059_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3152 _1614_.A a_10464_1385# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3153 vccd1 _1850_.CLK a_3983_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3154 a_27215_31274# _1464_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3155 vssd1 _1032_.C a_19189_13985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3156 vccd1 _1723_.A_N a_22015_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3157 a_19709_19631# a_19439_19997# a_19619_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3158 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3160 vssd1 _0963_.B a_14441_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3162 vssd1 a_27859_30186# _1456_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3163 a_8102_30511# a_7925_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3165 a_14144_27907# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3166 a_2750_1653# a_2582_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3167 vccd1 a_20303_1501# a_20471_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3168 vssd1 a_13057_8897# _1069_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X3170 a_10154_20495# _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X3172 a_27697_2223# a_26707_2223# a_27571_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3173 a_16904_3971# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3174 _1802_.X a_4116_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3176 vccd1 _1849_.CLK a_18703_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3179 _1835_.Q a_25623_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3180 vssd1 _1985_.CLK a_25235_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3181 _1858_.Q a_16055_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3182 a_13395_25615# a_12613_25621# a_13311_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3183 vssd1 a_27406_21919# a_27364_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3184 vssd1 _1074_.C a_17809_20513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3185 a_7939_13967# _1012_.Y _1175_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3187 a_18642_18793# _1405_.B a_18560_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3188 a_3593_24905# a_2603_24533# a_3467_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3189 vssd1 _1108_.X a_14287_13353# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3190 a_8498_20214# _1232_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3191 vssd1 _1269_.A1 _0951_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3192 vccd1 a_25531_9269# a_25447_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3193 vssd1 _1086_.Y a_4669_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3195 vssd1 a_9460_25847# _1337_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3196 a_20349_15279# _1127_.A a_20267_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3197 a_12893_12559# _1911_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3198 a_21695_17620# _1391_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3199 _1042_.B a_15411_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3200 a_13766_14735# _1107_.X a_13517_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3201 vssd1 a_18539_32117# a_18497_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3202 a_19487_4564# _1636_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3203 a_10423_9117# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3204 vssd1 _1186_.C1 a_11987_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3205 a_22983_19796# _1385_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3206 vssd1 a_2455_9295# a_2623_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3207 _0984_.A2 a_12295_20747# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3208 _1711_.X a_23299_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3209 a_10048_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3210 vccd1 a_20315_25236# _1838_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3211 _1775_.C1 a_7387_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3212 a_14920_15279# _1821_.Q a_14345_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X3213 vssd1 _1104_.C a_15115_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3215 a_22193_16367# a_21923_16733# a_22103_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3217 a_17673_31061# a_17507_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3218 a_6236_25071# _1306_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X3219 vssd1 a_22063_5162# _1960_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3220 vccd1 a_2382_4917# a_2309_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3221 a_12276_8585# a_11877_8213# a_12150_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3222 a_5165_2828# _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3223 a_26133_29423# a_25143_29423# a_26007_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3224 a_26225_27081# a_25235_26709# a_26099_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3225 vccd1 _1985_.CLK a_23947_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3226 a_26321_8029# a_25787_7663# a_26226_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3227 _0964_.A a_13183_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3228 vccd1 a_22707_18218# _1878_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3229 a_10213_15939# _2005_.Q a_10141_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3230 a_15538_32117# a_15370_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3231 a_15243_4943# a_14545_4949# a_14986_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3232 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3234 a_4800_7663# _1126_.Y a_4497_7637# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3235 vssd1 a_4587_24501# _1767_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3236 vssd1 a_21143_8916# _1605_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3238 _1646_.X a_13455_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3239 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3241 a_17845_21629# _1886_.Q a_17773_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3243 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_15750_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3244 vssd1 _0909_.X a_25695_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3245 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3247 a_18305_10749# _1080_.B a_18233_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3251 a_20004_29423# a_19605_29423# a_19878_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3252 a_3007_1679# a_2309_1685# a_2750_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3253 _2007_.D _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3255 a_20267_17455# _1969_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3256 vccd1 _1270_.A _1270_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3257 vssd1 a_23691_22075# a_23649_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3258 _1536_.A a_18699_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3259 a_25198_27359# a_25030_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3260 vssd1 a_12873_14337# _1038_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X3261 a_22181_1685# a_22015_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3262 a_28135_12778# _1713_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3263 a_21073_28169# a_20083_27797# a_20947_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3264 vssd1 _2023_.CLK a_1591_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3268 vssd1 a_11759_7338# _1657_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3269 a_27245_10927# _1586_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3270 a_4324_29673# a_4075_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3273 a_16934_31965# a_16661_31599# a_16849_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3274 a_19439_20719# _1184_.B1 a_19617_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3275 a_22879_31055# a_22015_31061# a_22622_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3276 a_19326_29967# a_19149_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3277 a_14901_19453# _1864_.Q a_14829_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3278 a_11413_3311# a_10423_3311# a_11287_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3279 vssd1 _1008_.X a_10021_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3280 a_2686_26703# clkbuf_0_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3281 a_16245_20747# _1053_.A a_16159_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3282 a_9489_5487# _2001_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3283 a_2198_6687# a_2030_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3284 vccd1 _1337_.S a_5203_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X3286 a_18107_21972# _1397_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3287 a_7885_17455# _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.212875 ps=1.305 w=0.65 l=0.15
X3288 vccd1 a_17573_4917# _1155_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3289 vccd1 a_20867_8426# _1599_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3292 a_24941_16367# a_24775_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3293 a_22856_18543# a_22457_18543# a_22730_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3294 a_18291_2388# _1628_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3295 a_12150_1501# a_11711_1135# a_12065_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3296 a_2340_7497# a_1941_7125# a_2214_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3297 a_11877_8213# a_11711_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3298 vssd1 _1353_.B a_11711_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3299 a_6186_21041# _1327_.A2_N a_6185_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X3300 vccd1 a_23266_3423# a_23193_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3301 a_7013_20495# _0911_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3302 a_22549_31055# a_22015_31061# a_22454_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3304 a_25030_13469# a_24591_13103# a_24945_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3305 vssd1 _1347_.Y a_7387_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3307 a_8118_13103# _1050_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X3308 a_8818_11703# _1104_.X a_8955_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3309 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3310 a_22963_25615# a_22181_25621# a_22879_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3311 a_5537_20541# _1313_.A a_5455_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3312 vccd1 _2005_.Q a_11711_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X3313 a_2539_1501# a_1757_1135# a_2455_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3314 a_20303_26525# a_19605_26159# a_20046_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3315 vccd1 a_15963_25589# a_15879_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3316 a_11938_9839# _0992_.A2 a_11848_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3317 a_12985_2767# _1955_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3319 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3320 a_25432_10927# a_25033_10927# a_25306_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3321 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3322 vssd1 _1771_.B _2007_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3323 vccd1 a_25455_24349# a_25623_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3325 a_8887_1679# a_8105_1685# a_8803_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3327 a_12873_14337# _1038_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X3328 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_15391_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3330 vccd1 a_17749_9269# _1120_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X3331 a_20131_30186# _1481_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3332 a_23649_27247# a_22659_27247# a_23523_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3333 vssd1 _0958_.B a_21249_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3334 _0913_.A1 a_2807_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3335 _1905_.Q a_10995_19899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3336 a_17170_14735# _1090_.X a_16921_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3337 vssd1 a_13663_2741# a_13621_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3338 vccd1 _1887_.CLK a_24407_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3339 a_3993_26409# _1769_.B1 a_4248_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3340 _1316_.X a_6870_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3343 a_23239_18909# a_22457_18543# a_23155_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3345 a_25497_9839# _1927_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3346 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3347 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3348 vssd1 _1190_.X a_19899_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3349 _1764_.Y _1764_.B a_3983_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3351 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3352 vccd1 _1639_.X a_13275_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3354 vssd1 a_10643_1679# a_10811_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3355 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3356 a_25455_24349# a_24757_23983# a_25198_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3357 vssd1 a_15059_7119# a_15227_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3358 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3359 a_12396_22057# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3360 vccd1 _1194_.B2 a_12535_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3361 a_15327_3855# a_14545_3861# a_15243_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3362 vccd1 _1850_.CLK a_12539_12565# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3363 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3364 a_8286_27247# a_8109_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3365 _1020_.D1 a_15483_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3366 a_7002_5263# _1208_.A1 _1226_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X3367 a_1941_7125# a_1775_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3368 vssd1 _1116_.C1 a_15081_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3369 _1081_.D1 a_18151_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3370 _1715_.X a_27347_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3371 vccd1 a_21207_4667# a_21123_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3372 a_19952_12533# _1293_.A1 a_20175_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3373 _1870_.Q a_21115_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3374 a_19605_1135# a_19439_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3375 a_9275_24746# _1547_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3376 a_25313_21807# _1877_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3377 a_22572_15055# _1190_.B1 a_22081_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3378 a_25401_23445# a_25235_23445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3379 vssd1 fanout37.A a_18703_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3380 a_15725_7809# _1040_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X3382 a_17113_6005# _0952_.A1 a_17366_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3383 vccd1 a_25823_8207# a_25991_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3384 _1549_.A a_9223_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3386 a_22093_6575# _1582_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3387 vccd1 _1234_.A2 a_2861_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X3388 a_10865_31599# a_10699_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3389 a_15750_28335# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3390 vssd1 a_7619_26324# _1818_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3391 vccd1 a_9889_15253# a_9919_15606# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3393 _1823_.Q a_27831_20987# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3394 vccd1 a_12500_15797# _1071_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3396 vssd1 a_2807_4917# a_2765_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3399 _1308_.Y _1308_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3400 a_18049_12925# _1110_.A a_17967_12672# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3401 vccd1 a_20947_28879# a_21115_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3402 a_11558_20969# _1537_.B a_11476_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3403 vccd1 a_15151_16733# a_15319_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3404 vssd1 _0963_.B a_11313_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3405 a_2673_17231# _1249_.A2 a_2589_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3406 _1033_.B1 a_14379_9408# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3407 vccd1 _1841_.CLK a_16863_29973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3408 a_15833_23983# a_15667_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3409 vccd1 _1817_.Q a_7015_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3410 vccd1 a_5199_1403# a_5115_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3412 a_27663_21085# a_26799_20719# a_27406_20831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3413 temp1.capload\[4\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3414 a_21143_21482# _1529_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3417 a_20819_17999# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3418 a_20349_14191# _1153_.A a_20267_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3419 a_16911_1300# _1640_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3420 a_19693_15113# a_18703_14741# a_19567_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3421 _1573_.A a_14467_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3422 vssd1 a_18539_31029# a_18497_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3423 a_12150_11471# a_11711_11477# a_12065_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3425 _0983_.A2 a_14043_20513# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3426 a_5908_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3427 vssd1 a_11023_5652# _1356_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3428 vccd1 a_12467_25339# a_12383_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3429 vssd1 _1024_.A2 a_17588_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X3430 a_7465_2223# _1952_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3431 _1015_.A1 a_10167_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3434 vccd1 a_12815_19631# _1489_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3435 a_25907_8207# a_25125_8213# a_25823_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3436 a_23224_27247# a_22825_27247# a_23098_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3437 _1421_.A a_12396_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3438 a_27333_21085# a_26799_20719# a_27238_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3439 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3440 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_4324_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3441 a_13919_19200# _1900_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3442 _1283_.B1 a_2695_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X3443 a_12625_2045# a_12355_1679# a_12535_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3444 _1040_.X a_17691_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3445 a_27931_3677# a_27149_3311# a_27847_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3447 a_20429_31599# a_19439_31599# a_20303_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3448 a_15255_23060# _1545_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3449 _1412_.A a_20171_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3450 vssd1 _1924_.CLK a_21739_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3451 vccd1 _1876_.CLK a_24591_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3452 vccd1 _1050_.Y a_8031_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X3453 a_17409_6575# a_17139_6941# a_17319_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3454 a_4529_6825# a_4341_6621# a_4447_6581# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3456 vssd1 a_6835_18543# _1768_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3457 _1523_.A a_19388_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3458 a_23193_3677# a_22659_3311# a_23098_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3459 a_18049_8751# _0935_.X a_17967_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3460 a_5639_10089# _1281_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3461 vssd1 _1119_.C1 a_15633_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3462 _1242_.A2 a_7111_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3465 vccd1 a_23691_4917# a_23607_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3466 _1267_.A1 a_4739_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3467 vccd1 a_7809_18517# _1257_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3468 a_20421_17455# _1969_.Q a_20349_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3469 vssd1 _1880_.Q a_19664_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3471 a_12337_10389# a_12171_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3472 vssd1 _0952_.A2 a_23573_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3473 a_15879_32143# a_15097_32149# a_15795_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3475 a_12797_2773# a_12631_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3476 a_24113_14741# a_23947_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3477 a_9994_13763# _1422_.B a_9912_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3479 vccd1 _1090_.C a_18979_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3481 a_22369_2767# _1993_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3482 _1138_.B1 a_19439_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3483 vssd1 _1873_.CLK a_26891_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3484 a_10133_8207# _1813_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3485 a_8447_7828# _1750_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3486 a_16481_8751# _1439_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3487 vssd1 fanout33.A a_19439_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3488 _1882_.CLK a_22751_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3489 vssd1 _0918_.A a_6847_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X3492 a_4064_9615# _1177_.B a_3761_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3493 a_24301_28879# _1895_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3494 a_12276_1135# a_11877_1135# a_12150_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3495 a_18777_3855# a_18243_3861# a_18682_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3496 a_24757_5487# a_24591_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3497 a_22747_10205# a_22567_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3498 vccd1 _1474_.A_N a_12355_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3501 vccd1 _1353_.A _1332_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3502 vssd1 a_11299_12180# _1847_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3503 vssd1 a_13698_31029# a_13656_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3504 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3505 a_22687_6941# a_21905_6575# a_22603_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3506 vssd1 a_24554_28853# a_24512_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3507 vssd1 a_11858_17973# _1133_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3508 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3511 vssd1 a_4859_5162# _1365_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3512 vccd1 a_22346_5599# a_22273_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3513 _1183_.B1 a_18979_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3514 vccd1 a_27463_24251# a_27379_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3515 a_24845_25993# a_23855_25621# a_24719_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3516 vccd1 _1038_.A1 a_13304_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X3517 vccd1 _1170_.A3 a_3063_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3519 _0994_.A2 a_19275_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3521 vccd1 _0909_.A a_7015_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3522 vccd1 _1242_.A2 a_5455_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X3523 vccd1 a_8051_4667# a_7967_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3524 _1156_.Y _1156_.D a_13999_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3525 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3527 vssd1 _1223_.A2 a_2040_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3529 a_24278_11445# a_24110_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3530 vssd1 a_15963_32117# a_15921_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3531 vccd1 a_19310_1653# a_19237_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3532 vccd1 a_17923_26922# _1859_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3533 a_1945_6575# _1777_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3534 vccd1 _2004_.Q a_10865_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X3536 a_27061_2223# _1731_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3537 a_1941_4949# a_1775_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3538 vccd1 a_24903_19087# a_25071_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3539 a_19107_3855# a_18409_3861# a_18850_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3540 vccd1 _1982_.CLK a_22369_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X3541 _1590_.X a_20815_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3543 _1474_.X a_13455_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3544 vssd1 a_11030_27359# a_10988_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3546 _1041_.A1 a_26267_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3548 a_11030_3423# a_10862_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3549 a_5503_4074# io_in[5] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3550 a_15882_11471# _1118_.X a_15633_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3551 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3552 a_13599_2388# _1625_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3553 a_2915_27613# a_2217_27247# a_2658_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3554 _1234_.A1 a_2807_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3555 a_16566_9117# a_16127_8751# a_16481_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3556 a_12030_9615# _1192_.A2 a_11940_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3557 vssd1 a_17841_17601# _1049_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X3558 vccd1 a_17381_7093# _1069_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X3560 a_9669_4765# a_9135_4399# a_9574_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3562 a_15732_29967# a_15483_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3563 a_2472_19605# _1310_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3564 a_24941_2767# a_24407_2773# a_24846_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3565 _0993_.X a_16159_9867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3566 _0925_.A2 _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X3567 _1056_.B1 a_14655_23552# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3568 vssd1 a_26283_18909# a_26451_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3569 _1750_.X a_9683_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3570 a_23573_12015# a_23303_12381# a_23483_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3571 a_20046_26271# a_19878_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3573 _1334_.A1 _1325_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3574 a_17722_15823# _1028_.X a_17473_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X3575 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_9772_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3576 a_11760_24759# _1305_.B a_11902_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3578 vccd1 _1816_.CLK a_7111_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3579 a_20046_5599# a_19878_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3581 a_21909_31599# _1842_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3582 a_2765_3311# a_1775_3311# a_2639_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3583 a_12889_29973# a_12723_29973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3584 a_8378_1679# a_7939_1685# a_8293_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3585 a_27590_19743# a_27422_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3586 vccd1 _1985_.CLK a_26431_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3587 a_22707_9514# _1601_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3588 a_27548_26159# a_27149_26159# a_27422_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3590 a_20046_5599# a_19878_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3591 _1130_.C1 a_18243_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3592 a_17388_27497# a_17139_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3593 a_1775_26703# _1775_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3594 a_10229_26409# _1464_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3595 a_18601_20719# _0958_.A a_18519_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3596 a_10287_2986# _1658_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3597 a_11877_6031# _1145_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3598 _1197_.D a_14287_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X3600 a_20768_22057# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3601 a_21089_5309# a_20819_4943# a_20999_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3602 vssd1 a_22567_25071# _1873_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3604 vccd1 fanout33.A a_20083_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3606 a_4534_30511# _1329_.X a_4035_30485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X3607 a_24087_6250# _1674_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3608 a_25271_2767# a_24573_2773# a_25014_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3609 _1623_.X a_12488_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3610 a_15097_32149# a_14931_32149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3611 vccd1 _1424_.A_N a_19991_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3612 a_2287_16885# _1230_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X3613 vssd1 _1985_.CLK a_26247_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3614 a_24025_10383# _1584_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3615 vccd1 a_21115_11445# a_21031_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3616 a_24420_25993# a_24021_25621# a_24294_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3617 a_9282_16341# a_9135_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X3618 vssd1 _1029_.X _1034_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3619 vssd1 _1353_.A _1353_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3620 a_6559_26703# _1242_.B1 _1287_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X3621 a_1643_23413# _1337_.S a_1925_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X3622 _1509_.A a_20308_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3623 vccd1 a_27406_20831# a_27333_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3624 _1113_.C a_11693_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X3625 vssd1 a_2807_3829# a_2765_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3626 _0913_.A1 a_2807_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3627 a_23837_11477# a_23671_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3628 vccd1 a_20947_27791# a_21115_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3629 a_16863_21376# _1838_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3630 vccd1 a_17139_9839# _1293_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3631 _1903_.Q a_10627_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3632 fanout33.A a_16863_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3633 _1100_.X a_14747_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3634 vssd1 a_23691_9019# a_23649_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3637 a_17841_17601# _1048_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X3638 a_3329_12925# _0929_.A a_3247_12672# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3639 vccd1 _1999_.CLK a_11711_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3642 vssd1 a_27675_29588# _1860_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3643 vssd1 _0921_.B _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3644 vccd1 _2005_.Q a_11711_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X3646 _1924_.CLK a_22015_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3647 a_5389_9633# _1172_.X a_5303_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3648 a_11877_11477# a_11711_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3650 vccd1 a_6927_19087# _1269_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3652 a_10791_23552# _1855_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3653 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3654 a_15197_9661# _0935_.X a_15115_9408# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3655 vssd1 a_7755_21263# _1762_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3657 vccd1 _1764_.B a_4248_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3659 a_14369_8207# _1149_.C1 a_14287_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3660 a_25869_28879# _1342_.B _1342_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3662 vssd1 a_23047_1403# a_23005_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3665 vssd1 _1141_.C a_13485_17483# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3666 vccd1 a_16911_1300# _1945_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3667 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3668 _1050_.Y _1050_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3669 vccd1 a_26295_18218# _1970_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3670 vssd1 a_9429_15033# a_9363_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3672 vssd1 a_1657_10901# _1177_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3673 a_7573_11791# _1158_.X _1279_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3674 vccd1 _1768_.A a_8031_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3675 vccd1 _1816_.CLK a_4167_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3676 _1941_.CLK a_13643_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3677 a_27180_16367# a_26781_16367# a_27054_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3680 a_11287_27613# a_10423_27247# a_11030_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3681 a_11877_6031# _1145_.B2 a_11793_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3682 a_20522_11471# a_20083_11477# a_20437_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3683 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3684 a_19471_16395# _0939_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3685 vccd1 _1760_.X a_27167_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3686 _1804_.Y _1281_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3690 a_22273_5853# a_21739_5487# a_22178_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3691 vssd1 a_22311_26427# a_22269_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3692 a_17139_18793# _1024_.A2 a_17221_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3693 vccd1 a_8307_16367# _0935_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3694 vccd1 _1424_.A_N a_10791_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3695 vccd1 _1532_.A a_9871_10391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3696 a_1674_30511# clkbuf_0_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3697 _1970_.Q a_26267_20149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3698 a_15845_24847# _1895_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3699 a_25198_15391# a_25030_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3700 a_26965_15279# a_26799_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3702 vssd1 a_13203_10357# a_13161_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3703 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE _1306_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3704 a_18455_1501# a_17673_1135# a_18371_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3705 a_23523_4943# a_22825_4949# a_23266_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3706 vssd1 fanout37.A a_15886_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3707 a_5169_13149# _0916_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3708 a_14747_28701# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3709 a_18673_21629# _1894_.Q a_18601_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3710 _1970_.Q a_26267_20149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3711 vssd1 a_12318_1247# a_12276_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3712 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3713 a_8454_15797# a_8307_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X3714 a_13202_14441# _1038_.C1 a_13122_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3717 _1086_.Y _1086_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3719 a_12249_15279# _1433_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3720 _1207_.B1_N a_4015_8779# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3721 _1705_.A a_27807_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3724 a_25953_7663# a_25787_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3725 vccd1 _1972_.Q a_23023_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3726 _1105_.X a_17231_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3728 a_4253_20719# _1328_.S a_4035_20693# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3729 vccd1 _1841_.CLK a_16495_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3730 a_27337_27247# _1836_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3731 vssd1 _1285_.B1 a_4863_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X3732 a_9773_1135# a_9503_1501# a_9683_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3733 fanout20.X a_23303_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3735 vccd1 _1117_.B a_10327_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3736 a_9999_7119# a_9135_7125# a_9742_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3738 a_13625_31055# a_13091_31061# a_13530_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3739 vssd1 a_11711_16919# _1422_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3740 vssd1 _1985_.CLK a_26983_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3741 a_17217_27791# _1899_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3742 _1270_.A a_10423_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3743 vssd1 _0918_.A a_7481_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3745 _1291_.B2 _1234_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3746 a_24554_14709# a_24386_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3747 _1816_.CLK a_3983_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3748 vccd1 a_2823_25437# a_2991_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3749 a_22653_7663# a_22383_8029# a_22563_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3750 a_13432_27497# a_13183_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3751 vccd1 a_7571_14191# _1374_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3752 clkbuf_0_temp1.dcdel_capnode_notouch_.A temp1.dcdc.A a_15732_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3755 a_15921_32521# a_14931_32149# a_15795_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3756 a_13429_17277# _1839_.Q a_13357_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3757 vccd1 a_1737_14165# _1277_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3758 vssd1 a_25623_2491# a_25581_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3759 vssd1 a_27739_2491# a_27697_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3760 a_26141_4399# _1959_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3761 vssd1 a_15963_31029# a_15921_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3762 vccd1 _1775_.C1 a_5349_3616# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3763 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_6927_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3764 _1195_.A2 a_23691_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3765 vssd1 _1138_.C1 a_19497_18689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3766 a_25800_22729# a_25401_22357# a_25674_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3767 a_2455_6941# a_1591_6575# a_2198_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3768 a_16692_8751# a_16293_8751# a_16566_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3769 _1323_.A2 _1277_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3770 vssd1 a_2807_7093# _1273_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3771 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8215_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3772 _1018_.X a_14379_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3773 a_1941_3861# a_1775_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3774 a_3325_2767# _1951_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3775 vssd1 _0993_.X a_16300_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X3776 vccd1 _0958_.B a_18367_25099# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3777 a_23063_20175# a_22365_20181# a_22806_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3778 a_25125_13469# a_24591_13103# a_25030_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3779 a_26927_25437# a_26063_25071# a_26670_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3780 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4988_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3781 a_8569_27247# a_8392_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3783 a_25842_12533# a_25674_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X3784 vccd1 a_24703_21237# a_24619_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3785 vccd1 _1830_.CLK a_18703_14741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3787 a_3830_3971# _1448_.A a_3748_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3788 a_26965_6941# a_26431_6575# a_26870_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3789 _1456_.A a_6968_25731# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3791 a_15851_22895# _1880_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3792 a_2723_7119# a_1941_7125# a_2639_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3794 vssd1 _0921_.A a_9871_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3796 vssd1 _0974_.A2 a_20676_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3797 a_21537_30511# a_21371_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3798 vccd1 _0917_.A a_2971_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3799 vssd1 a_16267_27412# _1542_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3800 a_6835_22351# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3801 a_17231_21807# _1893_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3802 vccd1 _1941_.CLK a_20175_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3803 a_4534_23983# _1304_.B a_4035_23957# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X3804 a_17727_17999# a_16863_18005# a_17470_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3806 a_17227_4765# a_17047_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3807 a_19069_12559# _1090_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3808 vccd1 clkbuf_0_net57.X a_1674_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3809 a_26597_25437# a_26063_25071# a_26502_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3810 a_6831_5853# a_6651_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3812 a_8504_2057# a_8105_1685# a_8378_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3813 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3814 vssd1 _1073_.A2 a_16565_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3815 a_25674_12559# a_25401_12565# a_25589_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X3816 vccd1 a_20671_32143# a_20839_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3817 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_8307_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3818 a_27421_23983# a_26431_23983# a_27295_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3819 a_10417_4221# a_10147_3855# a_10327_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3821 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3822 a_22103_16733# a_21923_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3823 vssd1 a_5871_23658# _1819_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3824 a_10593_22057# _0921_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3825 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3826 a_16267_27412# _1542_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3828 _1181_.X a_15667_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X3829 vccd1 _0913_.Y temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3830 a_26183_20175# a_25401_20181# a_26099_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3831 a_19191_2767# a_18409_2773# a_19107_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3832 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A _1274_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3833 a_27456_28335# a_27057_28335# a_27330_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3834 a_5713_28111# _0913_.A1 _0913_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X3835 _0909_.C _2009_.CLK a_6099_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3836 a_20315_25834# _1531_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3837 a_2129_3311# _1798_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3838 vssd1 _1850_.CLK a_14287_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3839 vccd1 _1852_.Q a_9350_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X3840 a_10681_6825# _1189_.B2 a_10597_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3842 vssd1 a_2623_9269# a_2581_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3843 vccd1 _1177_.B _1177_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3844 vssd1 a_25455_7119# a_25623_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3845 a_5720_18543# _1242_.A1 a_5417_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3846 a_25723_3855# a_24941_3861# a_25639_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3847 a_17397_17999# a_16863_18005# a_17302_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3848 a_19439_6941# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3849 vccd1 _1841_.CLK a_17507_32149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3850 vccd1 a_5048_14165# _1249_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3851 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3852 _1631_.X a_17227_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3853 vssd1 a_9963_15939# _0987_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X3854 a_27847_10205# a_27149_9839# a_27590_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3855 vssd1 a_24703_11445# a_24661_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3856 vssd1 _1218_.B _1301_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X3857 a_2281_31751# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3858 a_15097_31061# a_14931_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3859 vccd1 a_26175_26427# a_26091_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3860 a_5692_15253# _1325_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3863 _1730_.X a_23759_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3864 vccd1 a_18371_32143# a_18539_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3867 vccd1 _1113_.C a_17231_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3868 vssd1 a_28015_19899# a_27973_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3869 vccd1 a_7258_1247# a_7185_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3870 a_22369_26703# _1839_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3871 vssd1 _1880_.CLK a_23947_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3872 a_10279_16911# a_10667_16885# _1141_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3873 a_11793_21583# _1904_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3874 vccd1 _1982_.CLK a_26431_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3875 a_24941_16367# a_24775_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3876 a_10133_6031# _1563_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3878 a_23013_27247# _1893_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X3879 a_15698_18115# _1405_.B a_15616_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3880 vssd1 a_13551_8215# _1010_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3881 a_17996_24233# _1134_.B1 a_17894_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X3883 a_5233_11445# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3885 a_2382_3423# a_2214_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3886 vccd1 a_25455_1501# a_25623_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3887 vssd1 _1090_.C a_18305_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3891 a_26057_30287# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3894 vssd1 _1313_.X _1786_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3895 vccd1 a_20131_21972# _1889_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3896 a_10791_13647# _0987_.B _1071_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3897 a_25769_24527# a_25235_24533# a_25674_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3899 a_3548_20175# _1282_.A2 a_3087_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X3900 a_8027_19997# a_7847_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3902 vssd1 a_11306_31711# a_11264_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3903 _1101_.X a_13275_17024# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3904 a_13183_11177# _1197_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3905 a_25539_7119# a_24757_7125# a_25455_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3906 _1091_.B1 a_15207_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3907 vssd1 _1050_.Y a_8289_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X3909 vssd1 _1876_.Q a_18560_22467# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3910 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3911 vccd1 a_13311_25615# a_13479_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3912 a_8215_7119# _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3913 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_6736_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3915 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3916 vssd1 a_16274_24095# a_16232_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3917 vssd1 _0981_.B a_14901_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3919 a_15235_10205# a_14453_9839# a_15151_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3920 a_2122_9839# a_1945_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3921 vccd1 a_23707_29967# a_23875_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3922 vssd1 _1311_.B1 a_1644_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X3923 vccd1 _1301_.A1 a_3681_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3924 a_2313_25071# _1767_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3925 vssd1 _0975_.X a_15575_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3926 a_13161_10761# a_12171_10389# a_13035_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3927 a_13275_31965# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3928 _1198_.A1 a_6303_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3929 vccd1 a_4627_6031# _1782_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3930 a_17493_29423# _1475_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3931 vccd1 a_5693_16341# _1267_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3932 _1024_.A2 a_17541_15307# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X3933 vssd1 _1108_.C1 a_13517_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X3934 a_3835_2767# a_3137_2773# a_3578_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3935 a_2103_31573# _1329_.A1 a_2330_31921# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X3936 vccd1 a_13698_31029# a_13625_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3938 _1056_.C1 a_15851_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3939 a_18642_8323# _1577_.B a_18560_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3940 _1082_.X a_14379_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X3941 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3942 _2008_.Q a_3083_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3944 vssd1 a_27038_6687# a_26996_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3945 vccd1 a_21407_8029# a_21575_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3946 vssd1 a_14894_30623# a_14852_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3947 vssd1 _0958_.B a_16649_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3948 _1281_.A1 a_2807_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3949 a_20479_30877# a_19697_30511# a_20395_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3950 vccd1 a_20303_29789# a_20471_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3951 a_25382_16479# a_25214_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X3953 vccd1 _1043_.B a_9442_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X3954 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13432_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3955 vccd1 a_14979_17130# _1821_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3956 a_11601_2223# a_11435_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3957 a_23523_11293# a_22659_10927# a_23266_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3958 a_25674_12559# a_25235_12565# a_25589_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3959 a_6230_25321# _1242_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X3960 a_13643_22464# _1899_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3961 a_22227_26525# a_21445_26159# a_22143_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3962 a_9970_26742# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3966 _1821_.Q a_19735_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3968 vccd1 a_27590_12127# a_27517_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3970 vssd1 _2009_.CLK a_2603_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3971 a_20004_31599# a_19605_31599# a_19878_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3972 a_15921_25993# a_14931_25621# a_15795_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3974 a_14563_29967# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3975 vssd1 _1240_.X a_1643_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X3976 vccd1 _1816_.CLK a_7019_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3977 vssd1 a_11023_26922# _1858_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3978 _1852_.Q a_12467_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3979 vssd1 _0909_.B a_5731_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3981 vccd1 a_25198_13215# a_25125_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X3982 io_out[1] a_1643_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3983 vccd1 _1761_.X a_3514_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3984 vccd1 _2023_.CLK a_1775_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3985 _1897_.Q a_20471_31867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3986 a_23193_11293# a_22659_10927# a_23098_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3988 a_12079_12381# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3989 a_27663_21085# a_26965_20719# a_27406_20831# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3990 vssd1 a_24830_15797# a_24788_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3991 a_16565_3311# a_15575_3311# a_16439_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3993 vssd1 a_16734_8863# a_16692_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3994 vccd1 _1775_.C1 a_1683_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3995 a_8615_25953# _0911_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3996 vccd1 a_11115_7828# _1614_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3999 a_24087_6250# _1674_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4000 _1242_.A1 a_2623_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4001 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4002 a_12502_15391# a_12334_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4003 _1184_.X a_19439_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4004 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4006 vccd1 _1132_.C a_13643_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4007 vccd1 _1459_.A a_21187_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4008 a_6817_1135# a_6651_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4009 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4010 vssd1 _1342_.Y a_7755_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4011 vccd1 _1141_.C a_11895_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4012 vssd1 a_2807_6005# _1255_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4013 a_16986_25731# _1484_.B a_16904_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4014 vssd1 a_6705_16341# _1789_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4015 a_27437_14013# a_27167_13647# a_27347_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4016 vccd1 a_27859_29098# _1855_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4018 a_14839_26159# _0966_.B1 a_15017_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4022 a_9323_13103# _1198_.B2 a_9186_13255# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4023 vccd1 fanout21.X a_24775_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4024 a_15036_3145# a_14637_2773# a_14910_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4025 vssd1 _1179_.B1 a_16208_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X4026 a_2723_6031# a_1941_6037# a_2639_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4027 a_7387_31965# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4028 a_11563_31965# a_10699_31599# a_11306_31711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4029 _1837_.Q a_24887_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4030 vssd1 _1979_.Q a_22572_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X4031 a_14328_3561# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4032 a_2125_25071# a_1959_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4033 a_10515_19407# _0921_.A a_10765_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4034 a_19189_13985# _0958_.A a_19103_13985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4035 a_11752_13353# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4038 a_19204_28995# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4039 a_1965_19087# _1764_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4041 a_10317_19631# _1557_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4043 a_25581_5487# a_24591_5487# a_25455_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4044 a_5578_9001# _1279_.A1 a_5496_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4045 a_17305_29423# a_17139_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4046 a_16307_6941# a_16127_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4048 a_15630_29535# a_15462_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4049 a_7185_1501# a_6651_1135# a_7090_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4050 _1837_.Q a_24887_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4052 a_23115_19087# a_22935_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4053 a_24945_13103# _1980_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4054 _1286_.A1 a_2623_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4056 a_23377_16917# a_23211_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4057 a_12318_11445# a_12150_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4058 vccd1 _0952_.A2 a_23483_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4059 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4060 vccd1 _0958_.A a_18519_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4061 vccd1 _1459_.A a_16035_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4062 vssd1 a_15887_29789# a_16055_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4063 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4064 vccd1 a_1643_21237# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4065 a_17809_20513# _0958_.A a_17723_20513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4066 a_15483_13760# _1019_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4067 a_7636_32143# a_7387_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4068 vssd1 _1876_.CLK a_24591_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4069 vccd1 a_23395_17455# _1887_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4070 a_14287_13353# _1120_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4072 vssd1 _0903_.C _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4073 a_11233_31965# a_10699_31599# a_11138_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4074 _0951_.B _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4075 vssd1 a_24887_25589# a_24845_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4076 a_26099_4943# a_25235_4949# a_25842_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4077 a_17691_8320# _1040_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4079 vssd1 _1859_.Q a_7473_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4080 vccd1 _1249_.A1 a_2047_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4081 a_22081_14709# _1190_.B1 a_22238_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4082 vssd1 _1091_.C1 a_16921_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X4083 _1876_.CLK a_21831_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4084 vccd1 _1887_.Q a_17352_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4085 _1830_.Q a_19735_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4086 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4087 vccd1 a_21327_20394# _1888_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4090 vccd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4091 a_12150_11471# a_11877_11477# a_12065_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4092 vccd1 _1841_.CLK a_17507_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4093 _1609_.X a_16307_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4094 vssd1 a_22935_10383# fanout24.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4095 a_27149_26159# a_26983_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4096 a_19470_8323# _1577_.B a_19388_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4097 vccd1 _1140_.C a_12295_20747# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4098 _1144_.B a_4003_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4099 _1038_.A1 a_12743_13621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4101 vssd1 a_27295_24349# a_27463_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4103 _1767_.B a_4587_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4104 a_21327_20394# _1521_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4106 vccd1 a_22063_9514# _1578_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4107 _1038_.A1 a_12743_13621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4108 a_13238_2741# a_13070_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4110 a_14637_2773# a_14471_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R6 vccd1 temp1.capload\[13\].cap_43.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4111 a_21549_3311# a_21279_3677# a_21459_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4112 _1261_.A1 a_2715_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4114 vccd1 _1127_.A a_20267_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4115 vccd1 a_16083_14954# _1831_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4116 vccd1 _1132_.C a_15483_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4117 a_4244_30511# a_4213_30663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X4118 _1570_.X a_11752_13353# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4119 _1270_.Y temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4120 a_19928_18793# _1138_.B1 a_19826_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4121 vccd1 _1075_.C a_18427_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4122 vssd1 _1133_.C a_20421_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4127 vssd1 a_18355_28853# a_18313_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4128 _0906_.X a_8213_25335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X4129 a_23983_8207# a_23285_8213# a_23726_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4130 a_2405_27247# _2003_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4131 a_22238_13647# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4133 a_27167_12559# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4134 a_11874_25437# a_11601_25071# a_11789_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4135 _0909_.A _0903_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4136 a_13432_28879# a_13183_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4138 a_24554_14709# a_24386_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4139 a_8031_13353# _1052_.B1 _1324_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X4140 a_22270_29789# a_21997_29423# a_22185_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4142 _1141_.C _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4143 _1040_.B a_26175_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4145 a_23579_13469# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4146 vssd1 a_23799_3855# a_23967_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4147 vssd1 a_7699_3855# a_7867_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4148 temp1.capload\[3\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4149 a_19562_17705# _1506_.B a_19480_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4150 a_9400_13353# _1187_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X4151 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4152 a_9284_21781# a_9135_21807# a_9580_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4153 a_4627_18543# _1326_.A2 a_4533_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4154 vccd1 _1985_.CLK a_24775_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4155 a_24757_13103# a_24591_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4156 _1869_.Q a_22863_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4158 vssd1 _0965_.A2 a_15277_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4160 vssd1 a_12318_11445# a_12276_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4161 a_5908_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4162 a_16014_3677# a_15741_3311# a_15929_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4163 _1828_.Q a_23783_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4165 vccd1 a_9282_16341# _1090_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4166 vccd1 a_23266_11039# a_23193_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4167 _1261_.A2 a_8615_25953# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4168 a_25842_16885# a_25674_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4169 a_24386_14735# a_24113_14741# a_24301_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4170 a_7473_30333# a_7203_29967# a_7383_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4171 _1762_.Y _1764_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4172 a_26099_16911# a_25401_16917# a_25842_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4174 a_2778_15529# _1219_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4175 a_12065_1135# _1612_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4176 a_22879_25615# a_22015_25621# a_22622_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4177 vssd1 _1782_.A a_1816_11587# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4178 vssd1 a_24039_12559# _1985_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4179 _1828_.Q a_23783_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4184 vccd1 a_5692_15253# _1291_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X4185 vccd1 a_22879_1501# a_23047_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4186 a_22825_4949# a_22659_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4187 a_3993_26409# _1775_.C1 _1769_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4188 a_7828_6351# a_7295_6031# _1177_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4189 a_1820_10927# _1170_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X4190 vssd1 a_2807_3579# a_2765_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4191 a_17730_4943# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4192 a_2594_31055# clkbuf_0_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4193 vssd1 _1179_.B2 a_19480_15529# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4195 _0930_.A a_6559_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4196 a_2220_19087# _1257_.X a_1965_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4197 a_13238_2741# a_13070_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4198 vccd1 a_26267_23413# a_26183_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4199 _0951_.B a_10814_14709# a_10594_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4200 a_26387_1898# _1650_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4201 vssd1 a_10073_20693# a_10007_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4202 vccd1 a_2623_6843# a_2539_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4203 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4204 a_20492_20291# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4205 a_2048_19407# _0922_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X4206 a_24662_15823# a_24223_15829# a_24577_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4207 vssd1 a_27406_15391# a_27364_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4209 a_2582_1679# a_2143_1685# a_2497_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4210 a_26007_26525# a_25309_26159# a_25750_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4211 a_22549_25615# a_22015_25621# a_22454_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4212 vccd1 _1850_.CLK a_11895_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4213 vssd1 a_9871_10391# _1537_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4214 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4215 a_1841_23759# _1270_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4217 vssd1 _1086_.A a_6835_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4219 a_16106_24349# a_15833_23983# a_16021_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4220 a_26870_24349# a_26597_23983# a_26785_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4221 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4222 vssd1 a_25363_9295# a_25531_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4225 vssd1 a_10839_20884# _1851_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4226 _1216_.A2 _1246_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4227 a_24811_28879# a_24113_28885# a_24554_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4228 a_14776_24233# _0983_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X4229 a_25271_17999# a_24573_18005# a_25014_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4231 a_2769_27797# a_2603_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4232 vccd1 _1690_.A_N a_22015_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4234 _1483_.A a_16904_25731# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4235 vccd1 a_19027_25834# _1894_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4236 a_12123_23805# _1305_.B a_11760_23671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4237 _1697_.A a_23115_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4238 a_2673_13103# a_1683_13103# a_2547_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4239 vssd1 a_21407_8029# a_21575_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4240 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7636_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4241 _1232_.Y a_9963_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4242 vssd1 _1999_.CLK a_11711_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4243 _1636_.A a_18147_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4244 vssd1 a_20947_28879# a_21115_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4245 _1625_.X a_13408_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4246 vccd1 a_11306_31711# a_11233_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4247 a_17811_27791# a_17029_27797# a_17727_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4248 vssd1 _1999_.CLK a_9135_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4249 a_5261_10973# _0917_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4250 vssd1 _1887_.CLK a_25235_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4251 a_21905_5487# a_21739_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4252 vccd1 _0956_.C a_11693_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X4253 a_23119_14557# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4254 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_6651_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4255 _2004_.Q a_3635_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4256 _1219_.B1 a_7201_14851# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4257 vccd1 _1240_.B1 a_3299_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4259 vccd1 a_12318_8181# a_12245_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4260 a_19027_25834# _1534_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4261 a_18673_20719# _1837_.Q a_18601_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4262 a_20437_27791# _1875_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4263 a_4525_20175# _1327_.A1_N a_4443_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4264 a_22383_13469# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4265 vssd1 _1816_.CLK a_4167_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4266 a_19793_26159# _1542_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4267 a_16182_3423# a_16014_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4268 a_2589_17231# _1249_.A1 a_2287_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X4269 a_26854_14303# a_26686_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4271 a_2962_14735# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4272 vssd1 fanout33.A a_15667_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4273 vssd1 a_17727_17999# a_17895_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4274 _0975_.X a_18887_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X4275 vssd1 _1822_.Q a_20860_19203# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4276 _1532_.A a_2327_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4277 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4278 vssd1 a_15335_2767# a_15503_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4279 vccd1 a_27571_2589# a_27739_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4280 vccd1 _1860_.CLK a_9963_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4281 vssd1 a_25899_11195# a_25857_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4282 a_20690_11445# a_20522_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4283 a_22419_31965# a_21721_31599# a_22162_31711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4284 _0965_.A2 a_16159_20747# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4286 vccd1 a_23903_1300# _1991_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4288 vssd1 a_22015_7119# _1924_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4290 _1308_.B _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4292 a_12659_1501# a_11877_1135# a_12575_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4293 vccd1 a_9999_4765# a_10167_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4294 _1059_.X a_15299_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X4295 a_19605_29423# a_19439_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4296 a_27057_28335# a_26891_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4297 a_3111_5652# io_in[6] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4298 a_18551_11809# _1127_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4299 _1844_.Q a_20655_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4300 vccd1 a_17527_26427# a_17443_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4301 a_3553_13647# _1246_.A3 _1247_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.305 ps=1.61 w=1 l=0.15
X4302 a_25355_2767# a_24573_2773# a_25271_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4304 a_1735_29941# _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X4306 a_4244_23983# a_4213_24135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X4309 a_22567_10205# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4310 _1052_.B1 _1084_.C1 a_10331_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4311 a_19807_16911# _1179_.B1 a_19985_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4312 a_13445_31055# _1856_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4313 a_18509_15279# _1127_.A a_18427_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4314 _1479_.A a_14743_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4317 vssd1 _1027_.X a_17473_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X4318 a_12299_2589# a_11435_2223# a_12042_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4319 vccd1 a_21235_1898# _1992_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4322 a_12570_26409# _1422_.B a_12488_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4323 a_11299_11092# _1438_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4324 a_13974_21237# a_13806_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4325 _1279_.A1 _1164_.A2 a_7656_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4326 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13432_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4328 a_27663_15645# a_26799_15279# a_27406_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4329 a_25198_5599# a_25030_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4331 a_4064_21583# _1312_.B1 a_3759_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4332 a_4314_7093# a_4146_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4333 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4334 a_17470_29941# a_17302_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4338 vssd1 io_in[0] a_2962_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4339 a_22454_1679# a_22181_1685# a_22369_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4340 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4341 _0966_.X a_14839_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X4342 a_17381_14337# _1032_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X4344 vccd1 a_14491_24501# a_14407_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4345 vccd1 a_27095_23163# a_27011_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4346 a_22457_18543# a_22291_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4347 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4348 vssd1 a_21143_23658# _1833_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4349 vssd1 _1113_.C a_18673_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4350 a_27333_15645# a_26799_15279# a_27238_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4351 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4352 a_10331_23145# _0983_.B1 a_10413_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4353 vccd1 a_15633_19061# _1020_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X4354 vssd1 a_5417_18517# _1254_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4356 a_9761_22357# a_9595_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4357 a_6847_22057# _0921_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4358 vssd1 _1090_.C a_19133_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4359 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4360 vssd1 _2023_.CLK a_3707_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4361 a_14594_24233# _1056_.D1 a_14345_24129# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4362 a_4558_22895# _1284_.B1 a_4263_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X4363 vccd1 _1907_.CLK a_9135_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4366 a_27330_11293# a_26891_10927# a_27245_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4367 vccd1 _2009_.CLK a_2603_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4368 vssd1 _0918_.A _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X4369 a_18519_14191# _1696_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4370 vccd1 _1590_.A_N a_17967_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4371 fanout28.A a_1591_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4372 a_20230_28447# a_20062_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4373 _1332_.Y _1353_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4375 a_2309_7119# a_1775_7125# a_2214_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4377 vccd1 a_11759_29098# _1429_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4378 _1151_.X a_21463_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4379 a_25033_10927# a_24867_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4380 a_9970_27069# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4381 _1133_.C a_11858_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4382 a_26479_11690# _1715_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4383 vccd1 a_11287_3677# a_11455_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4384 vccd1 a_13495_2767# a_13663_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4385 vccd1 _0935_.X a_14839_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4386 a_9602_25981# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4387 vccd1 _1907_.CLK a_6283_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4388 vssd1 a_12927_4917# a_12885_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4389 a_14809_23805# _1874_.Q a_14737_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4390 vccd1 a_5503_4074# _0917_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4391 a_25156_27247# a_24757_27247# a_25030_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4392 a_13999_11471# _1156_.C a_13805_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4394 a_25401_16917# a_25235_16917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4397 vssd1 _1941_.CLK a_16863_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4398 vccd1 _1171_.Y a_7742_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X4399 vssd1 a_20690_11445# a_20648_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4400 vccd1 a_25750_9951# a_25677_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4401 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4402 a_6559_4943# _1202_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4403 a_3801_28981# _0909_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X4405 vssd1 _1123_.X a_6467_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X4406 _1074_.C a_9195_17973# a_8807_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4407 _1890_.Q a_27463_17723# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4408 a_2708_2057# a_2309_1685# a_2582_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4409 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4410 a_13533_21269# a_13367_21269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4411 a_10827_19997# a_10129_19631# a_10570_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4412 a_8706_17027# _1313_.X a_8624_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4413 a_25309_3855# a_24775_3861# a_25214_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4414 vssd1 _0921_.B _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4415 _1198_.B2 a_13183_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4416 vccd1 a_26267_22325# a_26183_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4417 vssd1 _1967_.Q a_21181_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4418 vccd1 _1249_.A1 _1265_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4419 a_12245_8207# a_11711_8213# a_12150_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4420 a_6743_10703# _1324_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4421 a_17578_29789# a_17305_29423# a_17493_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4422 a_13403_12559# a_12705_12565# a_13146_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4423 vssd1 _0925_.A2 a_4789_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4425 a_2547_8029# a_1849_7663# a_2290_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4426 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_17316_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4427 _1389_.A a_23483_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4428 a_4709_13647# _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X4429 a_1945_2223# _1793_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4430 vccd1 _1139_.C a_11711_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4431 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5816_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4432 a_16481_8751# _1439_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4434 vccd1 a_12815_9295# _1459_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4435 _1223_.A2 _1219_.A2 a_13257_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X4436 vccd1 _1234_.A1 a_6559_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4437 vccd1 a_3175_1653# a_3091_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4438 vccd1 _1047_.C a_15607_12043# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4439 a_7176_27497# a_6927_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4440 vccd1 _1374_.A_N a_23211_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4441 vssd1 a_5455_14735# _1231_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4442 vccd1 a_22339_19796# _1968_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4443 _1529_.A a_20860_19881# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4445 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4446 vccd1 _2005_.Q a_9195_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X4447 a_9602_15279# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4448 vssd1 _1982_.CLK a_26431_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4449 vssd1 a_25623_7093# a_25581_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4451 a_19041_19453# _1882_.Q a_18969_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4453 a_21695_17620# _1391_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4454 a_19973_16911# _1968_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4455 vccd1 a_26267_4917# a_26183_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4456 _1752_.X a_7659_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4457 a_13488_9001# _1057_.X a_13386_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4458 vccd1 a_7479_28887# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4459 a_18107_14954# _1574_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4460 vssd1 _1242_.A2 a_5713_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X4461 _1519_.A a_21091_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4465 _1540_.A a_14927_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4466 a_23098_9117# a_22659_8751# a_23013_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4468 vccd1 a_6151_22869# _1282_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X4469 a_25398_22173# a_24959_21807# a_25313_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4470 a_22983_19796# _1385_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4471 vccd1 _1822_.Q a_20942_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4472 a_17060_31599# a_16661_31599# a_16934_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4474 _1210_.B _1162_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4475 vssd1 a_20315_25236# _1838_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4477 a_10546_1385# _1607_.B a_10464_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4478 a_16408_5487# _0997_.X a_15917_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4479 a_14103_6031# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4480 vccd1 a_6927_19087# _1269_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4481 a_7366_15279# a_7189_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4482 _1308_.B a_9871_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4483 vccd1 _0935_.X a_18795_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4484 vccd1 a_23047_24501# a_22963_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4485 vssd1 a_2547_13469# a_2715_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4486 vccd1 a_8102_30511# a_8208_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4487 vccd1 a_10459_29789# a_10627_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4488 vccd1 _1273_.A1 a_4248_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4489 _1033_.A1 a_25623_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4490 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4491 vssd1 _1353_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4493 _1759_.A a_8947_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4494 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4495 vccd1 _1068_.A1 a_13120_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X4497 a_15235_30877# a_14453_30511# a_15151_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4498 _1375_.A a_8855_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4499 a_27379_6941# a_26597_6575# a_27295_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4500 a_10344_30345# a_9945_29973# a_10218_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4501 vssd1 _1830_.CLK a_15794_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4502 a_22244_13967# _1032_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X4503 a_11759_1898# _1662_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4504 a_14467_11293# a_14287_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4505 a_8464_32143# a_8215_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4506 _1243_.A _1242_.B1 a_5087_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4507 _1310_.B1 a_7481_23555# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4508 vssd1 _1889_.Q a_22285_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4509 a_2706_21583# _1259_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4510 a_26394_7775# a_26226_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4511 _1055_.C a_12027_20495# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X4512 a_19654_15823# _1130_.D1 a_19405_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X4515 vccd1 a_2715_13371# _1218_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4516 vccd1 a_23523_27613# a_23691_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4517 vssd1 _1893_.Q a_17548_25321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4518 vccd1 a_27406_15391# a_27333_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4519 a_25497_3311# _1990_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4521 _1717_.X a_23667_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4522 a_10839_20884# _1443_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4524 _1594_.X a_17456_7913# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4525 a_9761_29423# a_9595_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4526 a_26394_7775# a_26226_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4528 a_4337_1679# _1649_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4529 a_18751_5162# _1594_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4530 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7728_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4532 a_14972_26819# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4533 a_25582_26525# a_25309_26159# a_25497_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4534 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4535 vccd1 a_26099_20175# a_26267_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4536 _1850_.CLK a_2235_2775# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4537 a_25539_21085# a_24757_20719# a_25455_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4538 vccd1 a_22879_2767# a_23047_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4539 _1607_.X a_18468_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4542 a_25030_17821# a_24591_17455# a_24945_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4544 a_12425_25071# a_11435_25071# a_12299_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4545 a_5449_22895# _1306_.X a_5231_22869# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4546 a_21844_26159# a_21445_26159# a_21718_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4548 vssd1 a_26099_20175# a_26267_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4549 a_6277_11177# _1316_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X4550 vssd1 a_5015_1653# a_4973_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4551 a_17217_29967# _1477_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4552 a_27859_30186# _1456_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4553 a_18291_2388# _1628_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4554 vssd1 _1474_.B a_13545_32509# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4556 a_4968_28879# a_4719_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4557 a_14461_18793# _1082_.D a_14379_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X4558 vssd1 a_16607_3579# a_16565_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4559 vccd1 _1459_.A a_12815_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4560 vccd1 _1293_.A1 a_8859_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4561 _1246_.A2 _1226_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4562 _1398_.X a_15479_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4563 vccd1 _1170_.B2 _1205_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4564 vssd1 _1086_.A _1086_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4565 vccd1 a_25455_28701# a_25623_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4566 _1898_.Q a_20471_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4567 a_19991_24349# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4568 vssd1 a_7159_20884# _1557_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4569 a_12989_18543# _0964_.A a_12907_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4570 vccd1 _1308_.B a_2009_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4571 a_7980_9411# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4572 a_5693_19605# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X4574 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9595_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4575 a_24646_19061# a_24478_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4576 a_12575_29789# a_11711_29423# a_12318_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4579 vssd1 a_9135_25071# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4581 vssd1 a_9999_4765# a_10167_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4582 a_18877_7485# _0935_.X a_18795_7232# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4584 a_17647_2388# _1637_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4585 a_6817_1135# a_6651_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4586 _1270_.A _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4587 a_2309_6031# a_1775_6037# a_2214_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4589 a_25033_10927# a_24867_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4590 vccd1 _1448_.A a_8215_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4591 vssd1 _0987_.Y a_10953_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X4593 _1422_.B a_11711_16919# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4594 vssd1 _1816_.CLK a_2143_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4596 vssd1 _1856_.Q a_6968_25731# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4597 a_7481_23555# _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4598 vccd1 a_4571_7119# a_4739_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4600 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4601 _1771_.B a_2471_22869# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4602 _1703_.A a_27623_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4603 a_16127_16617# _1070_.A2 a_16209_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4604 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4605 _1070_.X a_17139_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4607 _1116_.D1 a_13183_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4608 _1081_.C1 a_21095_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4609 a_19439_12015# _1135_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4610 temp1.capload\[10\].cap.Y temp1.capload\[10\].cap.A a_14373_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4611 a_12245_29789# a_11711_29423# a_12150_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4612 _1374_.A_N a_7571_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4613 a_25581_31599# a_24591_31599# a_25455_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4614 a_2214_4765# a_1775_4399# a_2129_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4615 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4616 a_9037_19087# _0925_.A2 _1234_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4617 a_8300_25077# a_8113_25117# a_8213_25335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4618 _1972_.Q a_25623_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4619 a_19439_19997# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4620 a_22285_19453# a_22015_19087# a_22195_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4621 _0985_.A a_19807_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X4622 a_1945_9295# _1780_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4623 a_2009_21263# _0923_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.585 pd=2.17 as=0.135 ps=1.27 w=1 l=0.15
X4624 vssd1 a_14399_21237# a_14357_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4625 a_12570_4649# _1607_.B a_12488_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4626 temp1.capload\[13\].cap.Y temp1.capload\[13\].cap_43.LO a_23297_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4628 a_19605_5487# a_19439_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4630 a_12600_16367# a_12557_16600# a_12528_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X4631 _1590_.A_N a_16035_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4632 vssd1 _1762_.A a_9747_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X4633 vssd1 _1194_.A2 a_13408_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4634 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7176_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4636 vssd1 a_27647_16635# a_27605_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4637 a_16934_26525# a_16495_26159# a_16849_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4639 vccd1 a_27463_17723# a_27379_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4640 vccd1 clkbuf_0_net57.X a_1674_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4641 vssd1 a_15243_4943# a_15411_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4643 a_23650_23439# a_23211_23445# a_23565_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4644 a_20676_10499# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4645 a_4709_13647# _1217_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X4646 a_1975_29967# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X4648 a_8009_4399# a_7019_4399# a_7883_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4651 a_12189_24825# _1287_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4652 a_27149_26159# a_26983_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4653 a_3884_29239# _0909_.A a_3801_28981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4654 _0966_.A2 a_18367_25099# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4655 a_23473_8207# _1916_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4656 a_21917_9839# a_21647_10205# a_21827_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4657 a_14287_9001# _1196_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X4659 a_8941_6397# _1293_.A1 a_8859_6144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4660 a_20414_32117# a_20246_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4661 vccd1 _0921_.A a_10593_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4662 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4663 vssd1 a_19735_17973# a_19693_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4664 vccd1 a_21407_23261# a_21575_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4665 a_24025_21263# _1691_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4666 a_26099_20175# a_25235_20181# a_25842_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4667 vccd1 a_2991_25339# _2005_.Q vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4668 vssd1 _1899_.Q a_11476_20969# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4669 _1781_.B _1775_.A2 a_7013_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4670 a_23224_8751# a_22825_8751# a_23098_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4671 vssd1 a_6559_9295# _0930_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4672 _1177_.Y _1177_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4673 _1764_.A a_6927_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4674 a_27422_5853# a_27149_5487# a_27337_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4675 vccd1 _0984_.A2 a_12153_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4676 a_10865_18909# _2005_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X4677 a_20521_30511# a_19531_30511# a_20395_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4679 a_19310_14709# a_19142_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4680 _1544_.A_N a_8307_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4681 vccd1 _1010_.A a_11343_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4682 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8464_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4684 a_4149_1685# a_3983_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4686 _1649_.A a_7704_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4689 _0987_.B a_9963_15939# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4690 vccd1 _1830_.CLK a_22050_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4691 vssd1 _1329_.S a_2602_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X4692 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_7479_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4694 vccd1 a_2327_20183# _1775_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4695 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_10791_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4696 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_4811_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4697 vccd1 _1528_.A a_20942_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4698 vccd1 _1723_.A_N a_23487_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4699 a_22695_29789# a_21997_29423# a_22438_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4700 vccd1 a_12467_2491# a_12383_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4701 a_14287_11293# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4702 vssd1 a_17923_26922# _1859_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4703 a_21407_23261# a_20709_22895# a_21150_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4704 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4706 a_19142_14735# a_18869_14741# a_19057_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4707 _1743_.A a_20263_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4708 a_16566_9117# a_16293_8751# a_16481_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4709 _1881_.Q a_26175_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4710 a_11907_20175# _2004_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X4711 a_7650_17277# _1269_.A1 a_7561_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4712 vssd1 _1985_.CLK a_24775_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4714 _1156_.C a_11711_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4715 a_27548_19631# a_27149_19631# a_27422_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4716 a_18243_12015# _1128_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4717 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4718 a_21032_15823# _1081_.B1 a_20930_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4719 a_19623_7119# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4720 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4721 a_22963_2767# a_22181_2773# a_22879_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4722 a_12042_2335# a_11874_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4724 _1040_.B a_26175_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4725 _2019_.D a_4613_3916# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X4726 a_9999_31055# a_9135_31061# a_9742_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4727 _1786_.A1 _1313_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4728 vccd1 a_22622_1653# a_22549_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4729 a_20982_2589# a_20543_2223# a_20897_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4730 vssd1 _2006_.Q a_9894_17429# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4732 a_7479_28585# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4733 a_25497_29423# _1880_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4734 vssd1 a_23523_9117# a_23691_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4735 vssd1 a_24979_28853# a_24937_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4736 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4737 _1447_.A a_9268_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4738 vssd1 _0918_.A _0922_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4739 vccd1 a_12502_15391# a_12429_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4740 vssd1 _0983_.B1 a_14920_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X4741 a_11299_11092# _1438_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4742 a_4341_6621# _1210_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4743 a_22063_22570# _1509_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4744 a_15962_19087# _1018_.X a_15882_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X4745 _1800_.A2 _1317_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4746 a_21827_10205# a_21647_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4747 a_9669_31055# a_9135_31061# a_9574_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4748 vccd1 _1234_.A1 a_9037_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4749 _1089_.B a_21207_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4751 _1555_.A a_7935_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4752 a_27146_2589# a_26873_2223# a_27061_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4753 a_27590_12127# a_27422_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4754 a_27347_12559# a_27167_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4755 a_6553_17705# _1234_.A2 _1267_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4756 vssd1 _1850_.CLK a_11895_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4757 vccd1 _1782_.A a_7479_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4758 vssd1 _1287_.A fanout12.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4759 a_2382_4917# a_2214_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4760 a_21810_30877# a_21371_30511# a_21725_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4761 vssd1 a_27663_22173# a_27831_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4762 vccd1 _1890_.Q a_19562_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4764 a_4531_2589# a_4351_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4765 vssd1 _1177_.C a_4064_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4766 vssd1 a_27923_28603# a_27881_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4767 a_10791_13647# _1010_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4768 a_18409_3861# a_18243_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4770 vccd1 _1141_.C a_18243_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4772 a_25539_31965# a_24757_31599# a_25455_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4774 _1788_.X a_8624_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4775 a_21042_16617# _1113_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X4776 vssd1 _1793_.A2 a_8301_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4777 a_25401_13653# a_25235_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4778 a_19885_30511# _1871_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4781 vccd1 a_12318_29535# a_12245_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4783 a_19069_12559# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4784 _1760_.X a_2309_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X4785 vccd1 _1761_.X a_3514_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4788 a_13264_6575# _1068_.A1 a_12689_6721# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X4789 a_27422_10205# a_26983_9839# a_27337_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4790 vccd1 a_20471_26427# a_20387_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4791 vccd1 _1856_.Q a_7050_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4792 vccd1 _0906_.X a_7479_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4793 a_22063_8426# _1580_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4794 a_2281_31751# _1329_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X4796 vssd1 a_25823_8207# a_25991_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4797 a_24945_27247# _1835_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4798 a_8464_26409# a_8215_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4799 vccd1 a_23231_20149# a_23147_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4800 vccd1 _1040_.B a_21183_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4801 a_10229_26159# _1818_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4803 a_19671_25834# _1496_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4804 _1029_.B1 a_14747_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X4806 a_7101_14735# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4807 vssd1 a_12299_25437# a_12467_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4809 vccd1 _1344_.B a_4627_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4811 vssd1 a_20211_31055# a_20379_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4813 a_2340_4399# a_1941_4399# a_2214_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4814 a_23285_8213# a_23119_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4815 a_13449_22895# _0961_.A a_13367_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4817 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4818 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4819 vccd1 a_10811_29941# a_10727_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4820 a_8944_28111# _1347_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4821 vccd1 a_11711_15831# _1424_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4822 vssd1 a_25531_9269# a_25489_9673# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4824 a_27422_27613# a_26983_27247# a_27337_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4826 a_10160_29423# a_9761_29423# a_10034_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4827 a_25125_24349# a_24591_23983# a_25030_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4829 vssd1 _0909_.A a_8701_25953# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4830 a_25842_23413# a_25674_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4831 vssd1 _1764_.A _1764_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4832 vssd1 _1261_.A1 a_8624_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4834 vssd1 _1030_.B a_12441_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4835 _1583_.X a_18607_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4836 a_5888_32143# a_5639_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4837 vccd1 a_26295_2986# _1801_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4838 a_8440_10499# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4839 vssd1 _1050_.B _1050_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4841 vssd1 _1070_.A2 a_18048_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X4844 _1109_.B a_16791_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4845 a_23627_6740# _1592_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4846 a_2686_23439# clkbuf_1_1__f__0380_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4847 vssd1 _1823_.CLK a_22199_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4848 a_24573_2773# a_24407_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4849 _1015_.A1 a_10167_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4850 a_23707_29967# a_23009_29973# a_23450_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4851 a_25309_29423# a_25143_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4852 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4853 vccd1 _1110_.A a_16863_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4855 a_25674_23439# a_25401_23445# a_25589_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4856 a_3410_2767# a_2971_2773# a_3325_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4857 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4858 vccd1 a_19487_21972# _1828_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4860 vssd1 a_2382_6005# a_2340_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4861 a_27057_28335# a_26891_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4863 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4864 a_2382_4917# a_2214_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4865 a_13632_8751# _1568_.B a_13057_8897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X4866 vssd1 a_25455_31965# a_25623_31867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4867 vccd1 a_24719_25615# a_24887_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4868 a_6968_21379# _1448_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4869 vssd1 a_23443_7338# _1676_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4870 _1494_.A a_17088_26819# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4872 a_17496_15055# _1887_.Q a_16921_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X4873 vssd1 a_4495_11989# _1217_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4875 _1197_.B a_10515_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4876 vssd1 a_25455_2589# a_25623_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4877 vssd1 a_27571_2589# a_27739_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4878 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4879 _1267_.A1 a_4739_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4880 a_7159_20884# _1557_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4881 vssd1 _1768_.A a_7295_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4882 a_21273_3133# a_21003_2767# a_21183_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4883 vssd1 a_23266_8863# a_23224_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4884 a_11877_29423# a_11711_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4885 vccd1 a_3801_28981# _0909_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4886 vssd1 a_24719_25615# a_24887_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4887 vssd1 _1278_.X a_4036_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4888 vssd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4890 vssd1 _1074_.C a_18673_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4891 a_19487_21972# _1395_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4892 a_14226_17027# _1405_.B a_14144_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4893 a_24577_15823# _1701_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4894 a_12073_14191# _1231_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4896 a_2340_28335# a_1941_28335# a_2214_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4897 a_19697_30511# a_19531_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4898 _0909_.A _1255_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4900 _1732_.X a_22195_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4901 a_14733_4943# _1749_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4902 a_19709_6575# a_19439_6941# a_19619_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4903 a_4571_7119# a_3707_7125# a_4314_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4905 _0992_.A2 a_12927_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4906 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4907 vccd1 a_22622_26677# a_22549_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X4909 _1091_.C1 a_16863_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4910 a_9823_25981# _1332_.Y a_9460_25847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4911 _1141_.C _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4912 vccd1 a_17113_6005# _0999_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4914 a_1673_20969# _1283_.B1 a_1757_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4916 vssd1 _1842_.Q a_18329_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4918 a_21407_2589# a_20543_2223# a_21150_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4919 a_12165_22895# _1901_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4920 a_23523_2589# a_22659_2223# a_23266_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4922 a_19053_20175# _1836_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4923 a_20755_32143# a_19973_32149# a_20671_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4924 vccd1 a_25455_21085# a_25623_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4925 vccd1 a_10643_6031# a_10811_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4926 a_6230_25321# _1243_.A a_6073_25045# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4927 vccd1 a_16311_18543# fanout37.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4928 a_7659_8029# a_7479_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4929 a_8569_2767# _1614_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X4930 vssd1 a_16911_1300# _1945_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4931 vccd1 _1982_.CLK a_25787_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4932 a_4237_17231# _1291_.A1 a_3799_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4933 a_9742_4511# a_9574_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X4934 a_20211_31055# a_19347_31061# a_19954_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4935 a_10103_21046# _1334_.A1 a_9644_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X4936 vccd1 a_27295_13469# a_27463_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4937 _1459_.A a_12815_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4938 a_9223_21263# a_9043_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4939 a_9844_30761# a_9595_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4940 vccd1 _1840_.Q a_12570_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4941 vssd1 _0925_.A2 a_4351_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4942 a_4161_16367# _1231_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4943 a_8818_11703# _1120_.X a_9032_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X4944 vccd1 a_15299_21807# _1021_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4945 a_22825_3311# a_22659_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4946 vssd1 a_20395_30877# a_20563_30779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4947 vssd1 a_22898_24095# a_22856_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4949 vssd1 _1286_.A1 _1793_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4950 a_13455_32143# a_13275_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4952 _1300_.A2 _1325_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4953 _1146_.B a_20471_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4954 vssd1 a_19107_3855# a_19275_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4955 _1999_.CLK a_6283_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4957 a_4155_5487# _1267_.A1 _1804_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X4958 _1243_.A _1242_.A1 a_5174_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4959 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4960 a_16934_26525# a_16661_26159# a_16849_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4961 vccd1 _0958_.B a_17967_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X4962 a_18114_31029# a_17946_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X4963 _1418_.A a_16904_22467# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X4964 a_11902_23478# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4966 vssd1 a_11685_9813# _1008_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4967 _1324_.A _1052_.B1 a_8031_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4968 vssd1 a_20839_32117# a_20797_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4970 a_9823_15279# _1764_.A a_9460_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4971 a_17221_11837# _1010_.A a_17139_11584# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4972 _1322_.A a_5547_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4975 a_13399_17483# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4976 a_10727_6031# a_9945_6037# a_10643_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4977 a_18272_17705# _1049_.B1 a_18170_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4978 a_25674_23439# a_25235_23445# a_25589_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4979 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z _1243_.Y a_8464_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4981 a_23523_22173# a_22659_21807# a_23266_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X4982 a_5727_17999# _1780_.B1 a_5509_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X4983 a_6610_13879# _1175_.B2 a_6824_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X4985 a_14641_16367# _1850_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4986 vssd1 a_18850_2741# a_18808_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X4988 a_19605_31599# a_19439_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4989 _1405_.B a_17047_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4990 vssd1 fanout20.X a_23855_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4991 a_17017_8573# _1146_.B a_16945_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4992 a_12771_21482# _1549_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4993 a_11789_2223# _1647_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X4994 a_11957_6575# _1117_.B a_11885_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4995 _1033_.A1 a_25623_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4996 vssd1 a_25623_6843# a_25581_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4998 a_27548_9839# a_27149_9839# a_27422_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4999 _1467_.A a_14467_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5000 a_2398_25437# a_1959_25071# a_2313_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5001 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5002 vssd1 _1762_.A _1762_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5003 a_2594_31055# clkbuf_0_net57.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5004 a_17578_29789# a_17139_29423# a_17493_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5005 a_6914_28879# _1243_.A a_6611_29111# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X5006 vssd1 _2004_.Q a_6927_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5007 vssd1 a_9460_15431# _1199_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5008 a_22454_2767# a_22015_2773# a_22369_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5009 a_2615_31921# _1329_.A0 a_2103_31573# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X5010 a_21445_26159# a_21279_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5011 vccd1 a_25198_24095# a_25125_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5012 a_26502_23261# a_26229_22895# a_26417_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5013 a_13165_13103# _1199_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5014 a_1816_11587# _1781_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5015 a_15750_28335# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5016 _1985_.CLK a_24039_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5017 a_23791_29967# a_23009_29973# a_23707_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5018 vssd1 _0909_.C a_3956_29239# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
X5019 a_18329_27247# a_18059_27613# a_18239_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X5021 a_23193_22173# a_22659_21807# a_23098_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5022 a_23925_4233# a_22935_3861# a_23799_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5023 a_7825_4233# a_6835_3861# a_7699_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5024 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5025 vssd1 a_1828_19061# _1260_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5026 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5027 a_6829_29199# _1337_.S a_6611_29111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5029 vccd1 _1252_.A a_5731_12567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5030 a_11793_12925# _1110_.A a_11711_12672# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5031 _1090_.X a_16219_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5032 _1736_.X a_21183_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5033 a_22346_5599# a_22178_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5035 vssd1 a_28015_12283# a_27973_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5036 vssd1 a_24462_25589# a_24420_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5038 vssd1 a_25271_2767# a_25439_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5039 a_9920_25223# _1305_.B a_10062_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5042 _1077_.D1 a_12447_17024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5043 _1187_.A a_18519_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5044 a_21721_31599# a_21555_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5045 vccd1 _1261_.A1 a_8706_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5046 vccd1 a_9613_22869# a_9643_23222# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5048 a_21051_4074# _1743_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5049 _1537_.B a_9871_10391# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5050 vssd1 a_1643_23413# io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5051 a_22346_5599# a_22178_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5052 _1845_.Q a_16699_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5054 a_14825_2767# _1934_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5055 a_27406_20831# a_27238_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5056 _1820_.Q a_17895_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5057 vccd1 a_5169_13149# a_5269_13367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X5060 vssd1 a_6797_19605# _1325_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5061 a_23558_8207# a_23119_8213# a_23473_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5062 _1852_.Q a_12467_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5063 a_25842_22325# a_25674_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5065 vssd1 a_13587_29967# a_13755_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5066 vccd1 _1862_.Q a_14776_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5067 a_17685_3311# a_17415_3677# a_17595_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X5068 vccd1 a_10570_19743# a_10497_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5069 _1089_.B a_21207_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5070 vssd1 _1764_.B _1769_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5071 vccd1 a_16439_3677# a_16607_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5072 a_10585_22729# a_9595_22357# a_10459_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5073 a_2723_3677# a_1941_3311# a_2639_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5074 a_3536_3145# a_3137_2773# a_3410_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5075 vssd1 _1764_.A a_10814_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5077 a_21091_24349# a_20911_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5078 _1327_.A1_N _0925_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5080 _1577_.X a_20676_12265# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5081 vccd1 _1346_.A a_7790_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5082 _0921_.Y _0921_.A a_23205_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5083 a_17727_27791# a_16863_27797# a_17470_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5084 a_24386_14735# a_23947_14741# a_24301_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5086 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5087 a_2195_12533# _1301_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X5088 a_26969_16367# _1387_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5089 _1849_.CLK a_15794_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5090 _1464_.B a_10167_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5091 a_25674_22351# a_25401_22357# a_25589_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5092 vssd1 a_26854_14303# a_26812_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5094 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5095 a_23443_12778# _1711_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5097 vccd1 _1886_.Q a_21091_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5098 vccd1 a_27590_5599# a_27517_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5099 a_26628_25071# a_26229_25071# a_26502_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5100 _1395_.A a_18100_19203# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5101 a_22238_13647# _1006_.B2 a_22081_13621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5102 vccd1 a_12873_14337# _1038_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X5103 vssd1 a_23523_4943# a_23691_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5104 _1464_.B a_10167_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5105 _1121_.A1 a_5199_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5106 a_17317_13103# _1403_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5107 a_3065_11177# _1226_.B1 _1219_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5108 vccd1 _1723_.A_N a_22015_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5109 _1068_.C1 a_14287_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5110 a_17673_32149# a_17507_32149# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5112 a_17397_27791# a_16863_27797# a_17302_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5113 vssd1 a_14979_17130# _1821_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5114 vccd1 a_4003_2741# a_3919_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5115 vssd1 _0997_.X a_17956_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X5117 _1907_.CLK a_8307_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5118 a_7006_26409# _1306_.A2 a_6703_26133# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X5121 vccd1 a_28015_10107# a_27931_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5122 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_9844_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5123 a_14733_3855# _1622_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5124 a_6467_9001# _1086_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X5125 vccd1 a_20230_28447# a_20157_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5126 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_16127_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5127 a_14226_27907# _1484_.B a_14144_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5128 a_11030_27359# a_10862_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5129 a_9258_10089# _1198_.A2 a_9176_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5130 vssd1 _1020_.X _1034_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5131 a_22063_22570# _1509_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5132 vccd1 _0992_.A2 a_11842_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X5133 a_22622_24501# a_22454_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5134 vccd1 a_16734_8863# a_16661_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5135 _1438_.X a_12259_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5136 _0939_.A a_16863_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5137 a_7803_20884# _1445_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5138 vccd1 _1999_.CLK a_11435_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5139 _1639_.X a_12815_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X5140 vssd1 a_3759_21237# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X5141 a_2472_19605# _1311_.A1 a_2692_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5142 a_10331_10927# _1198_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5143 a_20429_26159# a_19439_26159# a_20303_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5144 vccd1 _1883_.Q a_20298_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5145 vccd1 _1833_.Q a_18642_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5146 _1982_.CLK a_22050_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X5147 a_22729_6575# a_21739_6575# a_22603_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5148 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5150 vccd1 _1289_.A2 a_5829_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5151 a_11760_23671# _1305_.B a_11902_23478# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5152 vccd1 a_26651_4765# a_26819_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5153 _1334_.A1 _1301_.A1 a_6671_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5154 vssd1 _1049_.X _1050_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5155 a_19981_13647# _1191_.B1 a_20065_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5156 _1782_.A a_4627_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5157 vccd1 _1744_.A_N a_21279_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5158 a_17221_18543# _1826_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5159 a_12973_5461# _0993_.X a_13130_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5160 a_22454_24527# a_22181_24533# a_22369_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5161 _1445_.A a_9176_19881# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5162 _1525_.A a_22195_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5163 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5165 a_16245_9867# _0939_.A a_16159_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5166 a_2769_22057# _1762_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5167 _1217_.A3 _1207_.B1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5168 vccd1 a_22799_7338# _1920_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5169 _1836_.Q a_28015_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5170 vssd1 a_22247_20884# _1879_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5171 vssd1 a_25842_22325# a_25800_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5172 _1067_.B a_8143_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5173 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5639_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5174 a_13495_2767# a_12797_2773# a_13238_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5175 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5176 vccd1 a_27663_21085# a_27831_20987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5178 vccd1 a_9937_4917# _1011_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5179 vccd1 _1121_.A1 a_9233_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5180 vccd1 a_27314_2335# a_27241_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5181 a_15017_26159# _1896_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5183 _0923_.Y _1775_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5184 _1689_.A a_21091_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5185 vccd1 a_22546_6031# a_22652_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5186 a_22247_20884# _1502_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5187 a_22935_19087# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5188 a_23303_15823# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5189 a_21978_30623# a_21810_30877# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5190 vssd1 _1860_.CLK a_9595_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5191 a_26651_8029# a_25787_7663# a_26394_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5192 _1968_.Q a_27095_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5193 _1038_.C1 a_16495_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5195 vccd1 a_23266_21919# a_23193_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5196 a_25309_9839# a_25143_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5197 vccd1 a_12743_11445# a_12659_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5198 a_23101_3861# a_22935_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5199 _1308_.B _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5200 vssd1 a_27590_9951# a_27548_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5201 vssd1 _2006_.Q a_12079_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5203 _1140_.C a_7442_17429# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5204 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5205 vccd1 _1242_.A2 a_2309_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5206 a_9949_29423# _1903_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5207 a_5015_17231# _1249_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X5208 a_22580_3145# a_22181_2773# a_22454_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5209 a_23523_2589# a_22825_2223# a_23266_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5213 vccd1 a_13599_2388# _1938_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5214 _1084_.C1 a_1626_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X5215 a_11023_7338# _1649_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5216 a_10083_31055# a_9301_31061# a_9999_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5217 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5218 vccd1 _1838_.Q a_16986_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5219 _1041_.C1 a_12907_7232# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5220 a_4529_18319# _1267_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5222 _0966_.B1 a_16711_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X5223 vssd1 _1823_.CLK a_25235_16917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5224 vssd1 _1130_.C1 a_19405_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X5225 vccd1 _1390_.B a_19836_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5227 vssd1 a_20601_15797# _1082_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X5228 _1306_.A2 _1305_.B a_5639_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5229 a_4035_20693# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X5230 vssd1 a_3635_27765# a_3593_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5231 vssd1 a_11115_7828# _1614_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5232 a_6600_24233# _0911_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5233 vccd1 _1424_.A_N a_14287_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5234 a_14361_7125# a_14195_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5235 a_22181_31061# a_22015_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5236 vccd1 fanout28.A a_9779_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X5237 a_16113_2223# _1947_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5238 a_21235_7338# _1597_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5240 vssd1 a_16035_7119# _1590_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5241 a_14725_8527# _1149_.A1 a_14287_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5242 a_21905_30877# a_21371_30511# a_21810_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5243 a_8372_25077# _0909_.A a_8300_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5244 vccd1 _1860_.CLK a_13367_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5245 vccd1 _1226_.A1 a_4709_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5246 _1084_.A1 a_12723_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5247 _1308_.B _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5248 a_25581_15279# a_24591_15279# a_25455_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5249 a_9761_2223# a_9595_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5250 a_3210_24501# a_3042_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5251 vssd1 _1888_.Q a_19388_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5252 vccd1 a_23523_9117# a_23691_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5253 vssd1 _1816_.CLK a_2971_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5256 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5257 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_7925_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5258 vccd1 _1762_.A a_7201_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5259 a_13783_5162# _1609_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5260 a_23684_8585# a_23285_8213# a_23558_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5261 vssd1 _1324_.A a_6743_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5262 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5263 vccd1 a_22863_29691# a_22779_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5264 a_12532_27023# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5266 a_24945_17455# _1914_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5267 _1381_.A a_14144_17027# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5268 vccd1 _1639_.X a_15207_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5269 vccd1 a_14231_21263# a_14399_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5270 _1292_.C1 a_3799_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5272 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5273 a_26225_14025# a_25235_13653# a_26099_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5274 vccd1 a_11030_3423# a_10957_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5275 a_16565_21807# _1530_.B a_16219_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5276 a_13130_5737# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5277 a_5448_10933# a_5261_10973# a_5361_11191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X5278 a_22879_24527# a_22181_24533# a_22622_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5280 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5281 vccd1 _1084_.C1 a_6559_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5284 a_22454_24527# a_22015_24533# a_22369_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5285 a_9326_22895# _0913_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X5286 a_6559_12559# _1234_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5287 a_3956_29239# _0909_.B a_3884_29239# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5288 a_3042_24527# a_2769_24533# a_2957_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5289 vssd1 _1222_.A1 a_2331_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5291 vccd1 a_24979_14709# a_24895_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5292 a_5542_28111# _1242_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X5293 a_27053_22895# a_26063_22895# a_26927_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5295 a_2037_7663# _1789_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5298 _1686_.A a_23759_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5299 a_22549_2767# a_22015_2773# a_22454_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5300 vccd1 a_26267_16885# a_26183_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5301 a_16366_2335# a_16198_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5302 a_2143_29789# _1760_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5303 a_12226_16341# _0956_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5304 vccd1 _1192_.A2 a_9683_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5305 vssd1 _1050_.Y a_8480_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5306 a_25030_1501# a_24757_1135# a_24945_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5307 a_16661_9117# a_16127_8751# a_16566_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5308 vssd1 a_18107_21972# _1829_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5309 a_18560_18793# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5313 a_26870_17821# a_26597_17455# a_26785_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5314 a_21459_3677# a_21279_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5315 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_7479_28887# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5317 _0909_.B a_6600_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5318 vccd1 _1979_.Q a_27347_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5319 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5320 a_27330_11293# a_27057_10927# a_27245_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5321 a_15749_24527# _0966_.B1 a_15833_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5322 _0925_.A2 a_10423_21807# a_10951_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5324 vssd1 _1820_.Q a_14144_17027# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5325 a_6651_11587# _1124_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5326 vssd1 a_22707_18218# _1878_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5327 _1337_.A0 clkbuf_1_1__f_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5328 a_10041_24527# _0921_.B a_10399_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5329 _1104_.X a_15115_14851# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5330 a_22379_14557# a_22199_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5331 vccd1 a_21575_2491# a_21491_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5332 vccd1 a_23691_2491# a_23607_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5335 vssd1 a_25623_27515# a_25581_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5336 vccd1 _1459_.A a_18611_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X5337 a_23281_28169# a_22291_27797# a_23155_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5338 vccd1 a_16699_24251# a_16615_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5340 a_18497_1135# a_17507_1135# a_18371_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5341 a_17673_31061# a_17507_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5343 _0925_.A2 _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5344 a_2129_4399# _1783_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5345 a_1827_32117# _1337_.A1 a_2054_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X5347 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE _1353_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5348 a_5996_16367# _1265_.A1 a_5693_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5349 a_21150_2335# a_20982_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5350 a_18427_26525# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5351 a_8178_12015# _1082_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X5352 vssd1 _1790_.Y a_7381_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X5353 _1619_.X a_14328_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5354 vssd1 a_23818_23413# a_23776_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5355 vssd1 a_21327_20394# _1888_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5356 a_4247_19407# _1232_.Y _1257_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5358 a_27241_2589# a_26707_2223# a_27146_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5359 a_5087_29967# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5360 _1476_.B a_18171_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5363 _1318_.X a_5487_5281# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5364 vccd1 _1238_.X a_4351_22359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5367 a_6135_2589# a_5437_2223# a_5878_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5368 a_2148_10927# _1170_.B1 a_1657_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5369 a_20947_28879# a_20083_28885# a_20690_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5370 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5371 a_2122_8029# a_1683_7663# a_2037_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5373 a_5629_7913# _1168_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X5374 a_25949_8585# a_24959_8213# a_25823_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5375 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5376 a_17548_25321# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5377 a_17217_29967# _1477_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5378 a_21327_20394# _1521_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5380 vccd1 _1568_.B a_13488_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X5381 vssd1 a_12318_29535# a_12276_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5382 vssd1 _1860_.CLK a_9595_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5383 vssd1 a_22063_9514# _1578_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5384 vccd1 a_5693_19605# _1780_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5385 a_2198_9269# a_2030_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5387 vssd1 _2023_.CLK a_1775_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5388 _0903_.C a_5639_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X5390 vccd1 _1269_.A1 _1766_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5391 a_24945_8751# _1924_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5393 a_7742_6031# _1173_.X _1177_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X5394 a_21643_12381# a_21463_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5395 a_4715_7913# _1168_.X a_4497_7637# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5396 _1068_.D1 a_11711_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5398 _1817_.Q a_10627_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5399 a_3467_24527# a_2769_24533# a_3210_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5403 a_1828_14709# _1230_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X5404 vccd1 a_24639_23060# _1886_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5405 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5406 a_8767_9295# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5407 _1817_.Q a_10627_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5408 _1042_.B a_15411_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5409 a_10083_4765# a_9301_4399# a_9999_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5410 vccd1 _0930_.A _1175_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X5411 _1075_.X a_17691_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5412 _1709_.X a_22563_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5413 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5414 _1272_.B1 a_1779_22453# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X5415 vssd1 a_25991_8181# a_25949_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5417 vssd1 _1881_.Q a_20308_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5418 vssd1 a_17527_31867# a_17485_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5420 a_16074_5737# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5421 vssd1 _1261_.A2 a_7928_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5422 a_26099_26703# a_25401_26709# a_25842_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5423 a_8815_20214# _1233_.A1 a_8356_20407# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X5424 a_25539_15645# a_24757_15279# a_25455_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5425 vssd1 _0918_.A _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5426 vccd1 a_21978_30623# a_21905_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5427 vccd1 _1347_.Y a_7387_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5429 vccd1 _1304_.B a_1765_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5430 _1278_.A1 a_3063_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5431 a_17302_1679# a_17029_1685# a_17217_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5432 vccd1 a_13571_12533# a_13487_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5433 vccd1 _1876_.CLK a_26983_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5434 vssd1 _2005_.Q a_12691_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X5435 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X5436 a_18597_2767# _1938_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5438 a_16209_16617# _1829_.Q a_16127_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5439 a_16523_3677# a_15741_3311# a_16439_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5441 vssd1 a_4590_25183# a_4548_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5442 _1534_.A a_17548_25321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5443 a_15370_31055# a_14931_31061# a_15285_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5444 vssd1 _1875_.Q a_19480_25321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5445 a_13625_24533# a_13459_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5447 vccd1 _1744_.A_N a_17139_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5448 vccd1 _1140_.C a_14379_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X5449 vssd1 _1924_.CLK a_23119_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5450 a_6644_5263# _1202_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X5451 a_15725_7809# _1071_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5452 vssd1 a_23047_31029# a_23005_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5453 vccd1 _1261_.A1 a_7843_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X5454 vccd1 _1846_.Q a_9994_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5456 vssd1 _0983_.X a_12171_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5457 a_11793_5487# _0939_.A a_11711_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5458 a_20690_27765# a_20522_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5459 a_9828_26935# _1775_.A2 a_9970_26742# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5460 vccd1 _0923_.Y a_2009_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5461 a_7896_11079# _2008_.Q a_8038_11254# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5462 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5463 a_23297_30511# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5464 _1006_.B2 a_25623_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5465 _0974_.B1 a_20267_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5466 a_20522_28879# a_20249_28885# a_20437_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5467 a_10209_21629# _1903_.Q a_10137_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5468 a_9747_16367# _1764_.A a_9656_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X5469 a_20188_28335# a_19789_28335# a_20062_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5470 vssd1 _0958_.B a_15637_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5472 a_2644_11587# _1221_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5474 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5475 a_14629_18793# _1073_.X a_14557_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5476 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5477 a_14634_7119# a_14195_7125# a_14549_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5479 vssd1 a_7896_11079# _1162_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5480 vssd1 _1850_.CLK a_12539_12565# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5481 a_10876_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5482 _1760_.B temp1.inv2_2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5483 _1890_.Q a_27463_17723# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5484 _0921_.A a_2971_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5485 a_9253_14219# _1286_.A1 a_9167_14219# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5486 a_7472_13353# _1790_.Y _1791_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X5488 a_24903_19087# a_24039_19093# a_24646_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5489 _1191_.A1 a_27923_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5490 a_2616_27247# a_2217_27247# a_2490_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5491 vccd1 _1032_.C a_19103_13985# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5493 a_11902_23805# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X5494 a_22898_24095# a_22730_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5495 _1654_.X a_6739_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5496 a_7295_6351# _1171_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X5497 a_19439_7663# _1111_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5498 vssd1 a_15151_30877# a_15319_30779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5499 _1141_.C _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X5500 vssd1 a_25455_15645# a_25623_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5501 a_26225_24905# a_25235_24533# a_26099_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5502 vccd1 a_5136_22583# _1303_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5504 vccd1 a_22081_14709# _1190_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5505 a_10957_27613# a_10423_27247# a_10862_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5507 _1070_.A2 a_16711_15307# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5508 a_11476_20969# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5509 a_26283_18909# a_25585_18543# a_26026_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5510 vccd1 _1820_.Q a_14226_17027# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5511 vccd1 _1074_.C a_17723_20513# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5512 a_8497_12015# _1084_.B1 a_8178_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X5513 a_24573_19087# a_24039_19093# a_24478_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5514 _1028_.X a_18427_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5515 a_7939_13967# _1175_.B2 _1175_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X5516 vssd1 a_18151_19631# _1032_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5517 vssd1 a_6927_17999# _1764_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5518 _0958_.A a_13551_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5519 vccd1 _1217_.A2 a_4351_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5520 a_10543_22351# a_9761_22357# a_10459_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5521 a_15265_21237# _1074_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5522 a_25198_13215# a_25030_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5523 vssd1 a_23903_1300# _1991_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5524 a_10125_7497# a_9135_7125# a_9999_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5525 a_24110_11471# a_23671_11477# a_24025_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5526 vssd1 a_17727_27791# a_17895_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5527 vssd1 a_20701_14709# _0953_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X5528 vssd1 a_2623_1403# a_2581_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5529 a_13545_4399# a_13275_4765# a_13455_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X5530 vccd1 _1153_.A a_19439_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5532 vccd1 _0913_.A1 a_13019_20495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X5534 clkbuf_0_net57.A temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5535 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5537 vssd1 a_21327_13866# _1986_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5539 a_19567_1679# a_18703_1685# a_19310_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5540 a_5087_10496# _1234_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5541 a_11987_22895# _0984_.B1 a_12165_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5543 a_26091_10205# a_25309_9839# a_26007_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5544 a_2405_9839# a_2228_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5547 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5550 vssd1 _1091_.X a_15115_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5552 vccd1 a_20690_11445# a_20617_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5553 vssd1 a_26927_23261# a_27095_23163# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5554 a_17967_8751# _1719_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5555 vssd1 a_10349_25045# a_10283_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5556 a_23266_11039# a_23098_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5557 vccd1 a_1779_22453# _1272_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5558 a_21327_13866# _1725_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5559 a_7465_2223# _1952_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5561 vccd1 a_15163_4564# _1622_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5562 vssd1 a_1644_18517# _1300_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5563 a_2248_7663# a_1849_7663# a_2122_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5564 vccd1 a_10073_20693# a_10103_21046# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5566 vccd1 _1872_.Q a_18607_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5567 a_27149_3311# a_26983_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5568 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5569 vssd1 a_10643_29967# a_10811_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5570 vccd1 a_4847_1679# a_5015_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5571 vccd1 a_25198_1247# a_25125_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5573 a_25030_28701# a_24591_28335# a_24945_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5574 a_20947_27791# a_20083_27797# a_20690_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5575 vssd1 a_19310_1653# a_19268_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5576 a_21445_26159# a_21279_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5577 _2007_.D _1771_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5578 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5579 vssd1 _1764_.A _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5580 _1122_.A1 _1104_.X a_9779_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5581 vccd1 a_17470_29941# a_17397_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5582 a_16013_29423# a_15023_29423# a_15887_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5583 vssd1 a_10627_22325# a_10585_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5584 a_12337_10389# a_12171_10389# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5586 a_11953_11073# _1045_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5587 a_9687_12919# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X5589 _1117_.B a_10627_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5590 vssd1 _1062_.X a_17381_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X5591 vssd1 a_20591_7338# _1996_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5592 vccd1 a_10827_19997# a_10995_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5593 a_24853_9295# _1678_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5594 vssd1 a_18114_32117# a_18072_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5595 a_20897_2223# _1944_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5596 a_17319_6941# a_17139_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5597 a_15277_28111# _1841_.Q a_14931_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5599 vssd1 _1924_.CLK a_26983_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5600 a_23013_2223# _1636_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5601 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_13275_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5602 a_23189_20553# a_22199_20181# a_23063_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5603 _1650_.X a_4531_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5605 a_17293_11837# _1977_.Q a_17221_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5606 a_3145_14191# _1277_.A a_3063_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5607 a_26133_26159# a_25143_26159# a_26007_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5608 _1877_.Q a_25991_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5610 a_23098_9117# a_22825_8751# a_23013_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5611 fanout12.A _1287_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5612 vccd1 a_14287_29423# _1841_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5613 vccd1 _1010_.A a_10791_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5614 a_2953_20969# _1268_.X a_2869_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5615 vccd1 _1830_.CLK a_25235_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5617 vccd1 _1858_.Q a_13398_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5620 a_23650_16911# a_23211_16917# a_23565_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5622 a_2639_6031# a_1941_6037# a_2382_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5623 a_2309_3677# a_1775_3311# a_2214_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5625 a_18371_32143# a_17673_32149# a_18114_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5626 a_19567_14735# a_18869_14741# a_19310_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5627 a_22829_6031# a_22652_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X5628 vssd1 _1459_.A a_22015_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X5629 a_6607_6250# _1782_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5631 _1747_.A a_20539_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5633 _1749_.A a_17319_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5634 vccd1 a_21150_7775# a_21077_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5635 vccd1 _1329_.S a_2615_31921# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X5636 a_20004_26159# a_19605_26159# a_19878_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5637 a_5047_21237# _1292_.C1 a_5478_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X5638 _1756_.X a_6555_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5639 vssd1 a_23047_24501# a_23005_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5640 vccd1 _0930_.B a_4059_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X5641 a_4533_18793# _1326_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X5642 _1734_.X a_21459_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5643 _1065_.B a_25623_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5645 _1429_.A a_18239_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5646 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5647 _1898_.Q a_20471_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5648 a_27337_9839# _1926_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5649 _1099_.D1 a_17323_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5650 a_11865_12925# _1092_.B a_11793_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5651 a_17812_14441# _1033_.B1 a_17710_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5652 vccd1 _1150_.A2 a_17730_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X5653 vccd1 a_2455_9295# a_2623_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5654 a_2455_9295# a_1757_9301# a_2198_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5655 vccd1 a_5015_25339# a_4931_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5657 _1424_.A_N a_11711_15831# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5659 vccd1 _1760_.A_N a_7847_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X5660 _1242_.B1 a_7479_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5662 a_2686_23439# clkbuf_1_1__f__0380_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5664 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5665 _1764_.Y _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5666 _1022_.X a_17415_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5667 vccd1 _1876_.CLK a_22291_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5669 _1794_.Y _1304_.B a_9129_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5671 a_4351_12559# _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X5672 vccd1 a_24547_24746# _1880_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5673 _1050_.Y _1050_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5674 a_14760_7497# a_14361_7125# a_14634_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5675 _0965_.B1 a_17539_22923# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X5677 _1551_.A a_8440_24643# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5678 vccd1 a_4035_10901# _1246_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5680 a_20522_27791# a_20249_27797# a_20437_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5681 a_18751_5162# _1594_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5682 vccd1 a_23983_8207# a_24151_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5683 a_6921_5487# a_6651_5853# a_6831_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X5684 _1210_.B _1279_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5685 vccd1 a_23155_27791# a_23323_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5686 vccd1 _0913_.A1 a_4338_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X5687 vssd1 a_22339_19796# _1968_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5688 a_10287_2986# _1658_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5691 a_7479_8029# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5692 a_24547_24746# _1504_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5693 vccd1 a_24646_19061# a_24573_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5694 a_1791_13967# _1301_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X5695 a_2765_7497# a_1775_7125# a_2639_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5696 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5697 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5698 a_22898_27765# a_22730_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5699 a_22825_27247# a_22659_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5700 _1569_.A a_10511_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5701 _1560_.X a_9591_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5702 a_24719_25615# a_24021_25621# a_24462_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5703 a_10593_24233# _0921_.A a_10951_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5705 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X5706 a_13360_27023# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5708 a_14747_19200# _1864_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5711 vssd1 a_22771_6843# a_22729_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5713 vccd1 a_15319_16635# a_15235_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5715 vccd1 a_9000_14967# _1298_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5716 a_23266_3423# a_23098_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5718 _1154_.A1 a_23691_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5719 a_9769_6575# _0952_.A1 a_9687_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5720 a_22073_12533# _1151_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X5722 a_19664_23555# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5723 a_12502_4917# a_12334_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5724 a_11796_26159# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5725 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5726 a_17139_13103# _1070_.A2 a_17317_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5727 _1740_.X a_19619_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5728 _1677_.X a_21827_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5729 _1289_.B1 _0930_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5730 vccd1 a_21187_9295# _1685_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5731 vssd1 _1337_.S a_2326_32509# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X5732 vccd1 a_23351_25236# _1836_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5733 a_23443_9514# _1681_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5734 vccd1 a_7755_21263# _1762_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5735 a_25842_13621# a_25674_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5736 _1720_.A a_22195_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5737 a_1757_20969# _1282_.X a_1673_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5738 a_25125_1501# a_24591_1135# a_25030_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5739 a_23837_11477# a_23671_11477# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5740 vccd1 _1941_.CLK a_20543_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5741 a_12049_19631# _1819_.Q a_11977_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5742 a_5625_2223# _1356_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5743 vssd1 _1242_.A2 a_5345_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X5744 vccd1 _1038_.X a_14195_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5746 a_24110_10383# a_23671_10389# a_24025_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5747 vccd1 _1218_.B _1301_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5748 a_27149_19631# a_26983_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5749 vccd1 _1864_.Q a_14226_27907# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5750 vssd1 a_26295_18218# _1970_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5752 vssd1 a_27663_15645# a_27831_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5753 vssd1 _0930_.A a_7939_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
X5754 vssd1 _1903_.Q a_8025_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5755 a_12318_13621# a_12150_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5756 a_4931_1679# a_4149_1685# a_4847_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5758 fanout37.A a_16311_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X5759 vccd1 _1782_.A a_6375_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X5760 a_9963_15939# _2005_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5761 vssd1 a_2290_7775# a_2248_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5762 a_19521_12015# _1153_.A a_19439_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5763 vssd1 a_10627_29691# a_10585_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5765 a_24301_14735# _1979_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5766 vssd1 _1849_.CLK a_16127_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5768 a_10120_28585# a_9871_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5769 a_12557_16600# _2004_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X5770 a_16616_14441# _1099_.B1 a_16514_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X5771 a_27215_1300# _1652_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5772 _1021_.A a_15299_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X5773 vssd1 a_24554_14709# a_24512_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5775 _1557_.A a_8027_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X5776 a_26026_18655# a_25858_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5777 a_13705_16189# _1851_.Q a_13633_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5778 a_22015_3855# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5779 a_18601_16911# _1179_.C1 a_18519_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5780 _1793_.A2 _1314_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5781 a_7636_29673# a_7387_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5782 a_20407_2986# _1732_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5783 a_27789_20719# a_26799_20719# a_27663_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5784 vssd1 a_6835_18543# _1768_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5785 vssd1 a_26267_13621# a_26225_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5786 _1675_.X a_22563_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5787 vccd1 _1047_.C a_12447_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X5788 a_8112_18543# _1255_.A1 a_7809_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5789 vccd1 a_25455_6941# a_25623_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5790 _1330_.X a_4035_30485# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5792 a_19973_29789# a_19439_29423# a_19878_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5793 a_15640_27497# a_15391_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X5794 vccd1 a_20131_27412# _1843_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5795 a_15059_7119# a_14361_7125# a_14802_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5796 a_15538_32117# a_15370_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5798 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5799 a_25401_24533# a_25235_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5800 vssd1 a_18114_31029# a_18072_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5801 _2008_.Q a_3083_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5802 a_12502_4917# a_12334_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5804 vssd1 a_15265_21237# _1077_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X5805 vssd1 a_10811_8181# a_10769_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5806 vccd1 _1836_.Q a_19619_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5807 a_25582_29789# a_25143_29423# a_25497_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5808 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5809 vssd1 _0921_.B a_8399_23492# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5811 vccd1 temp1.capload\[15\].cap.A temp1.capload\[15\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5813 a_13579_2767# a_12797_2773# a_13495_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5814 a_17647_2388# _1637_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5815 vssd1 a_2807_28603# a_2765_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5816 a_23155_27791# a_22291_27797# a_22898_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5817 a_4404_18517# _1232_.Y a_4627_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5818 vssd1 _0925_.A2 a_3799_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5819 a_13265_11177# _1197_.D a_13183_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X5820 vssd1 a_9184_23047# _1341_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5821 a_7939_13967# _1766_.A0 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5822 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5824 _1876_.Q a_23323_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5825 vccd1 a_17470_1653# a_17397_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5826 a_8297_9001# _1813_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5827 a_15370_32143# a_15097_32149# a_15285_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5828 vssd1 a_9871_24527# _1308_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5831 vccd1 a_19735_14709# a_19651_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5832 vccd1 _1882_.CLK a_24591_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5833 a_2639_4943# a_1941_4949# a_2382_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5834 vssd1 _1205_.Y a_4101_8779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X5837 a_23707_29967# a_22843_29973# a_23450_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X5839 vssd1 a_24639_23060# _1886_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5840 _1422_.X a_12488_26409# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5843 vccd1 a_22162_31711# a_22089_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5844 a_19970_30877# a_19531_30511# a_19885_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5845 a_19513_31061# a_19347_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5846 a_23013_4943# _1929_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5848 a_13599_13866# _1755_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5849 a_23558_8207# a_23285_8213# a_23473_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5850 _1023_.B a_24703_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5851 _1873_.CLK a_22567_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5852 a_25823_22173# a_25125_21807# a_25566_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5853 a_9683_1501# a_9503_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5854 a_18751_21972# _1497_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5855 a_4789_20495# _1273_.A1 a_4443_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5856 a_6651_11587# _1086_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X5857 a_16849_31599# _1859_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5858 vccd1 a_1827_32117# _1338_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X5859 _1189_.B2 a_12743_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5860 a_27548_12015# a_27149_12015# a_27422_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5861 vccd1 a_27215_31274# _1465_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5862 a_15660_30287# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5863 a_6369_22895# _1242_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5864 a_22015_10383# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5865 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X5866 a_7711_5652# _1564_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5867 a_23377_29967# a_22843_29973# a_23282_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5868 _1037_.B a_20471_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5869 _0932_.A a_3247_12672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5870 vssd1 _1325_.B1 a_5167_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X5871 a_18697_17231# _1179_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5872 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8215_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X5873 a_18325_12015# _1153_.A a_18243_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5875 vccd1 _1053_.A a_16863_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5876 a_22181_26709# a_22015_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5877 a_5812_18319# _1786_.A1 a_5509_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5878 _1143_.X a_14655_18115# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5879 vccd1 a_12299_25437# a_12467_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5880 vccd1 a_11777_9269# _1192_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5881 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5884 a_23075_11690# _1680_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5885 vccd1 a_22695_29789# a_22863_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5887 a_4983_16143# _1277_.A _1289_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X5888 vssd1 a_18539_1403# a_18497_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5889 a_25965_32463# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5890 a_22369_31055# _1874_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5891 a_22365_20181# a_22199_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5894 vccd1 a_24830_15797# a_24757_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X5895 a_4262_30833# a_4213_30663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X5896 _1839_.Q a_23047_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5897 a_11023_18218# _1376_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5898 vssd1 _1873_.CLK a_22843_29973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5899 vssd1 a_8215_23983# _1474_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5900 _1097_.X a_13551_15936# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X5901 vssd1 _1313_.X a_8295_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X5902 a_3041_23983# a_2051_23983# a_2915_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5903 a_12488_4649# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5904 vssd1 a_18059_9839# _1153_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5905 a_7373_4399# _1816_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5907 vccd1 a_2472_19605# _1312_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X5908 vssd1 a_15538_32117# a_15496_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X5909 vccd1 a_9999_31055# a_10167_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5913 vccd1 _1199_.X _1250_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5915 a_22917_22357# a_22751_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5916 a_25125_17821# a_24591_17455# a_25030_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5917 vssd1 _1810_.A2 a_6548_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5918 _1074_.X a_16863_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5920 a_4587_24501# _1766_.A0 a_4796_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X5921 a_25842_16885# a_25674_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X5922 a_26781_16367# a_26615_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5923 a_4897_15823# _1249_.A2 _1289_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5924 a_2455_2589# a_1757_2223# a_2198_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5925 vccd1 a_2639_3855# a_2807_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5927 a_25030_21085# a_24591_20719# a_24945_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5928 vssd1 a_9999_31055# a_10167_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5930 _1219_.A2 _1226_.B1 a_3065_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5931 a_4814_24527# a_4765_24759# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X5932 a_15269_9661# _1057_.B a_15197_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5933 a_13813_24527# _1819_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X5935 a_9945_8213# a_9779_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5936 vssd1 _1841_.CLK a_17507_32149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5937 a_11704_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5938 vccd1 _0913_.A1 a_5455_20541# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X5939 vccd1 a_19735_1653# a_19651_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5940 a_2217_27247# a_2051_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5942 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_10120_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5943 a_23483_15823# a_23303_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5944 _1217_.A2 a_1775_12265# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5945 vccd1 a_25455_31965# a_25623_31867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5946 a_24803_25615# a_24021_25621# a_24719_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5947 a_15795_32143# a_15097_32149# a_15538_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5948 vccd1 a_23323_24251# a_23239_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5949 a_22879_1501# a_22181_1135# a_22622_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5950 a_9312_26159# _1344_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X5951 vssd1 _1873_.CLK a_21371_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5952 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5953 a_25674_16911# a_25401_16917# a_25589_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X5954 vccd1 a_9079_2767# a_9247_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5955 a_25842_12533# a_25674_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5956 a_25674_16911# a_25235_16917# a_25589_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5957 _1034_.Y _1020_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5961 vccd1 a_28135_12778# _1980_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5962 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_7636_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5963 vccd1 a_27295_24349# a_27463_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5964 a_9949_27791# _1818_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X5965 a_10129_29789# a_9595_29423# a_10034_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5966 vssd1 a_5231_22869# _1307_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5967 a_5303_9633# _1172_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5968 _1221_.B a_3095_9867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X5969 _1079_.B a_25899_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5971 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5972 vssd1 a_10423_21807# _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5973 vssd1 _1111_.B a_21549_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5974 vccd1 _1198_.A1 a_8395_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5975 _1149_.C1 a_11711_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X5979 vssd1 _1047_.C a_15545_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5980 a_8654_29967# a_8477_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5982 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_15640_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X5983 _1050_.Y _1049_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5984 a_6607_6250# _1782_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5985 vccd1 _1768_.A a_8031_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5986 a_16109_3677# a_15575_3311# a_16014_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X5987 a_4161_19087# _1254_.B1 _1257_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5988 a_17489_28885# a_17323_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5989 a_17444_19881# _1024_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X5990 _0965_.X a_18703_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5992 a_17075_9117# a_16293_8751# a_16991_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5994 a_12176_9839# _0991_.X a_11685_9813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5995 a_27973_3311# a_26983_3311# a_27847_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5997 vssd1 _1876_.CLK a_26983_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5998 a_14066_24501# a_13898_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X5999 a_27295_24349# a_26597_23983# a_27038_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6000 vccd1 _1768_.A a_9135_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6001 a_12659_13647# a_11877_13653# a_12575_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6002 _1667_.X a_18239_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6003 vccd1 a_12189_23737# a_12219_23478# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6004 vccd1 a_19395_5162# _1668_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6005 vccd1 a_24639_7828# _1982_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6006 vssd1 _1071_.B1 _1156_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6007 a_5152_31849# a_4903_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6008 a_9275_10602# _1560_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6009 a_3065_11177# _1226_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6010 vccd1 a_7101_14735# a_7201_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X6011 _1368_.X a_5588_6825# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6012 vssd1 a_22073_12533# _1154_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X6013 vccd1 a_6607_30186# _1555_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6014 a_20614_4765# a_20175_4399# a_20529_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6015 vccd1 a_23266_8863# a_23193_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
R7 temp1.capload\[9\].cap_54.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6016 a_11067_15529# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6017 a_25401_11293# a_24867_10927# a_25306_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6018 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_10506_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6019 a_17493_29423# _1475_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6020 a_24937_29257# a_23947_28885# a_24811_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6021 _1795_.X a_6324_13353# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6022 a_19057_1679# _1643_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6023 a_16083_14954# _1401_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6024 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6026 vccd1 _1177_.C a_3095_9867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X6029 a_25397_18377# a_24407_18005# a_25271_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6030 a_24294_1679# a_24021_1685# a_24209_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6032 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6033 a_10419_28879# a_10239_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6034 vccd1 _1053_.A a_15851_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6035 vccd1 a_7442_17429# _1140_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6036 _1147_.X a_17139_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6037 _1274_.A _1273_.A1 a_7566_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X6038 vssd1 _1442_.A a_9360_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6039 a_20131_6250# _1744_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6040 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5816_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6041 a_14461_20719# _1021_.A a_14379_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6042 vccd1 a_8785_20473# a_8815_20214# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6045 a_1641_13879# _1246_.A3 a_1887_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X6047 vccd1 a_9920_25223# _1349_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6049 vccd1 _1489_.A_N a_21647_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6050 a_14726_16733# a_14287_16367# a_14641_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6051 a_22983_21482# _1515_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6052 a_16665_25071# a_16488_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6053 a_17013_19777# _1021_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X6054 _1270_.A a_10423_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6055 vssd1 _0998_.B2 a_19709_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6056 a_5639_25615# _1242_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6057 a_9595_31965# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6058 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6059 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6060 vccd1 _1873_.CLK a_22015_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6061 a_2864_19881# _1311_.B1 a_2609_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X6062 vccd1 _1191_.A1 a_21218_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X6063 vccd1 a_14427_12778# _1573_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6064 a_12604_26703# a_12355_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6065 a_15005_26409# _1476_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6067 a_17998_9295# _1112_.D1 a_17749_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6068 a_10968_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6069 _1120_.X a_14287_13353# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6070 a_2723_28701# a_1941_28335# a_2639_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6071 vccd1 _1898_.Q a_14467_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6072 a_10464_1385# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6073 vssd1 a_7993_11989# _1086_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X6074 a_23699_22351# a_22917_22357# a_23615_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6075 a_9677_8751# _0935_.X a_9595_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6076 vssd1 a_27859_29098# _1855_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6077 _1904_.Q a_11455_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6078 a_19605_26159# a_19439_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6079 vccd1 _1768_.A a_8307_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6080 a_19388_21379# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6081 vssd1 _1849_.CLK a_18703_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6082 a_22369_24527# _1834_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6083 vssd1 a_25455_6941# a_25623_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6084 a_23627_6740# _1592_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6085 io_out[3] a_4863_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6086 _1657_.A a_7199_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6087 a_14427_12778# _1573_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6088 a_11777_9269# _1293_.A1 a_12030_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X6089 a_13070_2767# a_12631_2773# a_12985_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6090 vccd1 _1010_.A a_15943_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6091 a_13882_1653# a_13714_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6092 vccd1 _1047_.C a_16863_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6093 a_15151_10205# a_14453_9839# a_14894_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6094 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_12263_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6095 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6096 a_25953_4399# a_25787_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6097 a_13035_10383# a_12337_10389# a_12778_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6099 vccd1 a_25198_17567# a_25125_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6100 a_13040_23555# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6101 vssd1 a_10938_16341# _1075_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6102 a_22181_25621# a_22015_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6105 vccd1 a_18539_31029# a_18455_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R8 temp1.capload\[15\].cap_45.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6106 a_24278_11445# a_24110_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6107 a_6923_27791# a_6743_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6108 a_26229_25071# a_26063_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6109 vccd1 a_4035_23957# _1773_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X6110 _1762_.A a_7755_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6111 vssd1 a_23231_20149# a_23189_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6112 a_8807_17999# _1762_.A a_8449_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6113 vccd1 a_12927_13103# _1223_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X6114 a_27623_11471# a_27443_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6116 a_23565_23439# _1892_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6117 a_12171_8751# _1043_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6118 a_13656_31433# a_13257_31061# a_13530_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6119 a_4811_26703# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6120 a_15531_15444# _1398_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6121 vssd1 _1985_.CLK a_23947_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6122 _1281_.A1 a_2807_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6123 a_22181_1135# a_22015_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6124 a_22504_12559# _1190_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6125 a_24512_29257# a_24113_28885# a_24386_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6126 a_17262_19881# _1024_.D1 a_17013_19777# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6127 _1129_.B a_28015_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6128 _1071_.B1 _0987_.B a_10791_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6130 a_24945_13103# _1980_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6131 a_16911_31274# _1538_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6132 _1062_.X a_17967_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6134 a_15795_25615# a_15097_25621# a_15538_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6135 a_4248_27497# _1764_.Y a_3993_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6137 a_26007_10205# a_25309_9839# a_25750_9951# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6138 vssd1 a_15538_31029# a_15496_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6139 a_7479_17277# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X6140 vccd1 _1020_.A2 a_19973_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X6141 vssd1 _1128_.B a_19388_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6143 _1287_.A _1286_.A1 a_6646_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X6144 a_17060_26159# a_16661_26159# a_16934_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6145 a_7993_11989# _1084_.C1 a_8497_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6146 _0913_.Y _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X6147 a_18560_22467# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6148 a_2966_19131# _1762_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X6149 a_10218_1679# a_9945_1685# a_10133_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6150 vccd1 a_26203_10602# _1728_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6151 vssd1 _1086_.A a_6651_11587# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6152 vccd1 a_23351_7828# _1927_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6153 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6154 vssd1 _1344_.Y a_8215_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6155 a_22825_8751# a_22659_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6158 a_20709_7663# a_20543_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6159 vssd1 _1532_.A a_9871_10391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6160 _1107_.X a_13091_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6161 _1269_.B1 a_4351_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6162 vccd1 _1316_.A a_6870_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6163 a_22181_1685# a_22015_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6165 vssd1 _1841_.CLK a_17507_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6166 _1880_.Q a_26175_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6167 _2007_.Q a_5015_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6168 _1237_.B2 _1233_.X a_4985_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X6169 vssd1 _0918_.A a_10423_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6170 _1037_.B a_20471_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6171 a_12440_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6173 vccd1 a_7515_1501# a_7683_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6174 vccd1 _1242_.A2 a_6559_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X6175 a_20169_13103# _1878_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6179 a_2195_12533# _1246_.B2 a_2413_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X6180 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6181 a_22143_26525# a_21279_26159# a_21886_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6182 _1112_.B1 a_15391_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6183 a_23193_9117# a_22659_8751# a_23098_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6184 vssd1 _1841_.CLK a_17139_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6185 a_22622_31029# a_22454_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6186 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5152_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6187 a_14894_9951# a_14726_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6188 a_9442_18793# _1422_.B a_9360_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6189 vssd1 a_12815_9295# _1459_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6190 a_2005_32375# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X6191 a_27517_27613# a_26983_27247# a_27422_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6193 a_12355_32143# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6194 a_13616_30761# a_13367_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6195 temp1.capload\[1\].cap.Y temp1.capload\[1\].cap.A a_24677_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6196 a_25198_7093# a_25030_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6197 vccd1 a_25474_11039# a_25401_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6199 a_18059_25615# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6201 vccd1 a_5731_7127# _1448_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6202 a_19326_29967# a_19149_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6203 a_10191_27069# _1775_.A2 a_9828_26935# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6204 vccd1 _1261_.A1 a_8209_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X6205 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4075_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6206 a_2037_7663# _1789_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6208 _1485_.A a_19204_28995# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6209 a_27931_26525# a_27149_26159# a_27847_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6210 a_8929_2057# a_7939_1685# a_8803_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6211 _1665_.A a_15387_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6212 a_16120_28111# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6214 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6215 a_9919_25654# _1336_.A1 a_9460_25847# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6216 _1170_.A2 _1126_.Y a_27253_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6217 a_9301_7125# a_9135_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6218 _1766_.A0 _1269_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6219 a_20740_4399# a_20341_4399# a_20614_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6220 vssd1 a_17727_29967# a_17895_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6222 vccd1 a_10459_22351# a_10627_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6223 vccd1 a_2836_19319# _1233_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X6225 vssd1 a_24278_11445# a_24236_11849# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6227 a_13529_12937# a_12539_12565# a_13403_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6228 _1035_.X a_13367_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6229 vssd1 _1032_.C a_17293_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6230 vccd1 _1685_.A_N a_23579_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6231 a_3861_6397# _1281_.A1 a_3789_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6232 vssd1 _1242_.A2 a_2585_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X6233 a_8293_1679# _1565_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6235 vssd1 a_10459_22351# a_10627_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6236 a_8464_29673# a_8215_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X6237 _1769_.Y _1769_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6238 a_24639_4564# _1670_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6239 a_25589_13647# _1986_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6240 a_1849_7663# a_1683_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6241 a_23374_3855# a_23101_3861# a_23289_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6242 vssd1 a_26267_4917# a_26225_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6243 a_7274_3855# a_7001_3861# a_7189_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6244 a_23281_23983# a_22291_23983# a_23155_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6245 vssd1 _1069_.C a_12723_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X6247 a_20308_21379# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6248 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12604_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6251 a_17595_3677# a_17415_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6252 vccd1 fanout21.X a_22659_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
D1 vssd1 _1807_.Y sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X6254 vssd1 a_21235_25834# _1513_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6256 vccd1 _2009_.CLK a_1959_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6257 a_12535_1679# a_12355_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6258 a_12065_13647# _1906_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6260 a_25455_7119# a_24757_7125# a_25198_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6261 vccd1 a_23726_8181# a_23653_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6262 vssd1 _1127_.A a_10648_12675# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6263 vssd1 a_6559_9295# _0930_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6264 _1125_.X a_6651_11587# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X6265 vssd1 clkbuf_0_temp1.i_precharge_n.X a_1674_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6266 _1034_.Y _1029_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6268 vssd1 _2023_.CLK a_1683_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6269 vssd1 a_7755_21263# _1762_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6271 vssd1 _1015_.A1 a_10693_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6272 vssd1 _1139_.C a_11865_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6275 a_15197_14851# _1104_.D a_15115_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6276 vssd1 a_9186_13255# _1199_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6277 a_22825_27247# a_22659_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6278 a_27590_3423# a_27422_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6280 io_out[1] a_1643_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6281 a_14634_7119# a_14361_7125# a_14549_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6283 a_19487_2388# _1740_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6284 vssd1 a_1591_5487# fanout28.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6286 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6287 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6288 a_9949_2223# _1657_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6289 vssd1 _1231_.B1 a_2489_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6291 a_24945_28335# _1894_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6292 _1473_.A a_14144_27907# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6294 vccd1 _1231_.B1 a_3345_19131# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6297 _1767_.Y _1767_.B a_1683_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6298 a_22645_27791# _1876_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6300 vssd1 _1056_.X a_12723_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6301 _1899_.Q a_17895_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6302 vssd1 _1217_.B1 _1230_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X6303 vssd1 _1985_.CLK a_24591_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6304 vccd1 a_5871_1898# _1816_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6305 a_9489_5487# _2001_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6306 a_2602_31599# _1329_.A1 a_2103_31573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X6307 vccd1 fanout20.X a_22935_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6308 a_13196_3145# a_12797_2773# a_13070_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6309 a_2639_7119# a_1775_7125# a_2382_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6310 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6311 _1775_.C1 a_7387_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6312 vccd1 _1816_.CLK a_6835_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6313 a_24945_8751# _1924_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6315 a_17967_12672# _1965_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6317 vssd1 a_27279_14459# a_27237_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6318 a_3945_4917# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X6319 vssd1 a_18611_15823# _1506_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6320 a_25677_3677# a_25143_3311# a_25582_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6321 vssd1 a_10643_6031# a_10811_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6322 a_12384_11177# _0987_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6323 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6324 a_9963_15939# _0956_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6325 a_10045_15939# _0956_.C a_9963_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6327 a_10528_19631# a_10129_19631# a_10402_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6328 a_14410_4649# _1607_.B a_14328_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6330 a_11888_30287# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6331 a_22580_27081# a_22181_26709# a_22454_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6332 vccd1 a_18751_24148# _1834_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6333 a_21095_13103# _1079_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6334 a_5392_23983# _1287_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6335 vccd1 _1126_.Y a_4601_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
R9 temp1.capload\[1\].cap_46.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6336 a_10331_23145# _0983_.B1 a_10413_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6337 vssd1 a_23818_16885# a_23776_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6339 a_24025_10383# _1584_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6340 vssd1 a_6927_19087# _1269_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6341 a_27149_12015# a_26983_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6342 a_26670_23007# a_26502_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6343 a_9309_13647# _1012_.B _1012_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6345 a_19103_13985# _0958_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6346 _1448_.A a_5731_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6347 a_19142_17999# a_18703_18005# a_19057_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6348 _1155_.B a_14287_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6349 vccd1 _1153_.A a_11711_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6351 a_1975_29967# temp1.inv2_2.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X6352 vccd1 _1639_.X a_10147_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6353 vssd1 _1864_.Q a_14144_27907# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6354 _1436_.X a_10971_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6355 vccd1 _0961_.A a_17691_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6356 vccd1 _1128_.B a_19470_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X6357 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6358 vccd1 _1090_.C a_16219_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6359 fanout21.X a_23246_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6360 vssd1 _0918_.A a_10154_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6361 a_25639_3855# a_24775_3861# a_25382_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6362 a_21039_4765# a_20341_4399# a_20782_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6363 vccd1 _1723_.A_N a_22383_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6364 a_25313_8207# _1578_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6365 a_17723_20513# _0958_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6366 vssd1 a_17013_19777# _1024_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X6367 _1184_.A2 a_17723_20513# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6368 _1032_.C a_18151_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6369 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_15391_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6370 a_10459_22351# a_9595_22357# a_10202_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6371 a_4351_12559# _1217_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6372 vccd1 a_12226_16341# _0963_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X6376 a_23443_12778# _1711_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6377 a_13019_20495# _1781_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X6381 a_2009_21263# _1260_.B1 a_1643_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6383 vssd1 _0988_.X a_13264_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X6385 vccd1 _1304_.B a_5087_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6386 vssd1 a_21235_1898# _1992_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6387 _1521_.A a_20492_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6388 _1170_.B1 a_5496_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6389 a_20775_27412# _1492_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6390 a_22898_18655# a_22730_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6391 vccd1 a_14139_1679# a_14307_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6392 vccd1 _1873_.CLK a_21831_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6393 a_16986_22467# _1405_.B a_16904_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6395 vssd1 a_7387_15823# _1775_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6396 a_15115_14851# _1095_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6398 a_12797_2773# a_12631_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6399 a_21463_12381# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6400 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13616_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6401 a_16074_5737# _1047_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X6402 a_25401_4949# a_25235_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6403 a_2823_25437# a_2125_25071# a_2566_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6405 vssd1 a_5509_17973# _1786_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6406 vssd1 _1184_.B1 a_17496_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X6407 a_2214_3855# a_1775_3861# a_2129_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6408 a_5893_7663# _1168_.X a_5547_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6409 vccd1 a_13183_20719# _0964_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6410 vccd1 io_in[4] a_1626_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6411 a_19593_12015# _1135_.B a_19521_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6412 _1776_.X a_6968_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6413 vssd1 a_25382_3829# a_25340_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6414 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6415 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6416 a_8105_1685# a_7939_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6417 vccd1 a_3635_24501# a_3551_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6418 a_27931_19997# a_27149_19631# a_27847_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6419 a_11141_18543# _2005_.Q a_11041_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X6420 vccd1 a_18371_1501# a_18539_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6424 a_20907_6031# a_20727_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6425 vssd1 a_20655_28603# a_20613_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6426 vssd1 a_23075_11690# _1680_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6427 a_6736_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6428 a_8945_22717# a_8675_22351# a_8855_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X6429 a_2547_13469# a_1849_13103# a_2290_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6430 a_20131_6250# _1744_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6431 vssd1 a_12815_6031# _1639_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6432 a_10021_9985# _1071_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X6433 vssd1 _1047_.C a_13705_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6434 a_10270_10089# _1071_.B1 a_10021_9985# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6435 vssd1 _1095_.C1 a_14345_15425# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X6436 _1194_.A2 a_17895_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6437 a_13783_5162# _1609_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6438 vccd1 _0935_.X a_14103_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X6439 a_1941_4399# a_1775_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6440 a_18918_23555# _1405_.B a_18836_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6441 _1141_.C _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6442 a_22093_6575# _1582_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6444 vccd1 _1347_.Y a_8215_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6446 a_8654_2767# a_8215_2773# a_8569_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6447 vssd1 _1880_.CLK a_16863_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6449 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8464_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6451 _1362_.X a_10603_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6453 a_14369_5487# _0939_.A a_14287_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6454 vccd1 a_27923_11195# a_27839_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6455 vssd1 a_11759_29098# _1429_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6456 vccd1 _1999_.CLK a_9595_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6457 a_23653_8207# a_23119_8213# a_23558_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6459 vccd1 _1047_.C a_14471_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6461 vccd1 a_24462_1653# a_24389_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6462 a_14287_9001# _1193_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6463 a_13146_12533# a_12978_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6464 _1180_.X a_14931_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6465 a_16198_2589# a_15925_2223# a_16113_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6466 a_12202_11177# _1044_.X a_11953_11073# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6467 a_7969_17455# _1764_.A a_7885_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.08775 ps=0.92 w=0.65 l=0.15
X6470 vssd1 a_5503_4074# _0917_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6471 a_1941_4949# a_1775_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6472 a_4248_27497# _1764_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6474 vssd1 a_5455_17455# _1234_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6476 vssd1 a_13599_2388# _1938_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6477 a_27847_5853# a_27149_5487# a_27590_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6479 a_2869_20969# _1270_.A a_2787_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6480 _1604_.X a_20447_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6483 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6484 a_15054_26819# _1484_.B a_14972_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6486 a_24811_14735# a_24113_14741# a_24554_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6487 vccd1 _1021_.A a_14379_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6488 a_14894_16479# a_14726_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6489 a_18940_12533# _0974_.B1 a_19069_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6490 vssd1 _1015_.A1 a_10515_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6491 _1500_.A a_20999_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6492 a_10147_14735# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6494 vssd1 a_12743_1403# a_12701_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6496 vssd1 _0921_.B a_10765_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6497 _1972_.Q a_25623_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6498 _1232_.Y _0921_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6499 a_25559_10602# _1720_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6500 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6501 a_2405_23983# _1773_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6502 a_13533_21269# a_13367_21269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6503 a_25769_20175# a_25235_20181# a_25674_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6505 a_10471_7828# _1362_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6509 a_26479_1300# _1616_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6510 a_10073_20693# _1282_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6511 a_28135_13866# _1703_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6512 a_22063_11092# _1684_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6513 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6514 vssd1 a_22155_23658# _1691_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6515 a_26781_16367# a_26615_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6516 vccd1 _2003_.Q a_7755_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6517 a_20860_19203# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6519 a_18519_16911# _1179_.B1 a_18697_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6520 a_18237_4399# a_17967_4765# a_18147_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X6521 a_2631_8029# a_1849_7663# a_2547_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6523 vssd1 a_23155_24349# a_23323_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6524 _1272_.A2 a_2787_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6525 _1282_.A2 a_9284_21781# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6527 a_18397_12015# _1128_.B a_18325_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6528 a_9129_12879# _1316_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6529 vccd1 a_16055_29691# a_15971_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6530 vssd1 fanout33.A a_20083_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6532 a_25125_8213# a_24959_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6533 a_5354_28335# clkbuf_0_temp1.i_precharge_n.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6534 _1170_.A2 _1159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6535 a_25030_5853# a_24757_5487# a_24945_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6536 _1601_.A a_20308_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6537 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6538 vccd1 _1222_.B1 a_2195_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X6539 a_2217_27247# a_2051_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6540 a_6559_2767# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6541 a_5031_1501# a_4333_1135# a_4774_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6542 vccd1 a_22603_6941# a_22771_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6543 vssd1 a_20775_30186# _1871_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6544 vssd1 a_2287_16885# _1231_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X6545 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X6546 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13360_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6547 a_7756_17277# _2004_.Q a_7650_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X6548 a_2639_6031# a_1775_6037# a_2382_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6549 a_1864_18543# _1311_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6550 _1461_.A a_13316_25321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6551 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X6552 a_12705_12565# a_12539_12565# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6553 vccd1 a_15265_21237# _1077_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6554 vssd1 a_1641_13879# _1230_.A4 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6555 a_3247_12672# _0917_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6558 vccd1 a_10167_7093# a_10083_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
D2 vssd1 io_in[3] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X6559 _1404_.A a_19619_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6561 a_14410_3561# _1607_.B a_14328_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6562 vssd1 _1140_.C a_13337_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6563 a_14747_19631# _1869_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6566 vssd1 a_2639_3677# a_2807_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6567 vccd1 a_25991_22075# a_25907_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6568 a_18869_18005# a_18703_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6569 vssd1 a_25439_17973# a_25397_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6570 vssd1 _1764_.B a_4441_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6571 a_10951_24233# _0921_.A a_10593_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6572 vssd1 _1261_.A2 a_7111_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6573 vccd1 _1132_.A a_14747_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6574 a_9574_5853# a_9135_5487# a_9489_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6575 vccd1 a_10386_1653# a_10313_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6576 vssd1 a_13495_2767# a_13663_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6577 vccd1 _1020_.A2 a_18685_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X6578 a_27498_11039# a_27330_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6579 _1252_.A a_5361_11191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X6580 a_5174_30287# _1242_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X6582 vccd1 a_21051_22570# _1832_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6583 a_1945_6575# _1777_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6585 a_22319_30877# a_21537_30511# a_22235_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6586 a_27222_16479# a_27054_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6587 _1059_.B a_25623_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6588 a_10603_9117# a_10423_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6589 _1451_.X a_7567_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6590 a_11391_23060# _1422_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6591 _1045_.B1 a_11343_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6592 vssd1 _1767_.B _1767_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6594 a_7663_8207# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6597 _1870_.Q a_21115_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6598 vccd1 _2007_.Q _1053_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6599 vssd1 _1907_.CLK a_9779_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6600 vssd1 _1132_.X a_17565_24129# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X6601 vccd1 _1685_.A_N a_22383_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6603 a_11759_1898# _1662_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6604 _1391_.A a_22195_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6605 a_6997_10383# _1298_.A1 _1126_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6607 a_23903_26922# _1341_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6608 a_23266_21919# a_23098_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6609 a_27747_21085# a_26965_20719# a_27663_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6610 a_2030_9295# a_1591_9301# a_1945_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6611 vccd1 _1021_.A a_13551_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6612 _1064_.D1 a_14471_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6613 vccd1 a_25455_15645# a_25623_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6614 vssd1 a_7479_24527# _1242_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6615 vccd1 _1184_.A2 a_19053_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X6617 a_2340_4233# a_1941_3861# a_2214_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6618 a_1910_10927# _1170_.A2 a_1820_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X6620 a_17730_4943# _1150_.B2 a_17573_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6621 a_2897_10927# a_2696_11177# _1219_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6623 _1316_.A a_9167_14219# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6624 vssd1 _1243_.A _1243_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6625 vssd1 _1234_.A2 a_4237_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X6627 vssd1 a_15531_15444# _1399_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6628 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6629 a_14818_4943# a_14545_4949# a_14733_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6631 a_8480_21807# _1293_.A1 a_8177_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X6633 a_5061_23759# _1308_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6635 vssd1 a_22898_18655# a_22856_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6637 a_21909_31599# _1842_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6638 _1020_.B1 a_13919_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6640 vssd1 a_2455_1501# a_2623_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6641 a_24757_27247# a_24591_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6642 a_22730_24349# a_22457_23983# a_22645_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6643 a_8780_3145# a_8381_2773# a_8654_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6645 a_15633_11445# _1071_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X6646 vssd1 _0925_.A2 a_1855_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X6647 vccd1 a_14399_21237# a_14315_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6649 _1768_.A a_6835_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6651 vccd1 a_25363_9295# a_25531_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6652 a_25363_9295# a_24665_9301# a_25106_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6653 a_14655_23552# _1874_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6654 _1284_.B1 a_1591_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6655 a_25156_13103# a_24757_13103# a_25030_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6657 vssd1 a_17895_1653# a_17853_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6658 a_17996_24233# _0965_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6659 vccd1 a_27847_10205# a_28015_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6660 a_8807_17999# _1762_.A a_8449_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6661 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6662 _1406_.A a_18836_23555# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6666 vssd1 a_25474_11039# a_25432_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6667 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_12801_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X6668 a_24945_20719# _1699_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6669 a_14829_19453# _1132_.A a_14747_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6670 vssd1 a_27111_14557# a_27279_14459# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6672 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5980_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6674 vccd1 _1873_.CLK a_25235_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6676 a_2601_25935# _1763_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6677 vccd1 a_23542_3829# a_23469_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6678 _1809_.B a_6223_3339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X6680 a_21213_12897# _1153_.A a_21127_12897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6681 vccd1 a_7442_3829# a_7369_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6682 _1566_.X a_8579_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6683 a_19605_26159# a_19439_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6684 a_14726_10205# a_14453_9839# a_14641_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6685 a_15387_14557# a_15207_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6686 vssd1 _1141_.C a_17569_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6687 a_26785_13103# _1707_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
R10 temp1.capload\[2\].cap_47.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6690 a_11413_27247# a_10423_27247# a_11287_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6691 a_18685_16911# _1967_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6692 vssd1 _0981_.B a_14129_20513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6693 a_1941_3861# a_1775_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6694 vssd1 _1226_.A1 a_2897_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6695 _0984_.X a_12171_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6696 vccd1 a_5416_21781# _1785_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X6697 a_14533_20719# _1858_.Q a_14461_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6699 a_24205_10383# a_23671_10389# a_24110_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6700 a_9301_31061# a_9135_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6701 _1231_.B1 a_5455_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6702 _1152_.B a_26267_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6703 clkbuf_0_temp1.dcdel_capnode_notouch_.A temp1.dcdc.A a_15660_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6704 vssd1 _1830_.CLK a_18703_14741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6706 a_2505_16911# _1230_.B1 a_2287_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6707 _1057_.X a_15115_9408# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6708 a_13999_11471# _1156_.D _1156_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6709 vccd1 a_14802_7093# a_14729_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6710 a_12771_3476# _1623_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6711 a_3210_27765# a_3042_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6712 vccd1 _1896_.CLK a_19347_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6714 vssd1 a_27463_6843# a_27421_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6716 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9135_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6717 a_22181_1135# a_22015_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6718 vccd1 _1889_.Q a_22195_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6719 vssd1 _0951_.B a_17627_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6720 _1489_.A_N a_12815_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6721 a_21091_16911# a_20911_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6722 a_8749_2767# a_8215_2773# a_8654_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6723 vccd1 a_8325_10901# a_8355_11254# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6724 _1338_.A a_1827_32117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6725 vccd1 _1424_.A_N a_19439_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6726 _1826_.Q a_25071_19061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6727 _1074_.C a_9195_17973# a_8807_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6728 vccd1 a_2807_7093# a_2723_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6729 vssd1 _1781_.B a_5996_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6731 a_14839_10499# _1007_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X6733 _1839_.Q a_23047_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6734 a_9613_22869# _0913_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6736 a_22879_1679# a_22015_1685# a_22622_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6737 a_11711_6031# _0988_.X a_11889_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6738 _1045_.C1 a_12171_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6739 a_23005_31433# a_22015_31061# a_22879_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6740 a_28043_16042# _1705_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6741 a_7295_6351# _1173_.X a_7295_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6742 a_3042_27791# a_2769_27797# a_2957_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6745 vccd1 _1489_.A_N a_14747_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6746 vccd1 _1876_.CLK a_22015_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6747 a_12299_25437# a_11601_25071# a_12042_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6749 vssd1 a_22879_2767# a_23047_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6750 a_10313_1679# a_9779_1685# a_10218_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6751 a_14729_7119# a_14195_7125# a_14634_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6752 _1053_.A _2007_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6753 vccd1 _1967_.Q a_21091_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6754 a_10129_27791# a_9595_27797# a_10034_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6755 vccd1 _1887_.CLK a_22751_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X6756 vccd1 _1194_.A2 a_13130_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6757 a_15759_28879# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6758 vccd1 a_22073_12533# _1154_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X6759 a_7749_7663# a_7479_8029# a_7659_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X6762 _1696_.B a_26451_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6763 a_20529_4399# _1941_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6764 vccd1 a_22879_26703# a_23047_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6765 a_25198_17567# a_25030_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6766 _1326_.A2 _0930_.B a_3155_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6767 vssd1 a_13571_12533# a_13529_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6768 a_6981_12559# _1255_.A1 a_6559_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6769 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11704_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6770 a_27337_27247# _1836_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6771 _1889_.Q a_23691_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6772 a_6565_21041# _1282_.A2 a_6056_20871# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X6773 a_9079_2767# a_8381_2773# a_8822_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6774 a_25398_8207# a_24959_8213# a_25313_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6776 _1695_.A a_22103_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6778 a_12276_11849# a_11877_11477# a_12150_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6779 vssd1 a_22622_1653# a_22580_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6780 a_9700_5487# a_9301_5487# a_9574_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6781 vccd1 a_25807_3829# a_25723_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6782 vssd1 _1775_.A2 a_8372_25077# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X6783 vssd1 a_8177_12533# _1123_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6784 a_6713_24893# _1304_.B a_6641_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6786 a_9312_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X6787 vccd1 _1844_.Q a_15696_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6788 vccd1 _1823_.CLK a_26615_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6789 a_26597_13103# a_26431_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6790 vssd1 a_23266_27359# a_23224_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6791 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z _1243_.Y a_9312_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X6792 vccd1 _1837_.Q a_18423_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6793 a_25842_24501# a_25674_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6794 _1691_.A a_22195_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6795 a_15369_5321# a_14379_4949# a_15243_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6797 vssd1 _1876_.CLK a_23855_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6798 vssd1 a_18751_24148# _1834_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6799 a_9919_15606# _1199_.A1 a_9460_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6800 a_14287_17455# _1852_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6801 _1144_.X a_9687_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6802 a_20249_27797# a_20083_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6803 a_10511_9295# a_10331_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6804 a_2312_31599# a_2281_31751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X6805 a_24110_21263# a_23671_21269# a_24025_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6806 vssd1 _1459_.A a_18151_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6808 vccd1 a_9735_9514# _1759_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6809 vccd1 _1744_.B a_19803_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X6810 a_25455_31965# a_24757_31599# a_25198_31711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6811 a_17946_31055# a_17673_31061# a_17861_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6812 a_15800_26819# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6813 a_1737_14165# _1223_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X6814 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_6927_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6815 a_2048_15055# _1277_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6816 a_2156_9673# a_1757_9301# a_2030_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R11 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6818 a_24719_25615# a_23855_25621# a_24462_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6819 a_26417_22895# _1968_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6820 _1034_.Y _1034_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6821 vccd1 a_25198_5599# a_25125_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6822 vccd1 _1222_.A1 a_4798_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X6823 a_12759_4943# a_12061_4949# a_12502_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6824 _1875_.Q a_21115_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6825 a_24757_2223# a_24591_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6826 a_26873_2223# a_26707_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6827 vccd1 _1907_.CLK a_9135_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6828 a_24938_9295# a_24665_9301# a_24853_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6830 a_17270_6031# _0998_.B2 a_17113_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6832 vccd1 _1132_.A a_18519_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6833 a_4161_19087# _1254_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X6834 a_17456_7913# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6835 a_25842_6005# a_25674_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6836 a_10953_6575# _1562_.A a_10515_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6837 _0925_.A2 a_10423_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6838 vssd1 a_9742_7093# a_9700_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6839 a_20591_1898# _1629_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6840 a_24639_18708# _1695_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6841 a_2497_1679# _1651_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6842 vssd1 a_22603_6941# a_22771_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6845 a_24389_25615# a_23855_25621# a_24294_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6846 _1153_.X a_21279_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6848 a_15005_2767# a_14471_2773# a_14910_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6849 a_7553_8751# _1165_.C a_7469_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6851 a_12323_18365# _2004_.Q a_12232_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X6852 _1434_.X a_9912_13763# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X6853 a_24025_4399# a_23848_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6854 vccd1 a_23323_18811# a_23239_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6855 a_8031_17999# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6856 vssd1 _0989_.A2 a_3748_3971# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6857 a_6639_17455# _1261_.A1 _1267_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X6859 a_16175_9514# io_in[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6860 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_10506_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6861 vccd1 _1828_.Q a_17444_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6862 vssd1 a_3175_1653# a_3133_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6864 a_25589_4943# _1960_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6865 a_13714_1679# a_13275_1685# a_13629_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6866 a_14625_6575# _1063_.B a_14553_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6867 a_25198_8863# a_25030_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6868 vccd1 a_27663_15645# a_27831_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6869 a_25497_29423# _1880_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6870 a_12381_20747# _0961_.A a_12295_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6871 a_18949_7485# _1061_.B a_18877_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6876 vccd1 a_16366_2335# a_16293_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6877 vccd1 _1590_.A_N a_19439_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6878 _1355_.X a_5404_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X6879 vccd1 a_24278_10357# a_24205_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X6880 _1059_.B a_25623_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6881 a_2030_2589# a_1591_2223# a_1945_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6883 a_20359_6941# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6885 vccd1 _1873_.CLK a_21555_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6886 a_20395_30877# a_19697_30511# a_20138_30623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6887 a_7625_26677# _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X6888 a_1757_9301# a_1591_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6889 vccd1 _1218_.B a_1955_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X6893 vssd1 _1086_.B _1086_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6894 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.A a_14370_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6895 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5980_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X6896 a_19885_30511# _1871_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6897 vccd1 _1347_.Y a_9043_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6899 a_21051_24746# _1519_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6900 vssd1 _1723_.B a_22285_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6901 a_10459_2589# a_9761_2223# a_10202_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6902 a_25030_21085# a_24757_20719# a_24945_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6903 a_18887_19200# _1882_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6904 a_26394_4511# a_26226_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6905 vccd1 _1042_.B a_12570_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X6906 vccd1 _1311_.A2 a_2609_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6907 a_23523_27613# a_22659_27247# a_23266_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X6908 a_21143_21482# _1529_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6910 a_4404_18517# _1325_.X a_4533_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6911 a_3042_27791# a_2603_27797# a_2957_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6913 vccd1 a_7619_26324# _1818_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6914 a_27153_20719# _1823_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6915 a_26394_4511# a_26226_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6916 a_6743_10703# _1125_.X _1126_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X6917 a_27149_12015# a_26983_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6918 a_25858_18909# a_25585_18543# a_25773_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X6920 a_17946_31055# a_17507_31061# a_17861_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6921 a_11977_19631# _0958_.A a_11895_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6922 a_16495_12015# _1685_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6923 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4075_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6925 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6926 a_22015_21263# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6927 vssd1 fanout21.X a_24775_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6928 vssd1 a_26295_2986# _1801_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6929 a_13261_27791# a_13084_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6930 a_4521_1135# _1367_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X6931 vssd1 _0951_.B a_18637_11809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6932 vccd1 a_5271_20719# _1353_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6933 _1321_.C a_3707_6144# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6934 _1845_.Q a_16699_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6935 a_12318_29535# a_12150_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X6936 a_23193_27613# a_22659_27247# a_23098_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6938 a_4059_15431# _1323_.A2 a_4293_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X6939 a_2539_2589# a_1757_2223# a_2455_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6940 vssd1 a_11287_27613# a_11455_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6941 vccd1 a_23903_24746# _1881_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6942 a_22334_13967# _1974_.Q a_22244_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X6944 a_15285_31055# _1465_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6945 vccd1 a_15917_5461# _1196_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X6946 vssd1 _1110_.X a_17749_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X6947 vssd1 a_21051_22570# _1832_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6949 vssd1 a_27590_26271# a_27548_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X6951 _1226_.B1 _1208_.A1 a_7002_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6953 vssd1 _1277_.A _1323_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6954 vccd1 _1474_.A_N a_13275_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6956 vssd1 a_4404_18517# _1327_.A2_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6957 _1662_.X a_12535_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X6958 vccd1 a_2807_6005# a_2723_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6959 a_5693_16341# _1325_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X6962 a_2309_28701# a_1775_28335# a_2214_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6963 vccd1 _1823_.CLK a_24591_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6964 _1047_.C a_8454_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6965 a_18869_14741# a_18703_14741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6966 vccd1 _1876_.CLK a_22015_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6967 a_14287_14557# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6968 a_22063_11092# _1684_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6969 a_15594_21263# _1075_.X a_15514_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X6970 vccd1 a_2715_13371# a_2631_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6971 a_21150_7775# a_20982_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X6972 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6973 a_8449_17999# _1762_.A a_8807_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6975 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6976 a_25125_28701# a_24591_28335# a_25030_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6977 _2004_.D _1775_.C1 a_3993_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6978 a_9184_23047# _1305_.B a_9326_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6980 a_22931_15645# a_22751_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6982 a_25524_8585# a_25125_8213# a_25398_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6984 vccd1 a_11269_16600# a_10938_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X6985 a_25125_5853# a_24591_5487# a_25030_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X6986 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_3983_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X6987 vccd1 a_15963_32117# a_15879_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6988 io_out[7] a_27811_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6989 vssd1 a_4847_1679# a_5015_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6991 vccd1 _1768_.A a_4811_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6992 vssd1 _1198_.A1 a_8485_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6993 a_7563_23555# _0921_.B a_7481_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6994 vccd1 a_21575_23163# a_21491_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6996 a_12259_12381# a_12079_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X6997 vccd1 _1154_.A1 a_22504_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X6999 a_9779_11791# _1120_.X _1122_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26975 pd=1.48 as=0.08775 ps=0.92 w=0.65 l=0.15
X7000 vssd1 a_8307_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7001 a_2869_20969# _1269_.B1 a_2953_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7002 a_2309_1685# a_2143_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7003 a_14921_26409# _0965_.X a_14839_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7004 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7005 a_13077_29967# _1456_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7006 vssd1 a_23351_25236# _1836_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7007 vccd1 _0921_.A a_10593_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7009 vccd1 a_16863_9295# _0939_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7010 a_12500_15797# _1070_.X a_12892_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X7011 a_22648_12879# _1154_.A1 a_22073_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X7012 vccd1 a_15255_23060# _1899_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7013 vssd1 a_13974_21237# a_13932_21641# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7014 a_22285_16189# a_22015_15823# a_22195_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7015 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7016 vssd1 _0956_.C a_10667_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X7018 _1587_.X a_21136_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7019 a_18140_23983# _1843_.Q a_17565_24129# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X7021 a_9687_6575# _1144_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7022 a_4590_25183# a_4422_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7023 a_25842_23413# a_25674_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7024 a_20303_1501# a_19439_1135# a_20046_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7026 vssd1 fanout24.A a_24867_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7027 a_5670_6825# _1782_.A a_5588_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7028 a_20648_11849# a_20249_11477# a_20522_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7029 vssd1 a_3983_17455# _0921_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7030 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7031 vssd1 a_18371_1501# a_18539_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7034 _1577_.B a_12539_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7035 vssd1 a_4847_25437# a_5015_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7036 vssd1 a_24979_14709# a_24937_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7037 a_13009_13103# _1219_.A2 a_12927_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X7039 a_2823_25437# a_1959_25071# a_2566_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7040 vccd1 a_11023_5162# _1647_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7041 vssd1 _1880_.CLK a_25143_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7042 vccd1 a_21235_7338# _1924_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7043 a_2030_8207# a_1757_8213# a_1945_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7044 _0930_.B _0921_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7045 vccd1 _1314_.X a_7472_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X7047 a_19619_6941# a_19439_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7048 vccd1 _1156_.Y a_7656_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X7052 a_23443_9514# _1681_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7053 a_23741_22729# a_22751_22357# a_23615_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7054 a_14231_21263# a_13533_21269# a_13974_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7055 vccd1 a_27590_9951# a_27517_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7056 a_5721_10089# _1218_.B a_5639_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X7057 vssd1 a_3299_22325# _1240_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7058 vccd1 a_14986_4917# a_14913_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7059 a_11391_23060# _1422_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7060 a_27215_1300# _1652_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7061 vssd1 _1090_.C a_19593_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7062 a_27590_27359# a_27422_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7063 a_18239_25615# a_18059_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7064 a_16293_2589# a_15759_2223# a_16198_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7066 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_16120_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7067 a_19057_17999# _1821_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7068 a_10125_4399# a_9135_4399# a_9999_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7069 a_4160_32463# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7071 a_2493_25437# a_1959_25071# a_2398_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7072 vssd1 _1459_.A a_11711_16919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7073 vccd1 _1474_.A_N a_7387_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X7074 vssd1 a_19310_17973# a_19268_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7075 a_9227_17705# _1269_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7076 vccd1 _1063_.B a_14651_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7077 a_24677_30511# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7079 vssd1 _1896_.CLK a_19531_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7081 a_13840_2057# a_13441_1685# a_13714_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7082 a_20858_14735# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X7083 _1597_.A a_19619_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7085 a_27847_26525# a_26983_26159# a_27590_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7088 vssd1 a_20131_27412# _1843_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7089 a_25171_15823# a_24389_15829# a_25087_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7090 a_2932_18517# _1300_.A1 a_3152_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7091 vssd1 a_15725_7809# _1050_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X7092 _1769_.Y _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7093 vssd1 fanout20.X a_22659_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7095 a_17904_15823# _1070_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7096 a_18682_3855# a_18409_3861# a_18597_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7097 vssd1 _0935_.X a_14839_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7099 vccd1 _2007_.Q a_8307_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7100 _0997_.X a_15883_13131# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7101 vccd1 a_2290_13215# a_2217_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7102 _1628_.A a_15432_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X7103 vccd1 _2023_.CLK a_1591_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7104 a_22622_25589# a_22454_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7105 a_2156_2223# a_1757_2223# a_2030_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7106 a_15081_12533# _1100_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7107 _1843_.Q a_23875_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7108 _1841_.CLK a_14287_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7110 a_15575_19881# _0966_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7111 _1110_.X a_18519_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7112 vccd1 a_12587_14954# _1850_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7113 a_25582_10205# a_25143_9839# a_25497_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7114 a_12441_4221# a_12171_3855# a_12351_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7115 a_19112_9411# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7116 a_5478_21583# _1328_.S a_5183_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X7117 vssd1 a_23983_8207# a_24151_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7119 _1031_.X a_14747_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7120 a_12701_14025# a_11711_13653# a_12575_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7121 a_10862_3677# a_10423_3311# a_10777_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7122 _0992_.A2 a_12927_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7123 vccd1 _1110_.A a_18059_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7124 vccd1 _1070_.A2 a_17221_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7125 vssd1 a_17527_26427# a_17485_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7126 a_11789_2223# _1647_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7127 a_20601_15797# _1081_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7128 _1582_.A a_18560_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7129 vssd1 clkbuf_0_temp1.i_precharge_n.X a_1674_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7132 _1864_.Q a_20471_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7133 vccd1 _1165_.A _1171_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7134 a_20959_26922# _1553_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7135 a_23607_11293# a_22825_10927# a_23523_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7137 a_12587_14954# _1441_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7138 vccd1 a_23266_27359# a_23193_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7140 a_2539_9295# a_1757_9301# a_2455_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7141 a_13882_1653# a_13714_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7142 a_21051_4074# _1743_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7143 a_10648_12675# _0987_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7144 a_2769_27797# a_2603_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7145 vssd1 _1139_.C a_10817_17483# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7146 vccd1 a_13203_10357# a_13119_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7148 vccd1 _1011_.A1 a_10452_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7150 a_25497_26159# _1881_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7152 a_5449_22895# _1270_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7153 vccd1 a_1643_21237# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7155 a_7711_5652# _1564_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7156 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7157 a_25030_31965# a_24757_31599# a_24945_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7159 a_7458_4765# a_7185_4399# a_7373_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7160 a_9574_4765# a_9301_4399# a_9489_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7162 a_1941_28335# a_1775_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7163 a_17773_22717# _1021_.A a_17691_22464# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7164 vccd1 _1274_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7167 a_19439_3677# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7168 a_7803_6740# _1752_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7169 vccd1 _0909_.A a_8615_25953# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7171 vccd1 a_25198_28447# a_25125_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7173 a_24067_8207# a_23285_8213# a_23983_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7174 vssd1 _1141_.C a_18397_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7175 vssd1 a_6927_19087# _1269_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7177 vssd1 a_27498_28447# a_27456_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7178 vssd1 _1448_.A a_7387_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7179 vccd1 _1110_.A a_17967_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7181 vccd1 _1103_.A1 a_20539_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7182 _1506_.B a_18611_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7185 vssd1 a_27215_31274# _1465_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7186 vccd1 _1072_.X a_14629_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7187 a_2455_6941# a_1757_6575# a_2198_6687# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7188 vccd1 _1572_.B a_12384_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7189 vssd1 _0952_.A1 a_17139_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X7190 a_22402_12559# _1154_.C1 a_22322_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X7191 a_27422_26525# a_27149_26159# a_27337_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7193 vccd1 _0939_.A a_21095_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7194 a_5177_14441# _1217_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X7195 a_25397_3145# a_24407_2773# a_25271_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7196 a_20046_29535# a_19878_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7197 vssd1 a_19395_5162# _1668_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7199 a_24945_23983# _1972_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7200 a_9584_16367# a_9135_16367# a_9282_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7201 a_11647_31965# a_10865_31599# a_11563_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7202 a_14066_24501# a_13898_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7203 vccd1 a_7718_2335# a_7645_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7204 a_14139_1679# a_13441_1685# a_13882_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7206 a_5437_2223# a_5271_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7207 vccd1 a_13955_31055# a_14123_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7208 vssd1 _1108_.A1 a_11752_13353# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7209 a_12065_1135# _1612_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7210 _1246_.B1 _1301_.A1 a_2505_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7212 vssd1 _1870_.Q a_19204_28995# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7213 vssd1 a_25842_26677# a_25800_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7214 vssd1 a_23875_29941# a_23833_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7215 a_2861_17999# _1280_.Y a_2777_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7217 a_15462_29789# a_15189_29423# a_15377_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7218 _1860_.CLK a_9779_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7219 vccd1 _1887_.CLK a_25419_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7220 vccd1 a_21695_17620# _1826_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7223 a_14913_4943# a_14379_4949# a_14818_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7224 vssd1 a_26651_8029# a_26819_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7225 a_16175_1898# _1665_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7226 a_16156_7913# _0993_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7227 a_10021_9985# _1011_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7228 vssd1 a_13955_31055# a_14123_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7229 a_18519_20719# _1837_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7231 vssd1 _1270_.A a_1591_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7232 a_25198_1247# a_25030_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7233 vssd1 a_24811_28879# a_24979_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7234 a_2009_21263# _1308_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7235 a_24757_27247# a_24591_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7236 vssd1 fanout33.A a_14931_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7237 a_2765_4399# a_1775_4399# a_2639_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7238 _0963_.B a_12226_16341# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7239 a_25030_7119# a_24591_7125# a_24945_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7242 vssd1 _1816_.CLK a_5271_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7243 a_17746_29535# a_17578_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7244 vssd1 _1132_.C a_16797_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7245 a_22369_1679# _1940_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7246 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7248 _1141_.C _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7249 a_5692_15253# _0930_.B a_5912_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7250 a_17352_14735# _1184_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7251 a_4466_8527# _1170_.B2 a_4167_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X7252 a_1643_21237# _1260_.B1 a_2009_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.585 ps=2.17 w=1 l=0.15
X7253 a_1941_3311# a_1775_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7254 vssd1 _1198_.A2 a_9779_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26975 ps=1.48 w=0.65 l=0.15
X7255 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12532_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7256 vssd1 _1300_.B1 a_2932_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7257 a_11759_7338# _1657_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7258 a_4253_10927# _1226_.B1 a_4035_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X7259 _1640_.X a_17595_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7260 vccd1 fanout24.A a_24867_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7261 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_16127_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7262 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7263 vccd1 a_2566_25183# a_2493_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7264 a_5534_23145# _1303_.X a_5231_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7265 a_25674_26703# a_25235_26709# a_25589_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7266 a_19233_4233# a_18243_3861# a_19107_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7267 _1479_.A a_14743_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7269 a_2225_17705# _1250_.B2 a_2143_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7270 a_7657_7439# _1162_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7272 a_17217_17999# _1820_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7273 a_23565_16911# _1831_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7274 _1744_.A_N a_18151_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7275 _1364_.X a_8855_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7277 vssd1 a_22403_30779# a_22361_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7278 a_23649_5321# a_22659_4949# a_23523_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7280 _1885_.Q a_27463_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7281 a_15457_6005# _0952_.A1 a_15710_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7282 vssd1 _1887_.CLK a_22659_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7283 a_27847_19997# a_26983_19631# a_27590_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7285 a_10459_22351# a_9761_22357# a_10202_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7286 a_18059_6941# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7287 vssd1 a_28135_12778# _1980_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7288 a_14726_30877# a_14453_30511# a_14641_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7289 a_10073_20693# _1282_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7290 _1830_.Q a_19735_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7292 a_20947_27791# a_20249_27797# a_20690_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7294 a_10034_22351# a_9595_22357# a_9949_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7295 a_5817_5487# a_5625_5792# _1798_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X7296 vccd1 _1924_.CLK a_24591_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7297 a_11287_3677# a_10423_3311# a_11030_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7298 vccd1 _1867_.Q a_14743_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7300 vccd1 _0998_.A2 a_17270_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7301 vssd1 a_24639_7828# _1982_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7302 a_25800_12937# a_25401_12565# a_25674_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7303 vccd1 _1261_.A1 _1789_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7304 temp1.capload\[6\].cap.Y temp1.capload\[6\].cap_51.LO a_25965_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7305 vssd1 a_11563_31965# a_11731_31867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7306 vccd1 a_4127_22869# _1285_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7307 vccd1 _1322_.A a_5271_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7308 a_9489_7119# _1812_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7309 _1573_.A a_14467_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7310 a_27755_28701# a_26891_28335# a_27498_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7311 _1145_.B2 a_10811_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7312 a_8289_13103# _1034_.Y _1324_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X7313 a_4248_27497# _1242_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7314 vccd1 a_24703_11445# a_24619_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7315 a_25014_17973# a_24846_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7316 vssd1 a_2198_2335# a_2156_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7317 vccd1 _1267_.A1 _1801_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7319 vssd1 a_28015_27515# a_27973_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7320 vssd1 a_16531_24349# a_16699_24251# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7321 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7322 vccd1 a_17727_17999# a_17895_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7323 vccd1 a_8803_1679# a_8971_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7325 vssd1 _1255_.A1 _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7327 a_25708_9839# a_25309_9839# a_25582_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7330 a_8392_29199# _1347_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7331 a_12532_27247# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7332 a_16301_17455# _0964_.A a_16219_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7333 vccd1 a_2198_8181# a_2125_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7334 a_20999_17999# a_20819_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7335 vssd1 _1269_.A1 _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7336 a_2472_15431# _1219_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X7337 a_10988_3311# a_10589_3311# a_10862_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7338 a_27215_4074# _1366_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7339 vccd1 _1719_.B a_22195_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7342 a_4443_20175# _1302_.B1 a_4525_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7344 vccd1 temp1.capload\[3\].cap_48.LO temp1.capload\[3\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7345 _1039_.B a_12467_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7346 a_9742_7093# a_9574_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7347 a_11040_32143# a_10791_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7348 a_16661_31599# a_16495_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7349 a_20157_13353# _1007_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7350 vssd1 a_22622_1247# a_22580_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7351 a_13806_21263# a_13533_21269# a_13721_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7352 vccd1 _2006_.Q a_12027_20495# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X7353 _0998_.A2 a_21575_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7354 _1195_.A2 a_23691_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7355 a_14345_24129# _1056_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X7356 vccd1 _1763_.A2 a_2983_23217# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X7357 vssd1 _1311_.A1 a_3155_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7359 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7360 _1147_.C1 a_16863_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7361 a_11759_32362# _1467_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7362 vssd1 _1764_.B _1762_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7363 vccd1 _1768_.A a_10147_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7364 vccd1 a_20131_30186# _1869_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7365 a_8440_24643# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7366 a_25581_2223# a_24591_2223# a_25455_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7368 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7369 a_26409_18543# a_25419_18543# a_26283_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7371 _1205_.A1 a_3063_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7372 io_out[7] a_27811_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7373 a_2153_25615# _1762_.Y a_2408_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7374 vccd1 a_27222_16479# a_27149_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7375 a_5361_11191# _0916_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X7376 a_22181_31061# a_22015_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7378 a_4985_19881# _1234_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7379 a_11834_13353# _1537_.B a_11752_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7380 a_1857_10749# _1208_.A1 a_1775_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7381 a_2962_29967# clkbuf_0_temp1.i_precharge_n.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X7382 vssd1 _1860_.CLK a_13367_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7383 a_1644_18517# _1231_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X7384 a_11711_5487# _1067_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7385 vssd1 fanout24.A a_26891_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7386 vssd1 a_20414_32117# a_20372_32521# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7387 a_7645_2589# a_7111_2223# a_7550_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7388 a_26870_6941# a_26597_6575# a_26785_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7390 vssd1 _1887_.Q a_20492_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7391 vssd1 _1823_.CLK a_26615_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7392 a_1769_15823# _1231_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X7393 a_14335_25834# _1431_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7394 a_9360_3971# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7395 _0909_.A _0903_.C a_6981_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7396 vssd1 _0983_.A2 a_10493_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7397 a_10129_19631# a_9963_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7398 a_27422_19997# a_27149_19631# a_27337_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7399 a_9489_31055# _1860_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7401 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7402 vssd1 a_14427_12778# _1573_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7403 a_18453_25099# _0958_.A a_18367_25099# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7405 _1700_.X a_28083_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7406 a_17102_31711# a_16934_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7408 a_24025_21263# _1691_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7410 _1471_.A a_14144_26819# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7411 vccd1 a_9275_24746# _1900_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7413 _1769_.Y _1273_.A1 a_4441_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7414 a_16127_16617# _1070_.A2 a_16209_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7415 _1044_.X a_11159_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7416 a_17470_1653# a_17302_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7417 a_14427_12778# _1573_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7418 a_20671_32143# a_19973_32149# a_20414_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7419 a_20263_3855# a_20083_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7420 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_9871_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7422 a_4351_12559# _1217_.B1 _1277_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X7423 vccd1 _0929_.A a_3247_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7424 a_25030_24349# a_24591_23983# a_24945_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7427 a_22799_7338# _1587_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7428 vccd1 a_9963_20175# _1232_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7429 vccd1 _0964_.A a_14747_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7430 a_16863_12559# _1070_.A2 a_17041_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X7431 vccd1 _1286_.A1 a_6565_21041# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7433 a_27422_5853# a_26983_5487# a_27337_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7434 vccd1 _1760_.A_N a_2143_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7435 a_2471_22869# _1286_.A1 a_2698_23217# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X7436 vssd1 a_2623_9269# _0911_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7438 vccd1 _1744_.A_N a_21003_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X7439 vssd1 _0909_.A a_6713_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7440 vssd1 a_23351_7828# _1927_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7441 vssd1 _1140_.X a_12321_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X7443 vssd1 a_6245_14165# _1810_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7444 vccd1 a_20471_1403# a_20387_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7445 a_6901_11587# _1124_.X a_6829_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7446 vssd1 a_21143_21482# _1892_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7447 a_4443_20175# _1302_.B1 a_4525_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7448 vssd1 _1113_.C a_17845_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7450 vssd1 _1109_.B a_13545_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7451 a_25156_7497# a_24757_7125# a_25030_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7452 vssd1 _1267_.A1 a_4116_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7453 a_17812_7119# _0997_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7454 _1054_.C a_12061_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7455 _1154_.C1 a_19439_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7456 vccd1 a_20563_30779# a_20479_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R12 vssd1 temp1.capload\[4\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7457 vssd1 clkbuf_1_1__f__0380_.A a_1766_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7458 a_13551_15936# _1851_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7459 vccd1 _1766_.A0 a_7025_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7460 a_7050_21379# _1448_.A a_6968_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7461 vccd1 _0929_.A a_3983_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7462 vssd1 _1171_.Y a_7828_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7463 a_16911_31274# _1538_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7464 a_2405_23983# _1773_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7465 a_19973_31965# a_19439_31599# a_19878_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7466 _1481_.A a_14604_27497# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7467 vssd1 a_12973_5461# _1196_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X7469 a_15151_30877# a_14453_30511# a_14894_30623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7470 vccd1 _1762_.A a_5639_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7471 vccd1 a_26927_23261# a_27095_23163# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7472 a_25455_15645# a_24757_15279# a_25198_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7473 _1243_.A _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7475 vccd1 _1850_.CLK a_11711_13653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7476 a_18497_32521# a_17507_32149# a_18371_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7478 vssd1 a_15255_23060# _1899_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7479 _1202_.Y _1170_.A2 a_27713_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7480 a_14821_16733# a_14287_16367# a_14726_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7481 vccd1 a_18383_3476# _1941_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7483 a_6230_25321# _1306_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X7484 a_26099_13647# a_25401_13653# a_25842_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7485 a_8378_1679# a_8105_1685# a_8293_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7486 a_24757_6575# a_24591_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7487 vssd1 _1054_.C a_16005_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7489 _1198_.A1 a_6303_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7492 a_2125_8207# a_1591_8213# a_2030_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7493 vccd1 clkbuf_0_temp1.i_precharge_n.X a_5354_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7494 vccd1 _1907_.CLK a_14379_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7496 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13452_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7498 a_24945_1135# _1668_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7499 a_15943_10496# _1102_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7500 vssd1 a_18171_29691# a_18129_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7503 a_27747_15645# a_26965_15279# a_27663_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7505 a_1781_18793# _1311_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7507 a_6056_20871# a_6186_21041# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X7508 vccd1 _1047_.C a_13551_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7509 a_14776_15529# _0983_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7511 vccd1 a_18850_3829# a_18777_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7513 a_2601_25935# _0913_.A1 _2003_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7515 _1049_.B1 a_20267_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7516 a_8449_17999# _1762_.A a_8807_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7517 a_23266_8863# a_23098_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7518 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_11040_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7519 a_2408_25615# _1763_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7520 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X7521 a_2382_4511# a_2214_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7522 _1769_.B1 _1764_.B a_4811_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7524 a_24757_7125# a_24591_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7525 vssd1 a_25750_9951# a_25708_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7526 a_12570_22351# _1142_.D1 a_12321_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7527 vccd1 _1132_.A a_14839_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7529 a_7008_16367# _1789_.A1 a_6705_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7530 a_7002_4943# a_6644_5263# _1226_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7531 a_23155_27791# a_22457_27797# a_22898_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7532 vssd1 a_4003_2741# a_3961_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7533 a_5448_27247# _1344_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7535 a_24788_16201# a_24389_15829# a_24662_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7536 a_22730_18909# a_22457_18543# a_22645_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7537 vccd1 a_27295_6941# a_27463_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7540 a_25743_1898# _1654_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7541 a_2769_24533# a_2603_24533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7542 vccd1 _1880_.Q a_19746_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X7543 vccd1 _1132_.C a_13919_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7545 a_13361_11177# _1191_.X a_13265_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X7546 a_14129_20513# _1053_.A a_14043_20513# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7547 vccd1 a_15299_18543# _0961_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7548 vccd1 _0951_.B a_15943_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7549 a_25842_6005# a_25674_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7550 vccd1 _1234_.A1 a_6559_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7551 a_22181_24533# a_22015_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7553 vccd1 _1860_.CLK a_9135_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7554 vccd1 _1830_.CLK a_15794_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7555 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7557 a_4248_5263# _1801_.Y a_3945_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7558 vssd1 _1823_.CLK a_24591_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7559 vssd1 _1763_.A2 a_5086_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X7560 vccd1 _1149_.A1 a_18239_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7561 a_1945_8207# _1786_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7562 a_25559_21482# _1699_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7564 _1158_.X a_9879_12675# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7566 vssd1 _1088_.B a_14373_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7567 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7569 a_15419_2767# a_14637_2773# a_15335_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7570 a_19487_2388# _1740_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7571 _1681_.X a_21643_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7573 vccd1 a_9742_4511# a_9669_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7574 vccd1 a_7626_4511# a_7553_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7575 _0930_.A a_6559_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7576 vccd1 _1907_.CLK a_9779_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7579 a_16849_26159# _1840_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7581 a_17627_15307# _0964_.A a_17541_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7583 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI a_9128_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7584 a_15833_24527# _1895_.Q a_15749_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7585 vccd1 a_10202_29535# a_10129_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7586 a_8807_17999# a_9195_17973# _1074_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7587 a_11241_14191# _1132_.A a_11159_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7588 vccd1 fanout24.A a_26891_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7589 vssd1 a_22879_26703# a_23047_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7590 vccd1 a_4590_25183# a_4517_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7592 a_11601_25071# a_11435_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7593 a_4621_2223# a_4351_2589# a_4531_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7594 a_4753_10089# _1086_.Y a_4669_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7595 a_1975_30287# _1242_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X7596 a_10100_5263# _1140_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7597 a_25398_8207# a_25125_8213# a_25313_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7598 a_8498_20541# _1232_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7599 vccd1 a_23167_14954# _1985_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7600 vccd1 a_27739_2491# a_27655_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7602 a_15143_7119# a_14361_7125# a_15059_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7603 a_2639_3677# a_1775_3311# a_2382_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7604 vssd1 _1086_.Y a_6743_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X7605 _1484_.B a_15207_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X7606 _1325_.B1 a_5269_13367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7607 vssd1 a_25623_13371# a_25581_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7609 vccd1 _1218_.B a_4709_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7611 a_17762_28879# a_17323_28885# a_17677_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7612 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7613 vssd1 a_12575_1501# a_12743_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7614 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_9312_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7615 a_16376_30761# a_16127_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7616 a_4149_1685# a_3983_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7617 a_7090_1501# a_6817_1135# a_7005_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7618 vccd1 _1242_.A1 a_5087_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X7619 a_27314_2335# a_27146_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7620 a_18324_9615# _1112_.A1 a_17749_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X7621 a_15741_3311# a_15575_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7623 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7624 a_23167_14954# _1723_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7625 _1780_.B1 a_4259_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7627 a_6559_12559# _1234_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7628 a_10195_13268# _1558_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7629 a_27548_5487# a_27149_5487# a_27422_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7631 a_4863_23413# _1285_.B1 a_5061_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7632 _1328_.S a_6847_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X7634 a_23005_3145# a_22015_2773# a_22879_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7635 a_16021_23983# _1431_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7636 vssd1 a_14345_24129# _1056_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X7637 a_7635_23555# _0921_.A a_7563_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7638 a_25198_2335# a_25030_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7639 vssd1 a_3210_27765# a_3168_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7641 a_13275_17024# _1839_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7642 a_27314_2335# a_27146_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
R13 vccd1 temp1.capload\[10\].cap_40.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7643 a_17316_27247# temp1.dac.vdac_single.einvp_batch\[0\].vref_55.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7644 a_14594_15529# _1094_.X a_14345_15425# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7645 vssd1 a_10167_4667# a_10125_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7646 a_14319_7691# _0935_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7647 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7649 a_15330_12559# _1103_.D1 a_15081_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X7650 a_5816_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7651 vssd1 a_1828_14709# _1311_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X7652 vccd1 _1132_.A a_14287_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7653 a_21407_8029# a_20543_7663# a_21150_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7654 vccd1 _1192_.X a_14537_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7656 a_14328_4649# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7657 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7658 vccd1 a_14894_16479# a_14821_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7659 a_15483_15823# _1024_.X a_15737_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7660 a_20775_27412# _1492_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7661 vssd1 _2007_.Q _1053_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X7662 vssd1 _1047_.C a_14441_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7663 vccd1 _2008_.Q _1772_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7664 a_22178_6941# a_21905_6575# a_22093_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7665 a_22185_29423# _1869_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7666 a_16105_24847# _1474_.B a_15667_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7667 a_10643_8207# a_9945_8213# a_10386_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7668 vccd1 _1762_.A a_9282_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X7669 a_9742_31029# a_9574_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7670 vccd1 _1841_.CLK a_15023_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7671 a_20982_23261# a_20709_22895# a_20897_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7673 a_5278_22717# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7674 a_3137_2773# a_2971_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7675 vssd1 fanout24.A a_26707_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7676 vssd1 a_3761_9269# _1208_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7678 vssd1 a_23047_2741# a_23005_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7680 vssd1 _1073_.A2 a_17301_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X7682 _0925_.A2 _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7684 vccd1 _0935_.X a_16863_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7685 _1723_.X a_22195_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X7686 a_13455_4765# a_13275_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7688 a_8325_10901# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7689 a_10386_29941# a_10218_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7690 vssd1 _1150_.A2 a_17180_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7691 _1887_.Q a_28015_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7692 a_8025_22717# a_7755_22351# a_7935_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7694 vccd1 a_11455_3579# a_11371_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7695 a_5087_29967# _1242_.B1 _1243_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X7697 _1048_.X a_18519_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7698 vccd1 a_26267_13621# a_26183_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7699 a_22101_32463# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7700 vssd1 a_9779_19087# _1860_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7701 a_27456_10927# a_27057_10927# a_27330_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7702 a_25401_13653# a_25235_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7705 vssd1 a_11953_11073# _1050_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X7706 a_25949_21807# a_24959_21807# a_25823_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7707 a_10938_16341# a_10791_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X7709 a_11759_32362# _1467_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7710 _1497_.X a_18560_22467# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X7711 a_11030_3423# a_10862_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7714 vccd1 _1855_.CLK a_13459_24533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7716 a_15265_21237# _1077_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7717 vccd1 _1999_.CLK a_14379_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7718 a_12978_27791# a_12801_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7720 a_15299_8751# _1059_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7721 a_5455_27791# _0913_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7723 a_25455_1501# a_24591_1135# a_25198_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7725 a_26099_24527# a_25401_24533# a_25842_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7726 vssd1 a_4351_22359# _1337_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7727 a_14894_30623# a_14726_30877# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7728 vssd1 a_25198_27359# a_25156_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7729 vssd1 _0965_.A2 a_19049_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7730 vccd1 _1690_.A_N a_23487_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X7731 a_20897_2223# _1944_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7732 a_12843_15645# a_12061_15279# a_12759_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7733 a_23013_2223# _1636_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7734 vssd1 a_24151_8181# a_24109_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7735 a_4167_8527# _1177_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7736 a_14747_12015# _1025_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7738 _1138_.C1 a_20267_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7739 _0999_.X a_16863_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X7742 a_13821_9615# _1801_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7743 a_10399_24527# a_9871_24527# _1308_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7744 _0985_.X a_15575_19881# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7746 a_19878_1501# a_19439_1135# a_19793_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7747 a_7553_4765# a_7019_4399# a_7458_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7748 a_1941_28335# a_1775_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7749 a_12061_19087# a_11895_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X7750 a_10202_29535# a_10034_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7752 a_24205_21263# a_23671_21269# a_24110_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7753 _1894_.Q a_25623_28603# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7754 vssd1 _2003_.Q a_7571_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7755 a_10055_21376# _1903_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7756 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7757 a_13120_6825# _1065_.X a_13018_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X7758 a_12679_31764# _1473_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7759 vccd1 _0923_.Y a_1769_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X7760 _1091_.B1 a_15207_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7761 _0983_.X a_10147_26409# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7762 a_12659_29789# a_11877_29423# a_12575_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7763 a_11865_5487# _1067_.B a_11793_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7764 a_8395_12559# _1052_.B1 a_8177_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X7765 a_8723_4074# _1566_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7766 _1192_.A2 a_15411_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7767 _1974_.Q a_25255_15797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7769 vccd1 _0983_.A2 a_10413_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7770 _1187_.X a_15299_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7771 _1182_.B a_25623_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7772 a_20537_9661# a_20267_9295# a_20447_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7773 a_6277_11177# _1234_.A1 _1797_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7774 vccd1 _1242_.A2 a_6230_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7775 vssd1 _0918_.A _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X7777 a_8785_20473# _1232_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7778 a_20911_16911# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7779 a_1827_32117# _1337_.A0 a_2036_32509# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X7780 a_2489_17455# _1250_.A1 a_2143_17705# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7781 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7782 vccd1 a_23903_19796# _1387_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7783 vccd1 _1985_.CLK a_24223_15829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7784 a_26870_13469# a_26431_13103# a_26785_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7786 a_23903_26922# _1341_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7788 a_11953_11073# _1044_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7790 a_9220_29199# _1347_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7791 a_13360_27247# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X7792 a_15514_1385# _1607_.B a_15432_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7793 a_10471_7828# _1362_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7794 a_23266_27359# a_23098_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7795 vssd1 a_2471_22869# _1771_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7796 a_22369_1135# _1957_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7798 a_26479_1300# _1616_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7799 vccd1 _1010_.A a_16495_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7800 a_12778_10357# a_12610_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X7802 vccd1 _0966_.A2 a_15005_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7803 _1353_.A a_5271_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7804 a_1757_2223# a_1591_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7806 vccd1 a_25087_15823# a_25255_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7807 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_16376_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7808 a_15887_29789# a_15189_29423# a_15630_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7810 a_7749_23145# a_7561_22941# a_7667_22901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7811 a_17845_22717# _1870_.Q a_17773_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7812 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7813 a_27517_12381# a_26983_12015# a_27422_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7814 vssd1 _0916_.A a_3983_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7815 a_25030_15645# a_24757_15279# a_24945_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7816 a_4760_5737# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7818 a_25064_9673# a_24665_9301# a_24938_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7819 a_2382_28447# a_2214_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7820 vccd1 _1347_.Y a_8767_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X7821 vssd1 a_14139_1679# a_14307_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7822 a_8062_9411# _1537_.B a_7980_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7823 vccd1 _1374_.A_N a_11803_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X7824 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7825 vssd1 a_2807_4667# a_2765_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7826 vssd1 _1744_.B a_19893_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7827 a_12027_20495# a_11711_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X7828 _1629_.X a_17180_2883# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7829 vccd1 _1059_.B a_17538_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X7830 _1810_.A2 a_6600_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7831 a_25198_28447# a_25030_28701# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7832 a_25524_21807# a_25125_21807# a_25398_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7833 vccd1 a_26819_4667# a_26735_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7834 a_12512_31055# a_12263_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X7835 a_21073_29257# a_20083_28885# a_20947_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7836 a_22181_2773# a_22015_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7838 vssd1 a_21115_27765# a_21073_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7839 a_12613_25621# a_12447_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7840 _0981_.B a_9894_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7841 vssd1 _2023_.CLK a_1591_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7842 vssd1 a_12815_9295# _1459_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7843 a_19899_19087# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7844 _1614_.A a_10464_1385# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X7845 a_8447_10004# _1563_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7846 a_13077_29967# _1456_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7847 vssd1 _1850_.CLK a_3983_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7850 vssd1 a_27590_5599# a_27548_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7851 a_13875_23658# _1421_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7852 a_17221_18793# _1832_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7853 vssd1 a_27295_6941# a_27463_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7854 io_out[4] a_4220_21959# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7855 vccd1 a_20315_25834# _1893_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7857 a_9656_16367# a_9613_16600# a_9584_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X7858 a_8102_30511# a_7925_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7859 vccd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7860 a_15285_25615# _1900_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7861 a_23190_22351# a_22751_22357# a_23105_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7862 _1094_.X a_12907_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X7863 a_25455_27613# a_24591_27247# a_25198_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7864 vccd1 _1277_.B a_4899_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7865 a_15620_6351# _0963_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7866 vssd1 _1800_.A2 a_4805_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X7867 vccd1 a_2103_31573# _1329_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X7868 vccd1 _1173_.X a_7295_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X7870 a_17727_1679# a_16863_1685# a_17470_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7871 vssd1 io_in[1] a_2327_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7875 vccd1 _0974_.A2 a_20758_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X7876 a_26479_11690# _1715_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7877 _1469_.A a_14972_26819# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7879 _1829_.Q a_21575_23163# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7881 temp1.capload\[10\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7882 vssd1 a_11711_25615# _1855_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R14 temp1.capload\[7\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7883 _1791_.Y a_7189_13408# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X7885 vssd1 a_6927_17999# _1764_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7886 a_20407_24746# _1414_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7887 a_22963_26703# a_22181_26709# a_22879_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7888 _0984_.A2 a_12295_20747# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7889 a_3873_7125# a_3707_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7890 vssd1 a_18940_12533# _0975_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X7891 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9016_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X7893 _0921_.B a_3983_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7894 vssd1 a_8307_14191# _1544_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7895 a_5625_2223# _1356_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7896 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4160_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X7897 vccd1 temp1.capload\[14\].cap_44.LO temp1.capload\[14\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7898 vssd1 a_28015_3579# a_27973_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7900 _1063_.B a_19735_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7901 a_24665_9301# a_24499_9301# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7902 vccd1 a_3635_27765# a_3551_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7903 vccd1 a_25823_22173# a_25991_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7904 a_11041_18543# _2004_.Q a_10969_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X7908 _0964_.A a_13183_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7909 a_25156_17455# a_24757_17455# a_25030_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7910 vccd1 _1332_.Y a_6463_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7911 a_25309_3311# a_25143_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7912 a_9176_10089# _1198_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7913 vccd1 _1459_.A a_23671_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7914 vccd1 a_3007_1679# a_3175_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7916 vccd1 a_8546_1653# a_8473_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7917 vssd1 a_21886_26271# a_21844_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7918 a_20407_2986# _1732_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7919 vssd1 a_17470_1653# a_17428_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7920 a_20046_31711# a_19878_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7921 a_10349_25045# _1274_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7922 a_4715_7913# _1159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7923 vccd1 _1532_.A a_9135_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7924 vssd1 a_12778_10357# a_12736_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7925 a_26502_23261# a_26063_22895# a_26417_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7926 vssd1 _1218_.B a_6600_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X7928 vccd1 a_25750_29535# a_25677_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7932 a_25539_9117# a_24757_8751# a_25455_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7933 _1685_.A_N a_21187_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7934 vccd1 _1269_.A1 a_9227_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7935 a_28043_16042# _1705_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7936 vccd1 a_26099_4943# a_26267_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7937 a_27655_9117# a_26873_8751# a_27571_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7939 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_7790_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7940 _1385_.A a_20860_19203# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7941 vssd1 fanout21.X a_25143_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7942 a_22073_12533# _1153_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X7943 _1492_.A a_18607_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7944 a_26785_17455# _1525_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7945 vssd1 a_7479_17277# _1139_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X7946 vccd1 _1349_.A a_12631_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7947 a_20775_30186# _1485_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7948 io_out[0] a_1643_21781# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7949 vccd1 _1768_.A a_7295_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7950 vccd1 _1782_.A a_9503_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X7951 vssd1 a_10667_16885# _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7952 a_25087_15823# a_24223_15829# a_24830_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7953 a_15327_4943# a_14545_4949# a_15243_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7954 _1274_.A _1242_.B1 a_7479_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7955 vccd1 a_24278_21237# a_24205_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7956 _1072_.X a_11711_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7957 _1713_.X a_27347_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X7958 _0998_.A2 a_21575_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7959 a_16863_8320# _1146_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7962 vccd1 _1834_.Q a_17904_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X7963 _0922_.Y _0921_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7964 vccd1 _1113_.C a_17171_16395# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7965 vccd1 io_in[2] a_1591_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7967 a_2214_7119# a_1941_7125# a_2129_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7968 vssd1 _1164_.A2 a_7749_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X7969 vssd1 _1143_.A a_14655_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7970 a_20004_1135# a_19605_1135# a_19878_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7971 a_16064_19087# _1020_.B1 a_15962_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X7972 _1179_.B1 a_18459_13131# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X7973 vccd1 _1140_.C a_8859_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7974 a_16373_17455# _1833_.Q a_16301_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7975 a_6645_6575# a_6375_6941# a_6555_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7976 vccd1 _0929_.A _0930_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7977 vccd1 fanout20.X a_22659_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7978 _1564_.X a_7843_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X7979 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7980 a_21533_22895# a_20543_22895# a_21407_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7981 a_4526_22057# _1294_.X a_4220_21959# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7982 a_23281_18543# a_22291_18543# a_23155_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7987 _1878_.Q a_27831_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7989 vccd1 _0932_.A a_5455_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7990 _1058_.B a_7683_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7991 vccd1 _1876_.Q a_18642_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X7992 vccd1 fanout33.A a_14287_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7993 vssd1 io_in[7] a_1591_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X7994 a_8301_15055# _1316_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7995 a_25497_9839# _1927_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7996 a_21511_28500# _1483_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7997 vssd1 _1144_.X a_11711_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7998 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7999 a_10777_3311# _1567_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8001 _1371_.A a_8440_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8002 vssd1 a_9828_26935# _1329_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8003 a_12771_3476# _1623_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8004 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8005 a_7935_22351# a_7755_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8006 a_27663_22173# a_26799_21807# a_27406_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8007 a_16439_3677# a_15575_3311# a_16182_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8010 vccd1 a_27399_16042# _1701_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8011 vccd1 _1876_.CLK a_22659_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8012 _1474_.B a_20379_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8013 a_23776_23817# a_23377_23445# a_23650_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8014 a_10817_17483# _0961_.A a_10731_17483# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8015 vccd1 _1274_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8016 a_25214_3855# a_24941_3861# a_25129_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8017 vssd1 a_16623_2589# a_16791_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8018 _0974_.A2 a_28015_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8019 a_19513_31061# a_19347_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8022 vssd1 a_19735_14709# a_19693_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8023 vssd1 a_4314_7093# a_4272_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8024 vssd1 a_23523_11293# a_23691_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8025 _1474_.B a_20379_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8026 a_12150_8207# a_11877_8213# a_12065_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8027 a_26513_31849# _1353_.B _1353_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8028 a_15293_14851# _1104_.C a_15197_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X8030 vccd1 _1242_.A2 a_1841_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8031 vccd1 _1113_.C a_18795_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8032 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_12512_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8033 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8035 _1387_.A a_23391_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X8036 vccd1 _2009_.CLK a_1775_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8037 a_27333_22173# a_26799_21807# a_27238_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8038 vssd1 _1165_.C a_6953_8545# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8040 vccd1 a_12539_7663# _1577_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8041 vccd1 a_25566_8181# a_25493_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8042 a_3517_22351# _0913_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X8043 a_27238_21085# a_26799_20719# a_27153_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8044 vccd1 a_2807_3579# a_2723_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8045 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8046 a_12528_16367# a_12079_16367# a_12226_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8048 a_1757_1135# a_1591_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8049 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8050 _1764_.Y _1764_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8051 vccd1 _1880_.CLK a_24591_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8052 a_11023_18218# _1376_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8053 vccd1 _1073_.A2 a_16209_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8054 a_20039_5162# _1607_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8056 a_9761_27797# a_9595_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8057 _2003_.D _1775_.C1 a_2153_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8058 _1410_.A a_19388_22467# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8060 a_12525_10383# _1848_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8061 vssd1 _1051_.A1 a_8440_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8063 vccd1 fanout21.X a_26707_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8065 a_2382_3423# a_2214_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8066 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8068 a_14641_16367# _1850_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8069 a_10911_19997# a_10129_19631# a_10827_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8070 _1139_.C a_7479_17277# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X8071 vccd1 _1941_.CLK a_18243_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8072 a_22365_20181# a_22199_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8073 vssd1 _2004_.Q a_9963_15939# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8074 a_10141_15939# _2004_.Q a_10045_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X8078 a_17831_30676# _1471_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8079 vccd1 a_13330_29941# a_13257_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8080 a_2957_24527# _1769_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8082 a_4519_9991# _1125_.X a_4669_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X8083 vssd1 a_8548_23413# _1329_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8084 vccd1 a_25623_20987# a_25539_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8085 a_23483_12381# a_23303_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8086 vssd1 _0989_.B2 a_10428_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X8087 a_7834_10089# _1164_.A2 a_7531_9813# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X8089 vssd1 a_5731_12567# _1325_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8090 _1873_.Q a_25623_31867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8092 a_20858_14735# _1824_.Q a_20701_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8093 a_27517_3677# a_26983_3311# a_27422_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8094 a_18233_10749# _0939_.A a_18151_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8095 a_22917_22357# a_22751_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8096 _1073_.A2 a_17171_16395# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X8097 vccd1 _1907_.CLK a_11711_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8098 vccd1 clkbuf_0_net57.X a_2686_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8099 _1116_.C1 a_13643_22464# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8100 a_2777_17999# _0925_.A2 a_2695_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8101 a_24757_6575# a_24591_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8102 vccd1 a_21575_7931# a_21491_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8103 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8104 vccd1 _1474_.A_N a_14287_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8105 a_8473_1679# a_7939_1685# a_8378_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8107 a_25750_29535# a_25582_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8108 a_5136_22583# _2008_.Q a_5278_22390# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8109 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8110 vssd1 a_27590_19743# a_27548_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8112 _1265_.A1 _1263_.A a_12073_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8113 vccd1 a_22346_6687# a_22273_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8114 a_17204_30761# a_16955_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8116 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8117 a_3435_22671# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X8118 _1088_.B a_19275_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8119 vssd1 _1306_.A2 a_6921_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X8120 a_16797_22923# _0961_.A a_16711_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8121 a_8059_2589# a_7277_2223# a_7975_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8122 vssd1 _1768_.A _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8123 a_7657_16617# _1325_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X8124 vccd1 a_19310_17973# a_19237_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8125 a_20571_28701# a_19789_28335# a_20487_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8126 a_5903_19407# _1273_.A1 _1280_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X8127 a_23833_30345# a_22843_29973# a_23707_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8128 a_13599_7828# _1749_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8129 vssd1 a_9735_9514# _1759_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8130 _1132_.A a_10883_21271# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8131 vccd1 _1221_.A _1246_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8132 temp1.capload\[15\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8133 a_24639_18708# _1695_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8134 _1127_.X a_20267_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8139 vssd1 a_12815_19631# _1489_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8140 a_17029_27797# a_16863_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8141 _1973_.Q a_25623_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8142 vssd1 _1766_.A0 a_7939_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8143 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_4252_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8145 _1152_.B a_26267_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8146 _1165_.A a_6467_9001# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X8147 a_13330_29941# a_13162_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8148 vssd1 _1894_.Q a_18789_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8149 vccd1 _2023_.CLK a_1683_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8150 vccd1 _1183_.A2 a_20081_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8151 a_20295_31055# a_19513_31061# a_20211_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8152 a_25589_26703# _1883_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8153 a_8548_23413# _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8154 _1977_.Q a_27463_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8155 vccd1 a_15081_12533# _1104_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8156 a_21936_30511# a_21537_30511# a_21810_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8157 a_23101_3861# a_22935_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8158 vccd1 _1999_.CLK a_10423_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8159 a_2030_6941# a_1591_6575# a_1945_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8160 vccd1 a_13057_8897# _1069_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X8161 a_25447_9295# a_24665_9301# a_25363_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8162 a_8937_29967# a_8760_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8163 a_8719_20541# _0913_.A1 a_8356_20407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8164 _1326_.A3 _1324_.A a_4161_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8165 vccd1 a_4847_25437# a_5015_25339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8166 vccd1 fanout37.A a_20543_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8167 _1658_.X a_10327_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X8168 a_9669_5853# a_9135_5487# a_9574_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8169 _1538_.A a_15800_26819# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8170 vccd1 a_5047_21237# _1294_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8173 vssd1 _1349_.A a_12631_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8174 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_8392_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8175 vssd1 a_7809_18517# _1257_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X8176 a_26969_16367# _1387_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8177 vccd1 a_25623_1403# a_25539_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8178 _1486_.B a_20563_30779# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8179 a_24945_23983# _1972_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8180 _1789_.A1 _1313_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8181 a_10386_1653# a_10218_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8184 vssd1 a_24535_10383# a_24703_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8186 a_10951_24233# a_10423_23983# _1270_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8187 a_26225_20553# a_25235_20181# a_26099_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8188 vccd1 a_20407_24746# _1837_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8189 a_24393_19087# _1826_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8190 _1164_.A2 _1198_.A2 a_8297_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8191 a_6559_12559# _1255_.A1 a_6981_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8192 _1818_.Q a_10627_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8193 a_5354_28335# clkbuf_0_temp1.i_precharge_n.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8194 a_25674_6031# a_25235_6037# a_25589_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8195 a_16175_9514# io_in[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8196 vccd1 a_17102_31711# a_17029_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8197 vccd1 a_23047_31029# a_22963_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8198 _0998_.B2 a_25439_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8199 vssd1 a_2639_3855# a_2807_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8200 vssd1 a_15227_7093# a_15185_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8201 vccd1 _0993_.X a_14453_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8202 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8203 a_8083_17455# _1269_.A1 a_7969_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.1365 ps=1.07 w=0.65 l=0.15
X8204 vccd1 _1141_.C a_13399_17483# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8205 vssd1 _1353_.A _1332_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8206 a_27548_27247# a_27149_27247# a_27422_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8207 a_2214_6031# a_1941_6037# a_2129_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8209 a_23607_22173# a_22825_21807# a_23523_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8210 vccd1 a_17541_15307# _1024_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X8211 a_5177_14441# _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X8212 vssd1 _1841_.CLK a_16495_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8214 _0918_.A a_3983_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8215 a_8675_8207# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8216 vccd1 _1896_.CLK a_20083_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8218 a_20499_23658# _1410_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8219 a_25198_20831# a_25030_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8220 a_11969_17455# _2006_.Q a_11869_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X8221 vccd1 a_17047_17455# _1405_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8222 a_13433_11177# _1197_.B a_13361_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
R15 temp1.capload\[6\].cap_51.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8223 a_2153_25615# _1775_.C1 _2003_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8224 a_25493_8207# a_24959_8213# a_25398_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8225 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.A a_14370_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8226 a_7100_19631# _0909_.A a_6797_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X8227 _1173_.X a_5547_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X8228 vssd1 a_9079_2767# a_9247_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8229 a_9595_8751# _1058_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8230 a_24025_11471# _1966_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
R16 vccd1 temp1.capload\[11\].cap_41.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X8231 a_27038_13215# a_26870_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8232 vssd1 _1202_.Y a_7002_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8233 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8235 vccd1 a_27406_21919# a_27333_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8236 a_10515_12015# _1198_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X8238 vssd1 a_11760_23671# _1346_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8240 _1250_.A1 _1199_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8241 a_5499_22717# _2008_.Q a_5136_22583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8242 vccd1 _1882_.CLK a_22751_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8243 vssd1 a_11023_5162# _1647_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8244 a_10133_8207# _1813_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8246 vssd1 _1873_.CLK a_22015_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8248 a_5187_16911# _1231_.B1 a_4932_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X8249 a_26007_10205# a_25143_9839# a_25750_9951# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8251 a_8785_15974# _0956_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X8253 a_21905_6575# a_21739_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8254 vssd1 _1973_.Q a_28173_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8255 a_19709_3311# a_19439_3677# a_19619_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8256 a_12253_8751# _1010_.A a_12171_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8258 a_18789_27069# a_18519_26703# a_18699_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8259 vssd1 a_23155_18909# a_23323_18811# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8262 a_20223_8426# _1582_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8263 a_6981_12559# _0903_.C _0909_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8265 vccd1 _2009_.CLK a_2051_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8266 vccd1 _1782_.A a_1898_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X8267 vccd1 _1690_.A_N a_27903_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8268 vccd1 _1122_.A1 a_6645_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X8269 _1762_.A a_7755_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8270 _1217_.A3 _1226_.A1 a_5449_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8271 a_25582_26525# a_25143_26159# a_25497_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8273 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8274 vccd1 _1861_.Q a_12752_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8275 vssd1 _1060_.C1 a_13057_8897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X8276 a_5269_13367# _0917_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8277 a_2949_25071# a_1959_25071# a_2823_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8278 a_25677_10205# a_25143_9839# a_25582_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8279 a_4173_14441# _1279_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8280 _1425_.A a_15939_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X8281 a_2047_16617# _1249_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8282 vssd1 _1924_.CLK a_25235_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8283 a_22273_6941# a_21739_6575# a_22178_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8285 a_20867_8426# _1598_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8286 vccd1 _1110_.A a_17323_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8289 vssd1 _1941_.CLK a_20175_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8290 a_12896_22671# _1861_.Q a_12321_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8291 vccd1 fanout20.X a_25787_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8293 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_6828_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8294 a_8385_30511# a_8208_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8296 vssd1 _0956_.C a_7756_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X8297 vssd1 a_25731_11293# a_25899_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8298 vccd1 _2006_.Q a_12079_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8299 a_16911_5162# _1633_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8300 a_20303_5853# a_19439_5487# a_20046_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8301 a_8178_12265# _1084_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X8302 a_6644_5263# _1208_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8303 vccd1 _0929_.A a_5361_11191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X8306 _0987_.Y _0987_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8307 vccd1 a_18114_1247# a_18041_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8308 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_17204_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8309 a_17013_19777# _1024_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X8310 vccd1 _1012_.Y a_7939_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8312 vssd1 a_10202_2335# a_10160_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8313 vccd1 a_17895_1653# a_17811_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8315 a_15115_9408# _1057_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X8316 a_27337_5487# _1728_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8317 vccd1 a_25623_31867# a_25539_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8318 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8321 a_11874_2589# a_11435_2223# a_11789_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8323 vssd1 _1216_.A2 a_4713_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X8324 a_20959_26922# _1553_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8325 io_out[2] a_1643_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8326 vssd1 _0994_.B2 a_15948_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X8327 _1458_.A a_10740_25731# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8328 a_5980_31849# a_5731_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8329 a_13146_12533# a_12978_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8330 a_17677_28879# _1469_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8331 _1186_.C1 a_10331_23145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8333 _0958_.A a_13551_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X8334 a_13432_28585# a_13183_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8335 a_19521_20969# _1184_.C1 a_19439_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8336 vccd1 _1823_.CLK a_24039_19093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8337 a_24945_17455# _1914_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8338 vssd1 _1438_.B a_12176_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X8339 _1034_.Y _1024_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8341 a_24937_15113# a_23947_14741# a_24811_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8342 vccd1 _1112_.A1 a_20999_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8343 vssd1 a_26175_29691# a_26133_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8344 vssd1 a_17930_28853# a_17888_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8345 a_28173_17277# a_27903_16911# a_28083_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8347 vccd1 a_8113_25117# a_8213_25335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X8348 _0918_.A a_3983_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8349 a_9360_18793# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8350 a_13061_7485# _1039_.B a_12989_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8351 a_12801_25615# _1901_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8352 a_4127_22869# _1274_.A a_4345_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X8353 _1111_.B a_23691_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8354 vssd1 _1344_.B a_4627_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8355 a_25800_23817# a_25401_23445# a_25674_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8357 vssd1 a_3983_19631# _0918_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8358 a_2156_6575# a_1757_6575# a_2030_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8359 vssd1 _1156_.Y a_7573_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X8360 _1431_.A a_13040_23555# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8361 vssd1 _1836_.Q a_19709_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8362 a_20390_9001# _1577_.B a_20308_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8363 a_2408_25615# _0913_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8364 a_5588_6825# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8365 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8366 a_7009_11177# _1084_.C1 _1086_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8367 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4988_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8368 a_25842_13621# a_25674_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8369 a_19609_29967# a_19432_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8370 vccd1 _1821_.Q a_14776_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8371 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4075_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8372 a_2524_25071# a_2125_25071# a_2398_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8373 a_17217_1679# _1624_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8375 a_17704_29423# a_17305_29423# a_17578_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8376 vccd1 a_2382_7093# a_2309_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8377 vccd1 a_10202_27765# a_10129_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8378 vccd1 _1103_.A1 a_15512_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X8379 a_24811_28879# a_23947_28885# a_24554_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8380 a_25800_6409# a_25401_6037# a_25674_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8381 a_27337_12015# _1978_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8382 a_2217_23983# a_2051_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8383 _1823_.Q a_27831_20987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8384 vccd1 _1968_.Q a_22195_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8385 a_12318_13621# a_12150_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8386 a_15081_22325# _1116_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X8388 a_15656_12879# _1103_.A1 a_15081_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8389 a_17029_31965# a_16495_31599# a_16934_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8390 vccd1 _1272_.A2 a_1841_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8391 vccd1 _0952_.A1 a_17139_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X8392 vssd1 a_26479_11690# _1716_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8393 vccd1 _1775_.A2 _0923_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8394 a_25674_13647# a_25401_13653# a_25589_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8395 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8396 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8397 a_14901_19631# _1869_.Q a_14829_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8398 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_15750_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8401 vssd1 a_19735_1653# a_19693_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8402 a_25674_4943# a_25235_4949# a_25589_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8405 a_19191_3855# a_18409_3861# a_19107_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8406 a_17029_12559# _1890_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8407 a_20315_26922# _1536_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8409 a_2129_4399# _1783_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8411 vccd1 a_11563_31965# a_11731_31867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8412 a_24481_28879# a_23947_28885# a_24386_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8413 vccd1 _1489_.A_N a_18427_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8414 a_13054_25589# a_12886_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8415 vccd1 a_7755_21263# _1762_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8416 _1230_.B1 _1249_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8417 vccd1 _0939_.A a_14471_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8418 a_20421_10927# _0973_.B a_20349_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8419 _0961_.A a_15299_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8420 vccd1 a_16607_3579# a_16523_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8421 a_23607_4943# a_22825_4949# a_23523_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8422 _1880_.CLK a_15886_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8423 vssd1 _1876_.CLK a_22015_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8424 a_12150_13647# a_11877_13653# a_12065_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8425 a_19521_7663# _1010_.A a_19439_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8426 _1038_.D1 a_16035_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8427 vssd1 _1882_.CLK a_26063_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8428 a_17673_1135# a_17507_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8429 vssd1 _1816_.CLK a_7019_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8430 a_9749_8751# _1058_.B a_9677_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8432 vssd1 a_25382_16479# a_25340_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8433 vccd1 a_25382_3829# a_25309_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8434 _1427_.A a_18239_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8435 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8437 vssd1 a_15115_5487# _1830_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8440 _1816_.CLK a_3983_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8441 vssd1 _1316_.X a_6363_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X8442 a_16182_3423# a_16014_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8443 vssd1 _1459_.A a_17047_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X8444 vssd1 a_5871_1898# _1816_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8445 vssd1 a_20885_16341# _1179_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8446 a_5639_25615# _1305_.B _1306_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8447 a_8031_17999# _1764_.A a_8449_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8448 a_17470_1653# a_17302_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8449 a_7803_6740# _1752_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8451 vccd1 a_23047_1403# a_22963_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8452 vssd1 _1775_.A2 a_6600_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8453 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_1860_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8454 a_24512_15113# a_24113_14741# a_24386_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8455 a_9949_2223# _1657_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8456 a_18041_1501# a_17507_1135# a_17946_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8457 vssd1 _1037_.B a_18237_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8458 a_15749_24527# _1180_.X a_15667_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8460 a_10693_8751# a_10423_9117# a_10603_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8461 a_17861_31055# _1467_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8462 vssd1 _1837_.Q a_18513_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8463 vccd1 a_23155_24349# a_23323_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8464 a_8395_22057# _1270_.A a_8177_21781# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X8465 a_8325_10901# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8466 a_16661_26159# a_16495_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8469 vssd1 a_20867_8426# _1599_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8470 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8471 vccd1 a_25455_2589# a_25623_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8473 vccd1 _1855_.CLK a_11435_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8474 a_19709_22895# a_19439_23261# a_19619_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8475 a_4669_10089# _1324_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X8476 a_23358_22325# a_23190_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8477 vccd1 _1242_.A2 a_5087_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8478 a_8569_27247# a_8392_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8479 vccd1 _1133_.C a_18519_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8480 vccd1 _2023_.CLK a_1775_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8482 vssd1 a_26670_25183# a_26628_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8484 a_5357_3087# a_5165_2828# _1808_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X8485 a_4061_7119# _2020_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8486 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8487 a_25401_20181# a_25235_20181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8489 a_21181_23983# a_20911_24349# a_21091_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8490 vssd1 a_12502_15391# a_12460_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8491 a_1674_28879# clkbuf_0_temp1.i_precharge_n.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8492 _1116_.D1 a_13183_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8493 _1637_.X a_16904_3971# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8494 vccd1 _0918_.A a_10041_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8495 a_25198_5599# a_25030_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8496 _1153_.A a_18059_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8497 a_7104_27247# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8499 a_24719_1679# a_23855_1685# a_24462_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8500 a_18072_31433# a_17673_31061# a_17946_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8501 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8502 vccd1 a_25439_17973# a_25355_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8503 vccd1 _1071_.B1 a_13433_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X8504 a_10839_10602# _1436_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8505 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_6559_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8506 vssd1 clkbuf_0_net57.X a_1674_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8508 a_23190_22351# a_22917_22357# a_23105_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8509 a_24573_18005# a_24407_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8510 vssd1 a_21695_17620# _1826_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8511 a_23155_24349# a_22457_23983# a_22898_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8512 vccd1 _2023_.CLK a_1591_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8514 vccd1 a_3983_19631# _0918_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8515 vccd1 _1021_.A a_13275_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8516 vssd1 _1074_.C a_14405_7691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8517 vccd1 _1177_.Y a_1857_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8518 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8520 _1607_.B a_9135_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8521 a_10413_23145# _1859_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8522 vccd1 _2005_.Q a_12226_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X8523 _1024_.D1 a_17415_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8525 a_12771_21482# _1549_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8526 vccd1 _1135_.B a_20447_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8527 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X8528 a_17727_1679# a_17029_1685# a_17470_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8529 a_26099_6031# a_25401_6037# a_25842_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8531 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13432_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8532 a_13464_5487# _0993_.X a_12973_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X8534 vccd1 fanout21.X a_24407_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8535 a_7656_11471# _1164_.A2 _1279_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X8536 a_10190_5263# _0989_.A2 a_10100_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X8537 a_12000_2223# a_11601_2223# a_11874_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8538 a_2103_13647# _1246_.B2 a_1641_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X8539 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4903_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8540 vssd1 _1049_.C1 a_17841_17601# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X8541 vssd1 _1123_.X a_6651_11587# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8542 a_10399_24527# _0921_.B a_10041_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8544 vssd1 a_24462_1653# a_24420_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8545 a_12701_29423# a_11711_29423# a_12575_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8546 a_7442_17429# a_7295_17455# a_8083_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X8547 a_2983_23217# _0958_.A a_2471_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X8548 a_6406_13353# _1316_.X a_6324_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8549 vssd1 a_15963_25589# a_15921_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8550 vccd1 _1882_.CLK a_26431_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8551 a_9282_16341# _1764_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X8552 vccd1 a_14335_2388# _1935_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8553 _1146_.B a_20471_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8554 _1674_.A a_20907_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X8555 a_19061_10749# _0952_.A1 a_18979_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8556 _1184_.B1 a_17999_16395# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X8557 a_18869_1685# a_18703_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8558 a_25639_16733# a_24775_16367# a_25382_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8559 vssd1 _0921_.A _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8561 a_15925_2223# a_15759_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8562 a_27590_26271# a_27422_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8563 a_4198_4649# _1801_.B a_4116_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8565 a_18850_2741# a_18682_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8566 a_5980_30761# a_5731_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8567 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_12482_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8568 a_27663_22173# a_26965_21807# a_27406_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8569 a_23098_11293# a_22659_10927# a_23013_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8570 a_7381_13103# _1314_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8571 vccd1 _0939_.A a_15299_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8572 a_9275_24746# _1547_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8573 vccd1 a_10839_20884# _1851_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8574 vccd1 a_13599_29588# _1469_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8575 vssd1 a_27847_26525# a_28015_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8576 vssd1 a_2198_6687# a_2156_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8577 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8578 a_18513_24893# a_18243_24527# a_18423_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8579 a_2490_24349# a_2051_23983# a_2405_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8580 vccd1 a_26283_18909# a_26451_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8581 a_20298_22467# _1506_.B a_20216_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8582 vccd1 _1328_.S a_3087_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X8583 vssd1 _1071_.B1 a_12500_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X8584 a_15410_12559# _1101_.X a_15330_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X8585 _0911_.A a_2623_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8586 a_17625_22923# _0964_.A a_17539_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8587 vssd1 _1801_.B a_3861_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8588 a_25773_18543# _1971_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8589 vssd1 _1830_.CLK a_25235_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8591 vssd1 a_23358_22325# a_23316_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8593 _1261_.A1 a_2715_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8594 a_16382_25071# a_16205_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8595 vssd1 a_15319_16635# a_15277_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8596 a_17811_29967# a_17029_29973# a_17727_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8597 vssd1 _1876_.CLK a_22659_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8598 vccd1 a_3835_2767# a_4003_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8599 vccd1 a_27859_30186# _1456_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8600 a_17029_18005# a_16863_18005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8602 a_8038_10927# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8603 a_1766_26159# clkbuf_1_1__f__0380_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8604 a_21235_25236# _1511_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8605 a_16021_23983# _1431_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8607 vssd1 a_2715_7931# a_2673_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8609 vccd1 a_24554_28853# a_24481_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8610 a_11874_25437# a_11435_25071# a_11789_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8611 _1337_.S a_4351_22359# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8613 vccd1 a_7111_25071# _1242_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8614 a_1657_10901# _1170_.B1 a_1814_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X8615 a_12759_15645# a_11895_15279# a_12502_15391# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8616 a_13357_17277# _1021_.A a_13275_17024# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8617 a_12637_15823# _1820_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8619 vccd1 _1010_.A a_14747_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8620 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8621 _1305_.B a_6559_24640# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8622 vccd1 a_17727_27791# a_17895_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8623 vccd1 a_2382_6005# a_2309_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8625 a_4973_25071# a_3983_25071# a_4847_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8627 a_25581_6575# a_24591_6575# a_25455_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8628 vssd1 a_22587_31867# a_22545_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8629 _1308_.B a_9871_24527# a_10399_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8630 vssd1 _1090_.C a_16373_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8631 a_25800_5321# a_25401_4949# a_25674_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8633 vssd1 _2009_.CLK a_1775_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8634 a_10270_14441# _1537_.B a_10188_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8635 vssd1 _1898_.Q a_14557_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8636 vccd1 _1690_.A_N a_27627_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8637 a_6223_3339# _1291_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8638 _1226_.B1 a_6644_5263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8639 _1486_.X a_13455_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8640 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9220_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8641 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13360_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8642 a_1757_1135# a_1591_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8644 vssd1 _1880_.CLK a_24591_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8645 a_15097_25621# a_14931_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8646 vssd1 _1876_.CLK a_22291_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8647 vssd1 _1140_.C a_10945_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X8648 a_19793_1135# _1945_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8649 a_17814_24233# _1133_.X a_17565_24129# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8651 a_10218_8207# a_9779_8213# a_10133_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8652 vssd1 a_25087_15823# a_25255_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8653 a_25750_3423# a_25582_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8654 vssd1 _1024_.A2 a_19980_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X8655 a_3919_2767# a_3137_2773# a_3835_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8656 vccd1 _1775_.C1 a_8215_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8658 a_7025_13647# _0930_.A a_6610_13879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X8660 a_12035_2986# _1617_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8661 a_18850_2741# a_18682_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8662 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8663 _1574_.X a_19480_15529# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8664 a_27149_27247# a_26983_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8665 a_8027_18793# _0925_.A2 a_7809_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X8667 a_5392_23983# _1294_.B1 a_5301_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X8668 a_22580_24905# a_22181_24533# a_22454_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8669 a_12299_2589# a_11601_2223# a_12042_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8670 a_25214_16733# a_24941_16367# a_25129_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8671 vccd1 _1353_.A a_26513_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8672 vccd1 _1068_.A1 a_14410_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X8674 a_15365_14851# _1095_.X a_15293_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8675 _1633_.X a_17319_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8676 a_9350_24233# _1422_.B a_9268_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8678 vccd1 a_15457_6005# _1008_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X8679 vccd1 _1217_.A3 a_4351_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8681 a_2677_1679# a_2143_1685# a_2582_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8682 a_26229_22895# a_26063_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8683 _1184_.X a_19439_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X8684 a_17262_2883# _1607_.B a_17180_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8685 vccd1 _1083_.A a_4842_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X8686 vssd1 a_27923_11195# a_27881_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8687 a_13713_30345# a_12723_29973# a_13587_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8688 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_13275_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8689 a_9786_23478# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8690 a_16005_22895# _1880_.Q a_15933_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8691 a_20885_16341# _1024_.A2 a_21042_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X8692 _1210_.B _1165_.A a_7637_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X8693 vssd1 _0992_.A2 a_7749_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8694 vssd1 _1221_.A a_2644_11587# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8695 _1855_.Q a_11731_31867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8696 vccd1 a_27095_25339# a_27011_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8697 vccd1 a_15163_2388# _1643_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8698 vssd1 _1325_.A2 a_6639_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X8699 vssd1 _0984_.A2 a_12057_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8700 _1121_.A1 a_5199_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8702 vccd1 _1855_.CLK a_12447_25621# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8703 vssd1 a_26267_20149# a_26225_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8705 vccd1 a_20471_5755# a_20387_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8706 a_4973_2057# a_3983_1685# a_4847_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8707 a_25769_4943# a_25235_4949# a_25674_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8708 a_23098_4943# a_22659_4949# a_23013_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8710 a_18147_4765# a_17967_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X8711 a_22238_14735# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X8713 a_12705_12565# a_12539_12565# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8714 _1294_.X a_5203_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8715 vccd1 _1011_.A1 a_7843_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8717 vssd1 _1314_.X a_9253_14219# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8718 a_23799_3855# a_22935_3861# a_23542_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8719 a_20727_6031# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8720 vssd1 a_25842_12533# a_25800_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8721 a_19470_21379# _1506_.B a_19388_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8722 a_24987_19087# a_24205_19093# a_24903_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8723 a_7699_3855# a_6835_3861# a_7442_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8724 a_19163_12879# _0974_.A2 a_19069_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X8727 vccd1 _1090_.C a_19439_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X8729 vssd1 a_4497_7637# _1170_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X8730 vccd1 _1794_.Y a_5451_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8731 _1580_.A a_19388_8323# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8732 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8734 vssd1 _1850_.CLK a_8307_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X8735 _1853_.Q a_15319_30779# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8736 vssd1 _1764_.A _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8737 _1975_.Q a_25623_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8738 a_14557_22895# a_14287_23261# a_14467_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X8739 a_13304_14441# _1035_.X a_13202_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X8740 _1145_.B2 a_10811_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8741 a_5496_9001# _1279_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8744 _1855_.CLK a_11711_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8745 vccd1 a_18107_21972# _1829_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8749 vccd1 _1342_.Y a_7755_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8750 vssd1 a_8803_1679# a_8971_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8751 a_10643_1679# a_9779_1685# a_10386_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8752 a_26099_4943# a_25401_4949# a_25842_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8753 a_4351_12559# _1217_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8754 a_22879_26703# a_22015_26709# a_22622_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8755 vccd1 clkbuf_1_1__f__0380_.A a_1766_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8756 a_2009_21583# _1242_.A2 a_2199_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8757 temp1.capload\[14\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8759 vssd1 a_23542_3829# a_23500_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8760 a_24945_5487# _1593_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8762 vssd1 a_7442_3829# a_7400_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8764 a_3761_9269# _1175_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X8765 a_1814_11177# _1170_.B2 a_1657_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8766 vssd1 a_19567_17999# a_19735_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8767 vccd1 a_21327_1300# _1990_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8768 _1008_.X a_14839_10499# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X8769 _1234_.A2 a_5455_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8771 a_5349_3616# _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8772 vssd1 a_18383_3476# _1941_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8773 vssd1 _1532_.A a_12815_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X8774 a_27057_10927# a_26891_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8775 vccd1 a_26267_24501# a_26183_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8776 vssd1 _1532_.A a_4627_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X8777 vccd1 _1010_.A a_17139_11584# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8779 a_27498_28447# a_27330_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8782 vccd1 a_2807_3829# _1304_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8784 a_15710_6351# _0994_.A2 a_15620_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X8785 a_22549_26703# a_22015_26709# a_22454_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8786 a_17381_7093# _1064_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X8788 a_22270_29789# a_21831_29423# a_22185_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8789 a_18048_16143# _1834_.Q a_17473_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8792 vssd1 a_27755_28701# a_27923_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8793 vssd1 a_15633_11445# _1120_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X8795 a_14323_24527# a_13625_24533# a_14066_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8796 a_19065_20495# _1884_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X8798 a_15882_26819# _1537_.B a_15800_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8799 a_2471_22869# _0958_.A a_2680_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8800 a_19497_18689# _1138_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X8801 vssd1 a_10386_1653# a_10344_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8803 _1451_.B a_10811_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8804 vssd1 a_12575_29789# a_12743_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8805 _1186_.X a_11987_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X8806 _1414_.A a_19619_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8807 vccd1 _2006_.Q a_10865_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X8809 vccd1 a_11685_9813# _1008_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X8810 vccd1 a_22063_22570# _1882_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8811 _1141_.C a_10667_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8812 a_9779_11791# _1104_.X _1122_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8813 a_10313_29967# a_9779_29973# a_10218_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8815 _1781_.Y _1781_.B a_13349_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X8816 a_23649_2223# a_22659_2223# a_23523_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8817 a_7932_25935# _1342_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8818 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A a_8004_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8820 temp1.capload\[8\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8821 _1175_.Y _1175_.B2 a_7939_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8822 _1075_.C a_10938_16341# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8823 a_17171_16395# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8824 a_2686_15823# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8825 vssd1 _1052_.B1 _1324_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8827 vccd1 a_8447_6740# _1812_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8828 vccd1 _1110_.A a_11711_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8829 a_14655_18115# _1134_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8830 vssd1 _1907_.CLK a_9135_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8831 a_21905_6575# a_21739_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8833 vssd1 _1080_.B a_18468_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8834 a_15496_31433# a_15097_31061# a_15370_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8835 _0930_.B _0929_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8836 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X8838 vssd1 a_15299_21807# _1021_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8840 a_22622_31029# a_22454_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X8841 vssd1 _1849_.CLK a_16113_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8842 _1967_.Q a_28015_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8843 vssd1 _1267_.A1 a_5639_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8844 vssd1 _2009_.CLK a_2051_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8845 a_26785_13103# _1707_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8846 a_20437_28879# _1870_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X8847 _1775_.B1 a_7847_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X8850 vccd1 _1474_.A_N a_7203_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X8851 a_4988_31375# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X8852 vccd1 a_19671_25834# _1876_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8853 a_10344_8585# a_9945_8213# a_10218_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8854 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_4252_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8855 a_5635_18793# _1325_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8856 vssd1 _1321_.C a_6309_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X8857 _1198_.A2 a_9779_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8858 a_9301_31061# a_9135_31061# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8860 vssd1 a_20230_28447# a_20188_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8861 _1517_.A a_20584_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8862 vccd1 _1941_.CLK a_15575_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8863 a_17749_9269# _1112_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X8864 vssd1 a_6610_13879# _1263_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8865 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12532_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X8866 a_12557_16600# _2004_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X8867 vccd1 a_20211_31055# a_20379_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8868 vccd1 _1880_.CLK a_16205_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8869 vssd1 _1802_.X a_4248_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8870 a_22454_31055# a_22181_31061# a_22369_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8872 a_3145_8751# _1263_.A a_3063_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8873 a_9644_23671# _0911_.A a_9786_23478# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8874 a_15477_20291# _1184_.X a_15381_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X8875 a_10147_14735# _1269_.A1 a_10397_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8876 vssd1 _1896_.CLK a_19347_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8877 a_10593_24233# _0921_.A a_10951_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8878 a_20081_12559# _0958_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X8879 a_22503_31965# a_21721_31599# a_22419_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8880 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8882 a_10493_26159# _1464_.B a_10147_26409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8883 vssd1 a_25623_17723# a_25581_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X8884 a_2581_8585# a_1591_8213# a_2455_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8886 vccd1 a_9999_5853# a_10167_5755# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8888 a_15013_27791# _1486_.B a_14931_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8889 a_1591_24527# _1775_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8890 vccd1 a_12318_1247# a_12245_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8891 a_23443_7338# _1675_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8892 a_20308_9001# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8893 a_8556_31055# a_8307_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X8894 _1310_.Y _1310_.B1 a_5731_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8895 a_20390_21379# _1506_.B a_20308_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8896 a_5451_11471# _1795_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8897 a_22235_30877# a_21371_30511# a_21978_30623# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8898 vssd1 a_2658_27359# a_2616_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8899 vccd1 _1876_.CLK a_25143_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8900 _1775_.C1 a_7387_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8901 vccd1 a_25014_2741# a_24941_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X8902 _1073_.X a_16219_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X8903 vccd1 _1300_.A2 a_3069_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8905 vccd1 _1154_.A1 a_23667_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8907 vssd1 _1879_.Q a_21917_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8908 a_25125_21807# a_24959_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8909 _1670_.A a_22195_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8910 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X8912 a_11299_12180# _1434_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8913 vccd1 _1146_.B a_14410_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X8914 a_9503_8029# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8915 vccd1 a_2971_16367# _0921_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8916 a_25198_6687# a_25030_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8917 vccd1 _1855_.CLK a_9595_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8918 a_22457_27797# a_22291_27797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8919 _0909_.C _1242_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8921 _1277_.A _1217_.B1 a_4351_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X8922 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8923 a_10413_22895# _1817_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8924 vssd1 _0975_.C1 a_18887_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8927 a_14357_21641# a_13367_21269# a_14231_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X8928 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8929 vccd1 a_24887_1653# a_24803_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8930 a_23224_5321# a_22825_4949# a_23098_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8931 vssd1 a_16863_23439# fanout33.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8933 vssd1 _1872_.Q a_18697_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8934 a_22454_2767# a_22181_2773# a_22369_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8935 vssd1 _1061_.B a_22285_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8936 a_14465_9001# _1196_.C a_14369_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X8937 a_10827_19997# a_9963_19631# a_10570_19743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8939 a_24236_11849# a_23837_11477# a_24110_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8940 vccd1 clkbuf_0_net57.X a_2686_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8942 _1625_.X a_13408_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8943 _1243_.Y _1243_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8944 vssd1 _1902_.Q a_7428_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8945 vccd1 a_7159_20884# _1557_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8947 _1876_.Q a_23323_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8948 a_11287_27613# a_10589_27247# a_11030_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8949 _1536_.A a_18699_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X8950 _1329_.S a_8548_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X8951 a_23282_29967# a_22843_29973# a_23197_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8952 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8954 _1325_.A2 a_5731_12567# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8956 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_8109_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8957 vssd1 _1568_.B a_10601_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X8958 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8959 a_1941_6037# a_1775_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8960 a_10951_24233# _0921_.A a_10593_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8961 a_10497_19997# a_9963_19631# a_10402_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8962 a_13517_14709# _1105_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X8963 vccd1 _1129_.B a_23759_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X8964 a_15330_22351# _1116_.D1 a_15081_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X8965 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_11711_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X8966 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8967 vccd1 a_6056_20871# _1328_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X8968 a_11969_2589# a_11435_2223# a_11874_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X8969 a_4213_24135# _1763_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X8970 _1513_.A a_20216_22467# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X8972 vccd1 a_28015_5755# a_27931_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8974 a_7277_2223# a_7111_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8975 a_2129_3855# _1796_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8976 a_16849_31599# _1859_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8977 a_2005_32375# _1337_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8978 a_25156_28335# a_24757_28335# a_25030_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X8979 vccd1 a_25623_15547# a_25539_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X8980 a_25030_2589# a_24757_2223# a_24945_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X8981 a_20591_1898# _1629_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8983 _1507_.A a_19664_23555# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8984 a_20782_4511# a_20614_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X8985 a_20487_28701# a_19623_28335# a_20230_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X8986 vccd1 _1301_.A1 a_5081_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X8987 _1060_.C1 a_9595_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X8988 vccd1 _1125_.X _1126_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8989 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9135_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X8990 vccd1 a_21831_25071# _1876_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8991 a_14195_13647# _1038_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8992 a_7619_2986# _1660_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8993 a_22879_31055# a_22181_31061# a_22622_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8994 _1099_.B1 a_18243_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X8995 a_13721_21263# _1851_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X8997 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_6808_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X8998 a_22454_31055# a_22015_31061# a_22369_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X8999 _1390_.B a_27831_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9000 a_7939_13967# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9001 a_25455_5853# a_24591_5487# a_25198_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9002 vssd1 _1887_.CLK a_24591_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9003 vssd1 _1816_.CLK a_7111_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9004 a_24209_1679# _1628_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9005 a_2897_10927# _1226_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9006 vssd1 _1486_.B a_13545_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9007 a_9772_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9008 vssd1 _2006_.Q a_9963_15939# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9009 vccd1 _2006_.Q a_10213_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X9010 a_27057_10927# a_26891_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9011 vccd1 a_10386_29941# a_10313_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9012 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9013 a_21917_21807# a_21647_22173# a_21827_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9014 _1382_.X a_15616_18115# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X9015 a_5727_17999# _1785_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9016 vssd1 a_25014_17973# a_24972_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9018 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9019 _1311_.B1 a_4899_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9020 a_20157_28701# a_19623_28335# a_20062_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9021 vssd1 _1985_.CLK a_26431_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9022 a_19878_5853# a_19439_5487# a_19793_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9023 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9024 a_2915_27613# a_2051_27247# a_2658_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9026 a_20315_25834# _1531_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9027 a_23776_17289# a_23377_16917# a_23650_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9028 a_17673_1135# a_17507_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9030 a_18685_16911# _1179_.B2 a_18601_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9031 a_11877_1135# a_11711_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9034 vssd1 _1140_.C a_14533_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9035 a_18697_28335# a_18427_28701# a_18607_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9037 _0984_.B1 a_10731_17483# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X9038 vccd1 a_22015_7119# _1924_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9039 vssd1 a_27847_3677# a_28015_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9040 _1562_.A a_12743_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9042 vssd1 a_10459_27791# a_10627_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9043 vccd1 a_15887_29789# a_16055_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9044 _0918_.A a_3983_19631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X9045 a_9961_12675# a_9687_12919# a_9879_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9046 vccd1 a_4035_30485# _1330_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X9047 vssd1 _1867_.Q a_14833_30333# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9048 vccd1 a_12042_25183# a_11969_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9049 a_11797_17455# a_11527_17821# a_11693_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9050 a_9613_16600# _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X9051 a_2585_27613# a_2051_27247# a_2490_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9052 vccd1 a_1673_22453# a_1779_22453# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9053 vssd1 a_12771_21482# _1901_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9054 _1250_.B2 _1249_.A1 a_5015_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9055 a_26870_17821# a_26431_17455# a_26785_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9056 vssd1 a_13643_3855# _1941_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9057 a_7002_4943# _1208_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X9058 a_5397_24233# _1294_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X9059 vssd1 _0958_.B a_14901_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9060 a_12245_1501# a_11711_1135# a_12150_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9061 _1332_.Y _1353_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9062 a_16661_26159# a_16495_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9063 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9066 _1151_.X a_21463_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9069 _0935_.X a_8307_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9070 a_26226_4765# a_25953_4399# a_26141_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9071 a_3041_21807# _1762_.A a_2603_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9072 vccd1 _1033_.A2 a_20157_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9073 vssd1 _0958_.B a_20421_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9074 a_23239_27791# a_22457_27797# a_23155_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9075 a_13398_25321# _1484_.B a_13316_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9078 vccd1 _0981_.B a_14043_20513# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X9079 a_1677_3087# _1221_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9080 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8556_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9081 vssd1 a_23903_19796# _1387_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9082 a_24462_1653# a_24294_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9083 vccd1 _1775_.A2 a_8120_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9084 vccd1 a_22983_19796# _1823_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9085 _0983_.B1 a_13399_17483# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9086 _1545_.A a_14467_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9087 a_3155_17455# _1323_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9088 a_2765_4233# a_1775_3861# a_2639_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9089 _0930_.Y _0930_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9090 _1722_.A a_22379_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9091 vssd1 a_23523_22173# a_23691_22075# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9092 vccd1 a_23047_25589# a_22963_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9093 a_13898_24527# a_13625_24533# a_13813_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9096 a_24757_23983# a_24591_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9098 a_16921_14709# _1091_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9099 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9101 vccd1 a_24075_23439# a_24243_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9102 a_2505_16911# _1249_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9105 vssd1 _2023_.CLK a_1591_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9106 a_23303_12381# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9107 vssd1 a_24075_23439# a_24243_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9108 a_26091_29789# a_25309_29423# a_26007_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9109 vccd1 a_27038_6687# a_26965_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9110 a_16054_7913# _1041_.C1 a_15974_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9114 a_8031_13353# _1034_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9115 _1273_.A1 a_2807_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9117 vccd1 a_23303_6031# fanout20.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9118 vccd1 _0958_.B a_20267_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9120 a_7626_4511# a_7458_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9121 vccd1 a_24547_5162# _1731_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9122 a_25125_21807# a_24959_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9123 a_9742_4511# a_9574_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9124 a_17102_26271# a_16934_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9126 vccd1 _1544_.A_N a_8399_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9127 vccd1 a_3983_3311# _1816_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9128 _1205_.Y _1177_.C a_4250_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X9131 vccd1 _1090_.C a_16711_15307# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X9132 a_7626_4511# a_7458_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9133 a_8259_10927# _2008_.Q a_7896_11079# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X9134 vccd1 a_23967_3829# a_23883_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9135 a_4774_1247# a_4606_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9136 vccd1 a_7867_3829# a_7783_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9137 _1869_.Q a_22863_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9140 a_24719_1679# a_24021_1685# a_24462_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9142 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9143 vccd1 a_23443_12778# _1979_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9144 a_2539_6941# a_1757_6575# a_2455_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9145 _0988_.X a_14319_7691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9146 a_24236_10761# a_23837_10389# a_24110_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9147 a_23009_29973# a_22843_29973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9148 vssd1 a_9247_2741# a_9205_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9149 a_4774_1247# a_4606_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9150 vssd1 _1183_.B1 a_19952_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X9151 _1056_.D1 a_13367_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9152 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9153 _1103_.A1 a_25807_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9154 vssd1 fanout21.X a_23565_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9155 vssd1 _1773_.B _1773_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9156 a_2581_1135# a_1591_1135# a_2455_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9158 vccd1 _1234_.Y _1237_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X9159 a_19310_1653# a_19142_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9160 a_8485_7485# a_8215_7119# a_8395_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9161 vccd1 _1474_.A_N a_9595_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9162 a_25589_20175# _1970_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9163 vccd1 a_10811_1653# a_10727_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9164 a_10218_6031# a_9945_6037# a_10133_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9165 vccd1 a_13517_14709# _1108_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9166 vssd1 a_2122_9839# a_2228_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9167 vssd1 _1265_.A2 a_5996_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9168 _1985_.Q a_25807_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9170 vssd1 a_9999_5853# a_10167_5755# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9171 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_3240_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9172 _1790_.Y _1273_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X9174 _1531_.A a_19619_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9175 a_19973_26525# a_19439_26159# a_19878_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9176 vssd1 a_22063_22570# _1882_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9177 a_24846_17999# a_24573_18005# a_24761_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9178 vccd1 a_1591_15279# _0929_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9179 _0952_.A1 a_19439_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9181 _0918_.A a_3983_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9182 a_2769_17231# _1277_.B a_2673_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9183 vccd1 _1304_.B a_6406_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9184 a_5632_3561# _1804_.Y _2021_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X9186 vssd1 a_27399_16042# _1701_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9187 vssd1 _0935_.X a_14103_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9188 _1873_.Q a_25623_31867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9190 a_8204_28111# _1775_.A2 _1775_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X9191 a_6705_16341# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X9193 a_13955_31055# a_13091_31061# a_13698_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9195 vccd1 a_25842_26677# a_25769_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9196 a_19133_10749# _1182_.B a_19061_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9197 a_21537_30511# a_21371_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9198 vssd1 _1006_.B2 a_27437_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9200 _1117_.B a_10627_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9201 vssd1 _1047_.C a_14625_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9202 a_13898_24527# a_13459_24533# a_13813_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9203 _1755_.A a_6831_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9204 a_10597_6825# _0988_.X a_10681_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9205 _1885_.Q a_27463_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9206 a_5047_21237# _1282_.A2 a_5265_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X9207 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9208 _0991_.X a_15607_12043# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9209 vssd1 a_13146_12533# a_13104_12937# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9210 _1182_.B a_25623_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9211 vccd1 _1829_.Q a_15479_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9212 a_13521_16367# _1840_.Q a_13449_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9215 _0925_.A2 a_10423_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9216 _1882_.Q a_27095_25339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9217 a_23289_3855# _1991_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9218 a_20004_5487# a_19605_5487# a_19878_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9219 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_6808_30761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9220 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_13367_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9221 a_5152_29673# a_4903_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9222 a_7189_3855# _1365_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9223 a_25708_29423# a_25309_29423# a_25582_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9224 vccd1 _1887_.CLK a_24591_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9225 a_14737_23805# _1053_.A a_14655_23552# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9226 a_24075_23439# a_23211_23445# a_23818_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9227 _1033_.B1 a_14379_9408# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9228 vccd1 _1374_.A_N a_8675_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9229 _1846_.Q a_12927_15547# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9230 a_4798_12265# _1216_.A2 a_4495_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X9231 a_19049_28111# _1842_.Q a_18703_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X9232 vccd1 a_2658_27359# a_2585_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9233 vssd1 _1031_.X a_17381_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X9234 a_20039_5162# _1607_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9236 _1190_.B1 a_21127_12897# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9237 a_9786_23805# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X9238 a_25815_11293# a_25033_10927# a_25731_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9239 a_8031_17999# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9241 vccd1 temp1.capload\[7\].cap.A temp1.capload\[7\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9242 a_25455_13469# a_24591_13103# a_25198_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9243 a_3707_6144# _1281_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9244 a_4064_21583# _1307_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X9246 _1084_.A1 a_12723_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X9247 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8307_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9248 a_16083_17130# _1382_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9250 vssd1 a_4035_20693# _1268_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9251 a_26597_6575# a_26431_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9252 a_16863_11177# _1155_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9253 a_27149_27247# a_26983_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9254 vccd1 _1723_.A_N a_22199_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9255 a_2143_17705# _1311_.A1 a_2225_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X9256 _0921_.A a_2971_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X9257 vssd1 a_13517_14709# _1108_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X9258 _1156_.Y _1143_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9259 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4903_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9260 a_19605_20969# _1835_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9261 a_10133_1679# _1616_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9262 a_8280_12265# _1071_.X a_8178_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X9263 _1433_.A a_10188_18115# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9264 a_7201_14851# _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9265 vccd1 a_25198_2335# a_25125_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9266 _1065_.B a_25623_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9267 vssd1 _0993_.X a_18324_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X9268 a_27859_30676# _1450_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9269 vccd1 _1344_.Y a_8215_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9270 a_2214_3677# a_1941_3311# a_2129_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9272 _1347_.Y temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9273 _1061_.X a_18795_7232# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9274 _1334_.A1 _1325_.A2 a_6843_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X9275 vccd1 _1905_.Q a_10270_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9276 a_21511_28500# _1483_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9277 a_11563_31965# a_10865_31599# a_11306_31711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9278 a_8579_4943# a_8399_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9279 a_20797_32521# a_19807_32149# a_20671_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9281 vssd1 a_27590_12127# a_27548_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9282 a_7561_22941# _0921_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9283 a_7015_22351# a_6835_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9285 vssd1 _2003_.Q a_7755_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X9286 vssd1 fanout20.X a_22935_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9287 a_21407_2589# a_20709_2223# a_21150_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9288 a_6559_24640# _1304_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9289 a_13257_13353# _1199_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X9290 _1293_.A1 a_17139_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9291 a_23615_22351# a_22917_22357# a_23358_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9292 vssd1 _1816_.CLK a_6835_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9293 a_16531_24349# a_15833_23983# a_16274_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9294 vccd1 _1723_.B a_22195_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9295 a_17999_16395# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9296 a_8381_2773# a_8215_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9297 vccd1 a_10643_8207# a_10811_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9298 a_23013_10927# _1716_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9299 vssd1 a_20471_29691# a_20429_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9300 _1081_.C1 a_21095_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9301 _1416_.A a_18423_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9302 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9303 a_14643_13647# _1050_.C a_14449_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9305 _1122_.A1 _1120_.X a_9779_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9306 a_12337_24233# _1451_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9307 _1019_.B a_21575_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9308 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_4811_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9309 a_15931_15823# _1029_.X a_15737_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9310 a_8449_17999# _1764_.A a_8031_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9313 vssd1 _1132_.C a_15969_13131# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9314 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X9316 a_5816_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9318 a_1674_28879# clkbuf_0_temp1.i_precharge_n.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9319 temp1.capload\[2\].cap.Y temp1.capload\[2\].cap_47.LO a_22745_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9320 a_20942_19203# _1405_.B a_20860_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9321 vccd1 fanout33.A a_16495_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9322 _1303_.A1 a_4443_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X9323 vccd1 _1744_.A_N a_19439_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9324 _1219_.A2 a_2696_11177# a_2897_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9325 a_15277_30511# a_14287_30511# a_15151_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9326 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7104_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9327 a_18751_21972# _1497_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9328 a_22063_18218# _1527_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9329 _1515_.A a_21412_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X9331 a_26203_10602# _1727_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9335 _1183_.B1 a_18979_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9336 _1823_.CLK a_22659_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X9337 a_18180_9295# _1112_.B1 a_18078_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X9338 a_25156_20719# a_24757_20719# a_25030_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9339 a_17473_15797# _1029_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9340 vssd1 clkbuf_0_net57.X a_1674_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9341 a_25198_27359# a_25030_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9342 _1238_.X a_7667_22901# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X9343 vccd1 a_22622_2741# a_22549_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9344 a_9301_4399# a_9135_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9345 a_7185_4399# a_7019_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9346 _1255_.A1 a_2807_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9347 vssd1 a_4863_23413# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9349 a_25674_13647# a_25235_13653# a_25589_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9350 vssd1 a_3007_1679# a_3175_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9351 a_8356_20407# _1233_.A1 a_8498_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9352 vccd1 _1887_.CLK a_25235_20181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9353 vssd1 a_6073_25045# _1344_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X9354 a_17831_30676# _1471_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9355 vccd1 a_9779_12015# _1198_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9357 vssd1 _1844_.Q a_13040_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9358 a_26927_23261# a_26229_22895# a_26670_23007# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9359 vssd1 _0981_.B a_15453_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9360 a_10727_8207# a_9945_8213# a_10643_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9361 a_1735_29941# temp1.inv2_2.Y a_2073_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X9362 vssd1 _1097_.X a_16185_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X9364 a_8038_11254# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X9365 a_12575_13647# a_11877_13653# a_12318_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9366 a_16175_1898# _1665_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9367 a_10202_22325# a_10034_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9368 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9369 a_20337_13967# _1191_.A1 a_19899_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9370 a_16366_2335# a_16198_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9373 _1116_.B1 a_17231_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9374 vssd1 _1887_.CLK a_24407_18005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9375 vccd1 _1888_.Q a_19470_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9376 a_25800_17289# a_25401_16917# a_25674_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9377 vccd1 _1121_.A1 a_5670_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9378 a_18416_17455# _1888_.Q a_17841_17601# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X9379 _1230_.B1 _1218_.B a_4877_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X9380 a_17730_4943# _0963_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9381 vccd1 _0911_.A a_5545_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X9382 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4896_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9383 a_27347_13647# a_27167_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9385 a_25401_4949# a_25235_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9386 vccd1 _0918_.A a_7635_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X9387 a_13490_24233# _1537_.B a_13408_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9388 vssd1 _1277_.B a_4989_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9390 a_10133_29967# _1450_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9391 a_26502_25437# a_26229_25071# a_26417_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9392 vccd1 a_27279_14459# a_27195_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9393 a_8105_1685# a_7939_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9394 vssd1 _1141_.C a_18545_13131# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9395 _1013_.X a_10648_12675# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9396 vccd1 a_17930_28853# a_17857_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9398 a_6645_9001# _1086_.A a_6549_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X9399 vssd1 a_5233_11445# _1796_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9400 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_1683_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9402 vssd1 _1242_.B1 _0913_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X9403 _1450_.A a_6923_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9404 a_14655_18115# _1142_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9405 a_2129_6031# _2019_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9407 a_6736_29423# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9409 a_7743_16367# _1286_.A1 _1291_.B2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X9411 _1649_.A a_7704_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9412 vccd1 _1982_.CLK a_26983_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9413 a_13599_7828# _1749_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9414 a_24945_28335# _1894_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9415 _1705_.A a_27807_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9416 vssd1 a_23691_2491# a_23649_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9417 vccd1 a_24547_31274# _1447_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9418 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5152_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9420 _1193_.X a_16127_16617# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X9421 vssd1 _0966_.A2 a_16105_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9422 a_17302_17999# a_17029_18005# a_17217_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9423 vccd1 a_25623_5755# a_25539_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9424 vssd1 _1528_.A a_20860_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9426 a_12720_16143# _0983_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X9428 vssd1 a_2807_3579# _1234_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9430 a_5136_22583# _1303_.A1 a_5278_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9432 vssd1 a_19027_25834# _1894_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9433 _1887_.CLK a_23395_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X9434 vccd1 a_11711_16919# _1422_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X9437 a_24547_31274# _1447_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9438 vccd1 _1440_.B a_14467_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9439 a_2037_13103# _1810_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9441 a_13629_1679# _1659_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9442 vccd1 a_2547_8029# a_2715_7931# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9444 a_25125_2589# a_24591_2223# a_25030_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9445 a_16290_4399# a_16113_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9446 a_2125_25071# a_1959_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9448 a_25842_24501# a_25674_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9449 a_18601_14191# _1110_.A a_18519_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9450 a_1766_26159# clkbuf_1_1__f__0380_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9452 a_17305_29423# a_17139_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9453 a_23013_4943# _1929_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9454 vccd1 a_22707_9514# _1926_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9455 vccd1 a_15081_22325# _1116_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9456 a_18887_20175# _1184_.B1 a_19065_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9458 vccd1 _1999_.CLK a_9779_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9459 vccd1 _1895_.Q a_15882_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9460 a_19027_25834# _1534_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9461 vccd1 a_7111_25071# _1242_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9462 a_15432_1385# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9463 a_9227_17705# _1764_.A a_9477_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9464 vssd1 _1721_.B a_22469_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9465 a_20617_11471# a_20083_11477# a_20522_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9466 a_11023_31274# _1479_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9468 a_2198_1247# a_2030_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9470 a_7515_1501# a_6817_1135# a_7258_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9471 vccd1 a_19567_1679# a_19735_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9472 a_26099_6031# a_25235_6037# a_25842_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9473 a_1673_16911# _1277_.B _1323_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9474 a_17727_29967# a_16863_29973# a_17470_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9475 vssd1 _1303_.X a_5449_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X9476 a_27215_4074# _1366_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9479 a_1860_31375# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9480 a_25674_24527# a_25401_24533# a_25589_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9481 a_16301_22057# _1898_.Q a_16219_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9482 a_25842_20149# a_25674_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9483 a_12219_23478# _1306_.A2 a_11760_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X9484 a_14852_16367# a_14453_16367# a_14726_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9485 vccd1 _1873_.CLK a_24591_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9486 a_16911_5162# _1633_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9487 a_15457_6005# _0993_.X a_15614_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X9488 a_2382_6005# a_2214_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9489 vssd1 a_2382_7093# a_2340_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9491 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9492 a_27038_17567# a_26870_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9493 a_26670_25183# a_26502_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9495 _1723_.A_N a_22015_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X9496 vssd1 _1876_.CLK a_25143_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9497 a_19619_3677# a_19439_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9498 vccd1 a_26394_4511# a_26321_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9499 vccd1 _1153_.A a_21279_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9500 vccd1 _1744_.A_N a_19623_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9501 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9135_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9502 vssd1 a_1829_16341# _1311_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X9503 a_17397_29967# a_16863_29973# a_17302_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9504 a_3042_24527# a_2603_24533# a_2957_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9505 a_19836_15823# _1024_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X9507 _0921_.Y _0921_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9508 a_17497_14013# _1127_.A a_17415_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9509 vccd1 a_2547_13469# a_2715_13371# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9510 vccd1 _1342_.B a_4719_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9512 a_2455_8207# a_1591_8213# a_2198_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9513 a_18584_31849# a_18335_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9515 a_6921_26159# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9517 _1142_.B1 a_10055_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9518 a_5817_5487# _1317_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9519 a_19786_31055# a_19513_31061# a_19701_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9521 vccd1 _2005_.Q a_11693_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X9522 a_7803_20884# _1445_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9523 a_24639_14356# _1722_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9524 a_25398_22173# a_25125_21807# a_25313_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9525 a_23523_3677# a_22659_3311# a_23266_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9526 a_15549_20291# _1181_.X a_15477_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9527 a_25589_12559# _1965_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9528 vccd1 a_11711_27791# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9529 vssd1 a_22143_26525# a_22311_26427# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9530 a_27167_13647# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9531 a_20897_22895# _1829_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9532 a_22806_20149# a_22638_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9533 a_16986_3971# _1607_.B a_16904_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9535 _1066_.B a_23047_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9536 a_9742_5599# a_9574_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9537 a_21218_11177# _1577_.B a_21136_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9538 vccd1 _1881_.Q a_20390_21379# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9539 _1090_.C a_9282_16341# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X9540 vccd1 a_15633_11445# _1120_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9541 vccd1 a_9963_15939# _0987_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X9542 a_14986_3829# a_14818_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9543 _1134_.B1 a_15483_23552# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9544 vccd1 _0918_.A a_7821_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X9545 _1095_.B1 a_11711_12672# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9546 vccd1 a_22247_20884# _1879_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9547 _1105_.X a_17231_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9548 vssd1 _1144_.B a_6829_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9549 a_11306_31711# a_11138_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9551 a_9949_27791# _1818_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9552 vssd1 a_24811_14735# a_24979_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9553 a_9016_27791# a_8767_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X9554 _1230_.B1 _1217_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.08775 ps=0.92 w=0.65 l=0.15
X9555 a_24757_13103# a_24591_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9556 a_22469_14191# a_22199_14557# a_22379_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9558 vssd1 a_6303_2491# a_6261_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9559 _1177_.C a_7295_6031# a_7828_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9560 a_6463_14441# _1780_.B1 a_6245_14165# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9561 a_17573_4917# _0997_.X a_17730_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X9562 a_22638_20175# a_22365_20181# a_22553_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9563 vssd1 a_7387_15823# _1775_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9564 vccd1 a_5878_2335# a_5805_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9565 a_25221_10927# _1680_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9566 vccd1 a_17473_15797# _1029_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X9567 a_22837_9839# a_22567_10205# a_22747_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9568 a_14345_24129# _1056_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9569 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9572 a_22247_20884# _1502_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9573 a_20942_19881# _1506_.B a_20860_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9574 a_9275_10602# _1560_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9575 a_27663_15645# a_26965_15279# a_27406_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9576 a_18114_32117# a_17946_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9578 a_11902_24566# _1287_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X9579 vssd1 _1329_.S a_5392_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9580 _1366_.X a_4760_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9581 _1133_.X a_17415_24640# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9582 vccd1 a_12743_13621# a_12659_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9584 vssd1 _1329_.S a_4263_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X9585 vccd1 _1882_.Q a_20850_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9586 _1101_.X a_13275_17024# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9587 _1205_.Y _1170_.B1 a_4466_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
X9588 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9589 vssd1 a_14307_1653# a_14265_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9590 _1136_.B a_25531_9269# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9591 vssd1 _0958_.A _1086_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9592 a_7258_1247# a_7090_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9593 a_10125_31433# a_9135_31061# a_9999_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9595 a_17381_7093# _1061_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X9597 vccd1 _1830_.CLK a_22935_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X9598 a_14901_12015# _1025_.B a_14829_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X9599 a_25674_24527# a_25235_24533# a_25589_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9600 a_16208_19407# _1972_.Q a_15633_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X9601 vssd1 _1246_.B2 _1216_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9602 vccd1 a_10386_6005# a_10313_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9603 _1049_.C1 a_14287_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9604 a_23023_21085# a_22843_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9605 a_11803_18909# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9606 vssd1 a_18850_3829# a_18808_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9607 a_11403_16367# _2006_.Q a_11312_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X9608 a_7649_15279# a_7472_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9611 a_17691_21376# _1886_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9612 a_12299_20495# _0956_.C a_12199_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X9613 a_4035_10901# _1226_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X9615 a_20315_26922# _1536_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9616 vccd1 a_2472_15431# _1249_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9617 _1441_.A a_14467_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9618 a_13846_14735# _1108_.C1 a_13766_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9619 a_18151_10496# _1080_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9620 a_4220_21959# _1294_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X9622 a_1591_20719# _1283_.B1 a_1769_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9623 a_11877_1135# a_11711_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9624 vssd1 a_22162_31711# a_22120_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9625 _1177_.Y _1175_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X9626 a_13054_25589# a_12886_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9627 a_22983_21482# _1515_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9629 vccd1 _1132_.A a_18887_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9630 vccd1 _1195_.B2 a_20539_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X9631 a_9999_4765# a_9135_4399# a_9742_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9632 a_5817_19087# _1325_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X9633 a_20591_7338# _1747_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9634 a_23098_22173# a_22659_21807# a_23013_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9635 vssd1 _1121_.A1 a_9779_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9636 a_1643_21237# _1259_.X a_2009_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9638 _1560_.X a_9591_11293# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9639 vssd1 _1873_.CLK a_21831_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9640 _1359_.X a_8395_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9641 vssd1 a_16311_18543# fanout37.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9643 a_21997_29423# a_21831_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9644 a_15387_1679# a_15207_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9645 a_22346_6687# a_22178_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9646 a_19786_31055# a_19347_31061# a_19701_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9647 a_10270_18115# _1422_.B a_10188_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9648 a_18607_28701# a_18427_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9649 a_20046_26271# a_19878_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9650 vssd1 a_17473_15797# _1029_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X9651 vccd1 _1246_.B1 a_2103_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X9653 _1895_.Q a_24979_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9654 vccd1 _1914_.Q a_20758_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9655 a_22546_6031# a_22369_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9656 a_22346_6687# a_22178_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9657 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9658 a_27406_21919# a_27238_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9659 a_26321_4765# a_25787_4399# a_26226_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9660 vssd1 a_2327_5487# _1532_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9661 _1118_.X a_17139_11584# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9662 vssd1 a_23450_29941# a_23408_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9664 vccd1 a_23783_22325# a_23699_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9665 vccd1 _1075_.C a_17691_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9666 a_7050_25731# _1422_.B a_6968_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9669 a_2686_15823# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X9670 vccd1 _1090_.C a_18151_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9672 vssd1 a_26651_4765# a_26819_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9673 _1084_.B1 a_9176_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9674 vccd1 a_5261_10973# a_5361_11191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9677 vssd1 _1133_.C a_19557_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9679 _1232_.Y _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X9680 a_2723_4765# a_1941_4399# a_2639_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9681 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9682 vccd1 _1875_.Q a_15512_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X9683 vccd1 _1823_.CLK a_26431_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9684 a_26413_14191# a_26247_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9685 a_7203_29967# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9686 vccd1 a_2382_3423# a_2309_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9687 a_7939_13647# _1012_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9688 a_22638_20175# a_22199_20181# a_22553_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9689 _1324_.A _1052_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9690 a_25743_1898# _1654_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9691 vccd1 _1316_.X a_5087_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9692 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_18584_31849# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9693 vccd1 a_27847_26525# a_28015_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9694 _1322_.A a_5547_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9695 a_25198_24095# a_25030_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9696 a_11869_17455# _0956_.C a_11797_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X9697 vssd1 _1860_.CLK a_9963_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9698 vccd1 a_9460_25847# _1337_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X9699 a_15656_22671# _1875_.Q a_15081_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X9700 a_27590_19743# a_27422_19997# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9701 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9703 _1021_.A a_15299_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X9705 a_5203_24233# _1294_.B2 a_5397_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X9706 a_15565_23805# _1132_.A a_15483_23552# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9708 vccd1 _1639_.X a_12171_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9710 vssd1 a_27847_19997# a_28015_19899# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9711 _1711_.X a_23299_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9712 a_7718_2335# a_7550_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9713 vssd1 a_21978_30623# a_21936_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9714 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9715 a_22238_14735# _1979_.Q a_22081_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X9716 _1191_.X a_19899_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X9717 a_25750_9951# a_25582_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9719 a_18519_26703# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9720 vccd1 _1374_.A_N a_22015_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9721 vccd1 _1685_.A_N a_20819_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9722 vssd1 _1135_.B a_20537_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9723 _1317_.X a_5087_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X9724 vssd1 _1860_.CLK a_9135_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9725 a_18969_19453# _1132_.A a_18887_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9726 vssd1 _1246_.A3 a_3247_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.219375 pd=1.325 as=0.10075 ps=0.96 w=0.65 l=0.15
X9727 vccd1 a_16991_9117# a_17159_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9728 a_15750_28335# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X9729 vccd1 a_4587_24501# _1767_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X9730 a_14379_20719# _1858_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X9731 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9732 a_13441_1685# a_13275_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9733 vssd1 _1207_.B1_N _1226_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9734 vssd1 a_2547_8029# a_2715_7931# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9735 vssd1 _1269_.A1 a_8919_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9736 a_19142_14735# a_18703_14741# a_19057_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X9737 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X9738 vssd1 a_24639_4564# _1959_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9739 vccd1 _1851_.Q a_9258_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X9740 a_10397_14735# _1269_.A1 a_10147_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9741 a_5805_2589# a_5271_2223# a_5710_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9743 vssd1 a_27095_25339# a_27053_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9744 vssd1 a_10570_19743# a_10528_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9745 a_3133_18319# _1281_.A1 a_2695_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9746 _1202_.Y _1170_.A3 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9747 a_15277_9839# a_14287_9839# a_15151_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9748 a_22419_31965# a_21555_31599# a_22162_31711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9749 a_7847_19997# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9750 vccd1 a_2932_18517# _1302_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X9751 _1376_.X a_11983_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9753 a_22603_5853# a_21739_5487# a_22346_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X9754 a_17250_14735# _1091_.C1 a_17170_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9755 a_22622_25589# a_22454_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9756 vccd1 _1775_.C1 a_1591_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9757 a_5731_24847# _1308_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9759 vssd1 _1804_.Y a_5541_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X9760 vccd1 _0921_.B _1232_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9761 a_14373_6397# a_14103_6031# a_14283_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9762 _1568_.B a_11455_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9763 a_19268_18377# a_18869_18005# a_19142_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X9764 a_23742_4399# a_23565_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9765 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_3983_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9766 vssd1 _1775_.C1 _1767_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9767 a_1841_22057# _1775_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9768 a_2047_16617# _1230_.A4 a_1829_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9769 vccd1 _0964_.A a_13551_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9770 _1194_.B2 a_13663_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9772 a_18090_17705# _1048_.X a_17841_17601# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X9773 a_11760_24759# _1306_.A2 a_11902_24566# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X9774 a_10313_6031# a_9779_6037# a_10218_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9775 vssd1 _0987_.Y a_12149_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X9777 a_22089_31965# a_21555_31599# a_21994_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9778 a_17113_6005# _0997_.X a_17270_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X9779 _1832_.Q a_23323_24251# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9780 a_3514_25615# _1761_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9781 a_22454_25615# a_22181_25621# a_22369_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9782 a_10007_23805# _0911_.A a_9644_23671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X9783 vccd1 a_9284_21781# _1282_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X9785 a_20249_27797# a_20083_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9786 _1023_.B a_24703_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9787 a_12065_11471# _1847_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9788 a_15299_20291# _1186_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9790 vssd1 a_25842_23413# a_25800_23817# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9791 vssd1 _1982_.CLK a_23303_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X9792 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_5639_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X9794 vssd1 _1289_.A2 a_4209_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X9795 vssd1 a_19487_11690# _1586_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9797 _1577_.X a_20676_12265# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9798 a_7428_24233# _1537_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9799 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_11711_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X9801 _1781_.B _0911_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9802 a_26133_3311# a_25143_3311# a_26007_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9803 a_5081_15279# _1250_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9804 a_4036_14165# _1325_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X9807 vccd1 a_16911_5162# _1942_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9809 a_22843_21085# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9810 a_19487_11690# _1586_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9811 _1408_.A a_18560_23145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9812 _1855_.Q a_11731_31867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9815 a_14465_8527# _1440_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X9816 a_20885_16341# _1293_.A1 a_21138_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X9817 a_1591_24527# _1771_.B _2007_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9818 a_9921_16911# _1269_.A1 a_9503_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9820 a_4669_9839# _1324_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X9821 a_23523_3677# a_22825_3311# a_23266_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9822 a_18114_1247# a_17946_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9823 vccd1 _1763_.A2 a_4547_24305# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X9826 a_24757_15823# a_24223_15829# a_24662_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X9827 vssd1 a_14335_2388# _1935_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9830 a_11789_25071# _1852_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9832 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_9772_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X9834 a_18114_1247# a_17946_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9835 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_5271_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9836 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9837 a_26597_6575# a_26431_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9839 vccd1 clkbuf_0_net57.A a_2594_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9840 a_22185_29423# _1869_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9842 vssd1 _0983_.A2 a_12896_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X9843 vssd1 a_11693_17821# _1113_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X9844 a_12337_19453# _0956_.C a_12237_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X9845 vssd1 _1132_.C a_15637_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9846 _1126_.Y _1298_.A1 a_6997_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9847 _1762_.Y _1764_.B a_5639_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9849 a_27406_15391# a_27238_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9851 a_1828_19061# _1764_.A a_2048_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9853 vssd1 a_13599_29588# _1469_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9854 a_19981_13647# _1190_.X a_19899_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9856 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9857 _1975_.Q a_25623_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9858 vccd1 _1924_.CLK a_24591_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9859 a_15381_8751# _0939_.A a_15299_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9860 a_12723_10089# _1069_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9861 vssd1 _1046_.B a_23389_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9862 a_7005_1135# _1755_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9863 a_12701_8585# a_11711_8213# a_12575_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X9866 vssd1 _1074_.C a_13521_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9867 vssd1 _1226_.B1 a_2897_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9868 a_20529_4399# _1941_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9869 a_14839_10499# _1008_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9870 a_20999_4943# a_20819_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9871 _1553_.A a_7428_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9872 a_15410_22351# _1116_.C1 a_15330_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9873 vssd1 _1834_.Q a_19388_22467# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9874 a_14379_18793# _1082_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9875 _1715_.X a_27347_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9876 vccd1 _0981_.B a_14747_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X9877 vccd1 fanout28.A a_2235_2775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X9878 a_7564_29423# _1347_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X9879 a_20081_12559# _1293_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9880 a_5145_23759# _1242_.B1 a_5061_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X9881 _1445_.A a_9176_19881# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X9882 vccd1 a_26267_6005# a_26183_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9883 a_21235_25236# _1511_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9885 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5980_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X9886 vssd1 a_8785_20473# a_8719_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X9887 vccd1 _1941_.CLK a_22015_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9888 a_17270_6031# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X9889 a_19286_28995# _1484_.B a_19204_28995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9890 a_2686_26703# clkbuf_0_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9891 a_13120_6825# _0988_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X9892 a_2658_27359# a_2490_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X9893 a_19793_5487# _1942_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X9894 vssd1 _1103_.A1 a_20629_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9896 vccd1 a_8818_11703# _1124_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X9897 _1095_.C1 a_17967_12672# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9898 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X9899 a_19619_23261# a_19439_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X9900 _0974_.A2 a_28015_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9902 vccd1 a_17102_26271# a_17029_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X9903 vssd1 _1058_.B a_6645_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X9904 vssd1 a_23691_27515# a_23649_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9905 vccd1 a_4059_15431# _1278_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X9907 a_26785_23983# _1885_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X9908 a_9643_23222# _1305_.B a_9184_23047# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X9909 a_9613_22869# _0913_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X9911 _1038_.C1 a_16495_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X9912 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X9913 a_8723_4074# _1566_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X9914 _1723_.B a_27279_14459# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9915 a_24619_10383# a_23837_10389# a_24535_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9916 vccd1 a_15795_31055# a_15963_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9917 vccd1 _1941_.CLK a_15759_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9918 vssd1 fanout33.A a_16495_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X9919 vccd1 a_7479_24527# _1242_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X9920 _0925_.Y _0922_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X9921 vccd1 a_2623_8181# a_2539_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9922 a_27031_29588# _1352_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X9923 vssd1 _1075_.C a_21213_12897# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9924 a_22244_15055# _1032_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X9925 _1744_.X a_19803_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X9926 a_2291_29967# _1775_.B1 a_1975_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X9927 vccd1 a_16382_25071# a_16488_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X9928 vssd1 _1133_.C a_17569_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X9929 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9930 a_5048_14165# _1217_.B1 a_5177_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9931 vssd1 a_15795_31055# a_15963_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9932 vssd1 a_2235_2775# _1850_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9933 a_19439_23261# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9934 vccd1 a_2623_9269# _0911_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9935 a_14043_20513# _1053_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X9936 a_14453_16367# a_14287_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9938 _0983_.A2 a_14043_20513# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X9940 vccd1 a_23691_3579# a_23607_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X9941 a_2897_10927# _1226_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X9942 vssd1 a_25623_28603# a_25581_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9943 a_4517_17999# _1267_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9944 vssd1 _1243_.A a_6829_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X9945 vssd1 a_23323_27765# a_23281_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9946 vccd1 a_18107_14954# _1914_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9947 vssd1 a_14986_4917# a_14944_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9948 vssd1 a_18751_21972# _1877_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9949 _1699_.A a_23023_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X9950 a_18869_14741# a_18703_14741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9951 _1496_.A a_19480_25321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X9953 vccd1 _1249_.A1 a_2505_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9954 _0994_.A2 a_19275_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9955 vssd1 _1562_.A a_7980_9411# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X9956 vssd1 a_26267_24501# a_26225_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9957 vssd1 a_5565_22649# a_5499_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X9959 a_23389_14013# a_23119_13647# a_23299_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X9960 vccd1 a_2639_4765# a_2807_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9961 vccd1 a_20395_30877# a_20563_30779# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X9962 a_9889_25913# _1329_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X9963 a_2382_7093# a_2214_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X9964 a_15962_11471# _1119_.C1 a_15882_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9965 vssd1 _0997_.X a_15656_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X9966 a_18325_14013# _1110_.A a_18243_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9967 vccd1 _0909_.C a_3801_28981# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X9968 a_25582_3677# a_25309_3311# a_25497_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9970 vccd1 _2006_.Q a_9894_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9971 vssd1 _1310_.Y a_4064_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9972 a_15825_19881# _0966_.X a_15753_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9974 vccd1 a_23075_11690# _1680_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9975 vssd1 a_15163_2388# _1643_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X9976 a_8807_17999# a_9195_17973# _1074_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9978 a_14686_27497# _1484_.B a_14604_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9979 _1772_.A0 _2008_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9980 a_2309_1685# a_2143_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R17 temp1.capload\[14\].cap_44.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X9981 a_4601_6825# _1159_.X a_4529_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X9982 vccd1 a_12978_27791# a_13084_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X9984 a_5625_20541# _0911_.A a_5537_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X9985 a_2962_14735# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9987 vssd1 a_25842_4917# a_25800_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X9988 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9989 vccd1 _1474_.A_N a_10239_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9990 a_19889_16911# _1179_.B1 a_19973_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9993 vccd1 a_11023_18218# _1820_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9994 vccd1 _1744_.A_N a_20359_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X9995 a_17802_15823# _1027_.X a_17722_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X9996 _1721_.B a_27739_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9997 a_23523_11293# a_22825_10927# a_23266_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X9999 a_21127_12897# _1153_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10000 vccd1 a_7571_20175# _0956_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10001 a_16711_15307# _1021_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10002 vssd1 _2023_.CLK a_1775_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10003 vssd1 _1191_.A1 a_21136_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10005 a_2915_24349# a_2217_23983# a_2658_24095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10006 a_4613_3916# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10007 a_19893_7485# a_19623_7119# a_19803_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10009 a_10740_25731# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10010 a_22063_8426# _1580_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10011 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10012 a_19671_25834# _1496_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10013 vssd1 _1257_.X a_1828_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X10014 _1301_.A1 _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10015 a_25382_3829# a_25214_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10016 vccd1 a_16035_7119# _1590_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10018 a_18642_23145# _1405_.B a_18560_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10019 vssd1 a_12189_23737# a_12123_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10021 a_12061_4949# a_11895_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10022 a_20437_11471# _1573_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10023 vssd1 a_20471_31867# a_20429_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10024 a_25455_9117# a_24757_8751# a_25198_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10026 a_27571_9117# a_26873_8751# a_27314_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10027 vccd1 _1544_.A_N a_18427_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X10028 _1046_.B a_28015_12283# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10029 vccd1 _1897_.Q a_13490_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10030 vssd1 _1234_.A2 a_3133_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X10031 a_14369_13353# _1120_.D a_14287_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X10032 a_22015_4765# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10033 _1192_.A2 a_15411_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10034 a_10083_5853# a_9301_5487# a_9999_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10035 vccd1 a_3111_5652# _0916_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10037 a_25382_16479# a_25214_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10038 a_23443_31764# _1474_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10039 _1021_.X a_17691_22464# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10041 vssd1 _1801_.B a_4155_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X10042 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4075_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10043 vssd1 a_25639_16733# a_25807_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10044 a_4521_1135# _1367_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10045 a_10331_9295# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10046 vssd1 a_12042_2335# a_12000_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10047 vssd1 _1900_.Q a_9313_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10048 _0929_.A a_1591_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X10049 a_9233_11471# _1198_.A2 a_8818_11703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X10050 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10051 vssd1 a_21327_1300# _1990_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10052 vssd1 a_10386_6005# a_10344_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10053 _1474_.X a_13455_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10054 _1464_.X a_9775_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10055 vssd1 _1895_.Q a_15800_26819# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10058 a_18597_3855# _1935_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10059 vssd1 a_25198_13215# a_25156_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10060 vssd1 _1034_.D _1034_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10061 a_25559_10602# _1720_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10062 vssd1 _1316_.X a_7189_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10063 a_15370_32143# a_14931_32149# a_15285_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10064 vccd1 a_16182_3423# a_16109_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10067 vccd1 a_9999_7119# a_10167_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10068 a_17853_28169# a_16863_27797# a_17727_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10069 a_18519_21376# _1894_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10071 vccd1 a_20223_8426# _1582_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10072 a_26686_14557# a_26413_14191# a_26601_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10073 a_18550_5737# _1607_.B a_18468_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10074 _1056_.B1 a_14655_23552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10075 vssd1 _1845_.Q a_10188_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10076 a_20690_28853# a_20522_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10077 a_27847_3677# a_26983_3311# a_27590_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10078 vccd1 _1226_.A1 a_4338_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X10079 a_12502_15391# a_12334_15645# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10080 _1283_.B1 a_2695_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X10081 a_18673_14191# _1696_.B a_18601_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10082 a_11343_8751# _1042_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10083 a_23351_32362# _1477_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10086 a_6645_10089# _1086_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X10087 a_7515_1501# a_6651_1135# a_7258_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10088 vssd1 a_12759_15645# a_12927_15547# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10089 vssd1 a_23671_15279# _1690_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10090 a_12689_6721# _1068_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X10092 vssd1 _1291_.A1 a_5639_10089# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10093 vssd1 _2006_.Q a_12323_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10094 vccd1 fanout28.A a_15115_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X10095 a_8215_8751# _1198_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X10096 vssd1 a_9275_10602# _1561_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10097 vssd1 a_5693_19605# _1780_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10098 vssd1 a_7531_9813# _1159_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10099 a_5060_31055# a_4811_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10100 a_7786_3561# _1448_.A a_7704_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10101 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10102 temp1.capload\[7\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10103 a_5545_22057# _0913_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X10104 vccd1 _1277_.A a_1673_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X10105 a_25382_3829# a_25214_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10106 vssd1 a_8447_6740# _1812_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10107 vssd1 _1057_.B a_18560_8323# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10108 _1390_.B a_27831_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10109 vssd1 a_16083_14954# _1831_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10110 vccd1 _1436_.B a_10971_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10111 _1219_.A2 a_2696_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X10112 vssd1 _1140_.C a_12381_20747# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X10113 vssd1 _1140_.C a_11865_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10114 vccd1 _0981_.B a_16159_9867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10115 vccd1 _1159_.X a_5629_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10116 a_6736_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10117 a_17029_26525# a_16495_26159# a_16934_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10118 vssd1 a_19952_12533# _1184_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X10119 vssd1 a_10167_31029# a_10125_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10120 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5888_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10122 vccd1 _1053_.A a_10883_21271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X10123 a_24846_17999# a_24407_18005# a_24761_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10124 vccd1 _1112_.A1 a_18180_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10125 a_1841_23439# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10126 a_24761_2767# _1992_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10128 a_15243_3855# a_14379_3861# a_14986_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10129 vccd1 a_7803_6740# _1753_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10130 _1326_.A2 _1323_.A2 a_3237_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X10131 vccd1 _0994_.A2 a_15514_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10132 a_20864_15055# _1113_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X10133 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11868_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10134 vssd1 _1762_.A _0981_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10135 a_17569_14013# _1023_.B a_17497_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10136 a_12701_1135# a_11711_1135# a_12575_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10138 a_22015_19087# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10139 vssd1 io_in[0] a_2962_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10140 a_20539_6941# a_20359_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10141 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X10142 a_27973_26159# a_26983_26159# a_27847_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10144 vssd1 a_3083_27515# a_3041_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10145 a_6555_6941# a_6375_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10147 a_10777_3311# _1567_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10148 vssd1 a_2623_2491# a_2581_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10149 vssd1 _1067_.B a_7289_2045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10150 a_9313_21629# a_9043_21263# a_9223_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10152 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10153 vssd1 _1255_.A1 _1800_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10154 vccd1 a_22771_5755# a_22687_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10155 a_5520_27497# a_5271_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10156 a_23607_27613# a_22825_27247# a_23523_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10157 a_8522_24643# _1537_.B a_8440_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10158 vssd1 _1272_.B1 a_1643_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X10159 _1032_.X a_18887_19200# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10160 vccd1 _1562_.A a_8062_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10162 vssd1 a_6703_26133# _1306_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10163 a_9460_25847# _1336_.A1 a_9602_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X10164 a_14467_23261# a_14287_23261# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10165 a_19480_17705# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10166 a_21376_16367# _1024_.A2 a_20885_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X10167 a_14449_13647# _1050_.C a_14643_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10168 _1149_.A1 a_23047_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10169 a_13545_32509# a_13275_32143# a_13455_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10170 _1329_.X a_2103_31573# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10171 a_5157_1135# a_4167_1135# a_5031_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10173 vccd1 _1158_.X _1279_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10175 vccd1 a_27831_20987# a_27747_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10177 vccd1 fanout24.A a_26983_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10178 a_2685_22057# _1270_.A a_2603_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10179 vssd1 a_14986_3829# a_14944_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10180 vccd1 _0989_.A2 a_3830_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10181 vccd1 _2023_.CLK a_1775_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10182 a_11842_10089# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X10183 a_11299_12180# _1434_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10184 vssd1 a_26099_4943# a_26267_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10185 vssd1 _1982_.CLK a_22369_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10186 a_12057_21583# _1856_.Q a_11711_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X10187 vssd1 a_10021_9985# _1012_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X10188 a_12150_29789# a_11877_29423# a_12065_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10189 a_21463_18543# _1879_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10191 vccd1 a_2639_3677# a_2807_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10192 a_2382_6005# a_2214_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10193 vssd1 a_3983_17455# _0921_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10194 vccd1 _1819_.Q a_11983_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10195 vccd1 _1823_.CLK a_23211_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10196 _1902_.Q a_12743_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10198 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10199 a_19310_1653# a_19142_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10200 clkbuf_0_temp1.i_precharge_n.A a_25695_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10201 a_12978_12559# a_12705_12565# a_12893_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10203 vccd1 _1113_.C a_19439_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10204 a_24236_21641# a_23837_21269# a_24110_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10205 _1558_.X a_10188_14441# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10206 vccd1 a_15531_15444# _1399_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10207 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10208 a_25401_26709# a_25235_26709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10209 a_10133_29967# _1450_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10210 a_24757_17455# a_24591_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10211 vssd1 a_8454_15797# _1047_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10214 vccd1 a_24075_16911# a_24243_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10215 a_23013_3311# _1989_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10216 a_23155_18909# a_22457_18543# a_22898_18655# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10217 a_2723_3855# a_1941_3861# a_2639_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10218 vssd1 a_4571_7119# a_4739_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10220 vccd1 _1970_.Q a_21032_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10221 a_4877_13967# _1218_.B _1230_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10222 vssd1 a_4036_14165# _1281_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X10223 vccd1 _1089_.B a_17319_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10224 _1850_.CLK a_2235_2775# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10225 vssd1 _1139_.C a_14901_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10226 vssd1 _1853_.Q a_7013_28157# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10227 _1883_.Q a_26267_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10229 vccd1 _0921_.A a_9963_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X10230 vccd1 a_13599_13866# _1755_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10232 a_9460_15431# _1199_.A1 a_9602_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X10233 vccd1 a_18151_6031# _1744_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10234 vccd1 _1448_.A a_8307_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X10235 _1119_.C1 a_11803_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10237 vccd1 _1032_.C a_21463_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10238 _1527_.A a_19480_17705# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10239 a_23098_2589# a_22659_2223# a_23013_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10240 vssd1 _1136_.B a_22653_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10241 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_12801_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10242 a_15005_26409# _1896_.Q a_14921_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10243 a_25497_26159# _1881_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10244 vssd1 a_26175_3579# a_26133_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10245 a_2309_4765# a_1775_4399# a_2214_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10248 _1782_.X a_1816_11587# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10250 vssd1 _0921_.B a_9284_21781# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10252 a_15370_25615# a_14931_25621# a_15285_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10254 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X10256 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X10257 vssd1 a_2639_4765# a_2807_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R18 temp1.capload\[11\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10258 vssd1 a_23047_25589# a_23005_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10259 vssd1 _1823_.CLK a_26431_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10260 _1744_.B a_25623_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10261 vccd1 a_2455_1501# a_2623_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10262 a_20359_3677# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10263 a_19567_1679# a_18869_1685# a_19310_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10264 vccd1 _0930_.A _1164_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X10265 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10267 a_14931_27791# _0965_.B1 a_15013_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10268 vccd1 _1879_.Q a_21827_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10269 a_2907_25437# a_2125_25071# a_2823_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10270 a_25489_9673# a_24499_9301# a_25363_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10271 a_25309_29423# a_25143_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10272 a_19405_15797# _1127_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X10273 vssd1 _1149_.A1 a_18329_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10274 vccd1 _1845_.Q a_10270_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10275 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_5060_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10276 _1422_.B a_11711_16919# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X10277 a_10195_13268# _1558_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10278 _1246_.B1 _1222_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10279 _1456_.A a_6968_25731# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10282 a_4655_7119# a_3873_7125# a_4571_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10283 vccd1 _0921_.A a_9871_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10284 _1985_.Q a_25807_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
D3 vssd1 _1367_.X sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X10286 a_14818_3855# a_14379_3861# a_14733_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10288 vccd1 a_21115_28853# a_21031_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10289 vccd1 a_18291_2388# _1628_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10290 a_25455_24349# a_24591_23983# a_25198_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10291 vssd1 a_25623_20987# a_25581_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10292 a_27406_20831# a_27238_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10294 a_3281_20175# _1257_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10295 _1074_.C _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10296 vccd1 _1217_.A2 a_4709_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X10297 a_23607_2589# a_22825_2223# a_23523_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10298 vssd1 a_24547_5162# _1731_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10299 vssd1 _1308_.B a_4598_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
X10300 a_9477_17705# _1764_.A a_9227_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10301 _0985_.A a_19807_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10302 vccd1 _1057_.B a_18642_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10304 a_19697_30511# a_19531_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10306 vssd1 a_27463_13371# a_27421_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10307 _1011_.A1 a_10811_6005# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10308 vccd1 _1813_.Q a_8855_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10311 a_9742_31029# a_9574_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10312 a_1841_22057# _1308_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10313 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10314 _1617_.X a_11707_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10315 _1477_.A a_12535_32143# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10319 a_13018_6825# _1068_.C1 a_12938_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10320 a_7896_11079# _1124_.X a_8038_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X10321 a_3168_28169# a_2769_27797# a_3042_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10322 vssd1 a_15319_10107# a_15277_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10324 a_12355_1679# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10325 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A _0913_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10326 a_12978_12559# a_12539_12565# a_12893_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10327 vccd1 a_14345_24129# _1056_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X10328 _1438_.B a_13203_10357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10329 a_1775_10496# _1177_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10331 a_10137_21629# _1132_.A a_10055_21376# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10332 a_5635_18793# _1234_.A2 a_5417_18517# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X10333 a_8392_29423# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10334 vssd1 a_14287_29423# _1841_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10335 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_5520_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10336 _1846_.Q a_12927_15547# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10337 a_15637_23805# _1867_.Q a_15565_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10338 vssd1 a_8356_20407# _1233_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X10341 a_25773_18543# _1971_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10342 vccd1 a_6283_4399# _1999_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10343 vssd1 _1982_.CLK a_25787_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10344 vssd1 a_22983_19796# _1823_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10345 a_14557_18793# _1077_.X a_14461_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10346 a_22653_12015# a_22383_12381# a_22563_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10347 a_9574_31055# a_9301_31061# a_9489_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10348 vssd1 a_19954_31029# a_19912_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10350 a_24075_16911# a_23211_16917# a_23818_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10352 _1135_.B a_26175_10107# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10353 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10354 a_23013_21807# _1889_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10355 _1693_.A a_23667_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10356 _1568_.B a_11455_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10357 a_27881_28335# a_26891_28335# a_27755_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10358 a_27421_6575# a_26431_6575# a_27295_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10359 a_11793_21263# _1904_.Q a_11711_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10360 a_4533_18543# _1326_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X10361 _1734_.X a_21459_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10362 fanout20.X a_23303_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X10363 vccd1 a_13551_8215# _1010_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10364 a_26183_26703# a_25401_26709# a_26099_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10366 a_8654_2767# a_8381_2773# a_8569_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10367 vccd1 _1685_.A_N a_18059_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X10368 a_5451_11471# _1780_.B1 a_5233_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X10369 a_16274_24095# a_16106_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10370 vssd1 _1882_.CLK a_22751_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10371 vssd1 a_22799_7338# _1920_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10372 _1099_.D1 a_17323_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10373 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_11711_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X10375 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10377 a_22622_1653# a_22454_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10378 a_27563_16733# a_26781_16367# a_27479_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10379 vccd1 a_25750_3423# a_25677_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10381 a_10452_10089# _0987_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X10382 a_22063_29098# _1490_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10383 _1247_.B1 _1246_.B1 a_3247_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X10385 vssd1 _2009_.CLK a_2603_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10388 _0987_.B a_9963_15939# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X10389 vccd1 _1091_.X a_15365_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10391 _1022_.X a_17415_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10392 a_13136_5487# _0963_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X10393 vssd1 a_22806_20149# a_22764_20553# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10394 vccd1 _2023_.CLK a_1775_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10395 vccd1 _1165_.C a_6867_8545# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X10398 a_26099_20175# a_25401_20181# a_25842_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10400 a_19194_9411# _1577_.B a_19112_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10401 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_6808_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X10403 a_11061_13103# a_10791_13469# a_10971_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10405 vccd1 _1127_.A a_10730_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10406 a_6817_27023# _1286_.A1 _1287_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X10407 _1743_.A a_20263_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10408 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10409 a_27789_21807# a_26799_21807# a_27663_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10410 a_3247_13967# _1246_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.219375 ps=1.325 w=0.65 l=0.15
X10413 _0998_.B2 a_25439_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10414 a_25589_24527# _1513_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10415 a_4253_20719# _0913_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10417 vccd1 fanout33.A a_16863_27797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10418 a_12318_1247# a_12150_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10419 vccd1 a_11455_27515# a_11371_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10421 a_16083_17130# _1382_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10425 a_4517_1679# a_3983_1685# a_4422_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10426 vssd1 _1763_.A2 a_2970_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X10428 a_19057_14735# _1399_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10429 a_11023_7338# _1649_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10431 _1234_.Y _0925_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10432 vccd1 a_25071_19061# a_24987_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10434 vssd1 a_8548_23413# _1329_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10435 a_12189_18150# _0956_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X10437 a_25589_4943# _1960_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10438 vssd1 _1850_.CLK a_11711_13653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10439 _1282_.A2 a_9284_21781# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X10440 vssd1 a_19310_14709# a_19268_15113# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10441 vccd1 _1065_.B a_22195_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10442 _1856_.Q a_14123_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10443 a_20230_28447# a_20062_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10444 a_19107_2767# a_18243_2773# a_18850_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10445 a_21108_2223# a_20709_2223# a_20982_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10446 a_23351_32362# _1477_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10447 a_2777_17999# _1281_.B1 a_2861_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10448 a_6219_2589# a_5437_2223# a_6135_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10449 a_23224_2223# a_22825_2223# a_23098_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10450 a_25585_18543# a_25419_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10451 _1401_.A a_15387_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10452 a_10597_6825# _1189_.C1 a_10515_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10453 vssd1 _1775_.B1 a_1735_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X10454 a_3799_16911# _1291_.B1 a_3977_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10455 _1740_.X a_19619_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10456 _1562_.A a_12743_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10457 vssd1 a_23443_12778# _1979_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10459 a_5813_24527# _0909_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X10460 vccd1 _2005_.Q a_11895_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10461 a_17470_27765# a_17302_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10462 vccd1 a_13238_2741# a_13165_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10463 _1856_.Q a_14123_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10464 vssd1 _1907_.CLK a_14379_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10465 a_9999_31055# a_9301_31061# a_9742_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10466 vccd1 a_20775_27412# _1874_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10467 _1895_.Q a_24979_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10468 a_8004_25615# a_7755_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X10470 _1257_.X a_3087_20175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10471 a_27425_11293# a_26891_10927# a_27330_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10472 a_23535_23060# _1697_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10474 a_12575_8207# a_11711_8213# a_12318_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10475 a_9574_31055# a_9135_31061# a_9489_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10476 vssd1 a_5687_4564# _2001_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10477 a_12249_4943# _1751_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10478 _1905_.Q a_10995_19899# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10479 _1788_.X a_8624_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10480 a_18107_14954# _1574_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10483 vccd1 fanout37.A a_23395_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X10484 a_2658_27359# a_2490_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10485 vssd1 _1882_.CLK a_24591_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10486 vccd1 _1888_.Q a_18272_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10487 a_13130_5737# _0963_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X10488 vccd1 _0911_.A a_5455_20541# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10489 vssd1 _1768_.A _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10490 a_9779_11791# _1198_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10491 a_20421_15279# _1046_.B a_20349_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10492 vccd1 _0958_.B a_21095_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10493 a_20303_1501# a_19605_1135# a_20046_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10495 vssd1 _1823_.CLK a_24039_19093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10496 fanout37.A a_16311_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X10497 a_20267_14191# _1136_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10498 vssd1 a_2915_27613# a_3083_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10499 a_14910_2767# a_14637_2773# a_14825_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10500 _1112_.D1 a_19439_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10501 a_2143_17705# _1311_.A1 a_2225_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10503 vssd1 a_16290_4399# a_16396_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10504 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_8158_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X10505 vccd1 a_24811_28879# a_24979_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10506 vccd1 a_19405_15797# _1143_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X10507 _1010_.A a_13551_8215# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X10508 a_14944_4233# a_14545_3861# a_14818_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10509 vccd1 a_7683_1403# a_7599_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10510 _1721_.B a_27739_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10511 a_10386_29941# a_10218_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10512 a_10133_6031# _1563_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10513 _1557_.A a_8027_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10514 vssd1 _1969_.Q a_23757_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10516 vssd1 a_8307_5487# _1907_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10517 a_27590_3423# a_27422_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10518 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_9871_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10520 vccd1 clkbuf_1_1__f__0380_.A a_2686_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10521 _1511_.A a_20768_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10522 temp1.capload\[0\].cap.Y temp1.capload\[0\].cap.A a_26517_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10523 a_14453_16367# a_14287_16367# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10524 vccd1 _1894_.Q a_18699_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10525 a_25750_26271# a_25582_26525# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10526 a_20897_7663# _1996_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10528 vccd1 a_21115_27765# a_21031_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10529 a_18239_6941# a_18059_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10530 vccd1 _1870_.Q a_19286_28995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10531 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10532 a_19557_16395# _0939_.A a_19471_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10533 a_9889_15253# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X10534 a_2122_13469# a_1683_13103# a_2037_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10535 vssd1 a_23523_2589# a_23691_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10536 _1330_.X a_4035_30485# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10537 vccd1 _1985_.CLK a_26247_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10538 _1273_.A1 a_2807_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10539 a_27859_30676# _1450_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10541 a_27839_28701# a_27057_28335# a_27755_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10543 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10544 vccd1 a_15411_3829# a_15327_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10545 _0909_.A _0903_.C a_6981_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10546 vccd1 _1873_.CLK a_22843_29973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10547 vccd1 _1125_.X a_5578_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10548 a_16080_5487# _1047_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X10549 vccd1 _1590_.A_N a_20635_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X10550 vssd1 _1316_.X a_5241_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10552 vssd1 a_4627_6031# _1782_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10553 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10556 vssd1 _0987_.Y a_13632_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X10558 vccd1 a_17895_17973# a_17811_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10559 a_21923_16733# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10560 vccd1 a_2639_4943# a_2807_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10561 _1592_.X a_18560_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10562 a_18271_28879# a_17489_28885# a_18187_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10563 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10564 _1494_.A a_17088_26819# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10565 vssd1 _1999_.CLK a_11435_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10566 vccd1 a_25842_12533# a_25769_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10568 vccd1 a_9186_13255# _1199_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X10569 a_25589_23439# _1888_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10570 vccd1 _1985_.Q a_21042_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10571 vssd1 a_19405_15797# _1143_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X10572 vccd1 _1977_.Q a_22563_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10573 a_2649_23047# _1763_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X10575 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10576 _1767_.B a_4587_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10577 vssd1 a_25559_10602# _1720_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10578 a_10062_25398# _1274_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X10579 a_8919_16189# _1764_.A a_8828_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X10580 a_14039_31055# a_13257_31061# a_13955_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10581 a_26735_8029# a_25953_7663# a_26651_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10582 vssd1 fanout12.A a_7606_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10583 _1242_.B1 a_7479_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X10584 vccd1 fanout20.X a_21739_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10586 a_20982_8029# a_20543_7663# a_20897_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10587 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10588 vssd1 _1901_.Q a_8440_24643# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10589 a_2778_15529# _1219_.B1 a_2472_15431# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10590 a_24945_1135# _1668_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10591 vccd1 a_22063_11092# _1966_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10592 vccd1 a_27663_22173# a_27831_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10593 vssd1 _1018_.X a_15633_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X10595 vccd1 a_28135_13866# _1975_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10596 a_9123_19407# _1234_.A1 _1234_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X10597 vccd1 _1768_.A a_9503_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10598 vssd1 fanout24.A a_24039_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X10600 a_6733_11587# _1086_.B a_6651_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X10601 a_3514_25615# _1761_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X10602 a_18397_14013# _1721_.B a_18325_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10603 a_22162_31711# a_21994_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
R19 temp1.capload\[0\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10604 vccd1 _1010_.A a_11803_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10605 _1767_.Y _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10607 a_10543_29789# a_9761_29423# a_10459_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10608 vssd1 a_5416_21781# _1785_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X10609 a_23757_18365# a_23487_17999# a_23667_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10610 a_1855_16143# _1298_.A1 _1300_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X10611 vccd1 _1973_.Q a_28083_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10612 a_18682_2767# a_18243_2773# a_18597_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10614 vccd1 _1868_.Q a_14686_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10616 a_6981_12559# _0903_.C _0909_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10617 a_3965_16911# _1291_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X10618 a_20982_23261# a_20543_22895# a_20897_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10619 a_5345_30287# _1242_.A1 _1243_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X10620 vssd1 _0958_.B a_18453_25099# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X10621 a_25401_20181# a_25235_20181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10623 vssd1 _1880_.CLK a_16205_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10625 a_13165_2767# a_12631_2773# a_13070_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10626 vccd1 a_22143_26525# a_22311_26427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10628 a_4209_15279# _1278_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X10629 vccd1 a_12189_24825# a_12219_24566# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10632 io_out[6] a_21371_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10633 a_1769_15823# _1325_.A2 _1300_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10634 a_14449_24905# a_13459_24533# a_14323_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10635 vssd1 a_22081_13621# _1006_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X10637 a_27038_6687# a_26870_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10638 vssd1 _1152_.B a_18560_7913# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X10639 vssd1 a_2472_19605# _1312_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X10640 a_25800_27081# a_25401_26709# a_25674_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10641 a_24021_25621# a_23855_25621# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10642 a_3137_2773# a_2971_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10643 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10644 a_15461_3145# a_14471_2773# a_15335_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10645 vccd1 a_27498_11039# a_27425_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10646 vssd1 a_8818_11703# _1124_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10647 vssd1 _1199_.X _1250_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10648 a_10593_24233# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10649 vssd1 a_21150_2335# a_21108_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10650 vssd1 a_23266_2335# a_23224_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10651 vccd1 a_11391_23060# _1841_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10652 a_13633_16189# _0964_.A a_13551_15936# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10653 a_2309_29789# a_2143_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10654 a_4015_8779# _1177_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X10655 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10657 vccd1 clkbuf_0_net57.A a_2594_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10658 _1129_.B a_28015_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10659 _1177_.C a_7295_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10660 vssd1 _1532_.A a_12539_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X10661 a_12165_19453# a_11895_19087# a_12061_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10663 vssd1 a_6135_2589# a_6303_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10664 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_5816_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10665 a_6324_13353# _1316_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10666 _1830_.CLK a_15115_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X10667 vssd1 _1047_.C a_13061_7485# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
R20 temp1.capload\[3\].cap_48.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10668 a_16849_26159# _1840_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10669 vccd1 _2009_.CLK a_2051_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10670 _1781_.Y a_13019_20495# a_13257_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X10671 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_10048_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10672 a_10160_22729# a_9761_22357# a_10034_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10675 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4903_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X10676 a_5357_3087# _1809_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10683 a_1841_23439# _1270_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10684 vssd1 a_25271_17999# a_25439_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10686 vccd1 _1182_.B a_20390_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10687 vccd1 a_23691_11195# a_23607_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10688 a_24811_14735# a_23947_14741# a_24554_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10689 vssd1 _1999_.CLK a_14379_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10690 a_6917_7119# _1086_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X10691 vssd1 a_9889_25913# a_9823_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10692 a_18121_12925# _1965_.Q a_18049_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10693 a_17302_27791# a_17029_27797# a_17217_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10694 a_16734_8863# a_16566_9117# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10695 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_7564_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10696 _1467_.A a_14467_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10697 a_1673_22453# _2009_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X10699 a_5639_26703# _1762_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10701 a_15633_11445# _1118_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X10702 vssd1 _1242_.B1 _1243_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X10703 _1867_.Q a_17895_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10704 a_15939_28879# a_15759_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10705 vccd1 _0916_.A a_3247_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10706 vssd1 _1249_.A2 _1230_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X10707 a_11877_13653# a_11711_13653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10708 vssd1 a_24547_31274# _1447_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10710 vccd1 _0958_.B a_14747_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10711 a_20421_14191# _1136_.B a_20349_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10714 a_2686_26703# clkbuf_0_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X10716 _1170_.A3 a_4447_6581# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X10717 vssd1 a_10643_8207# a_10811_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10718 vccd1 _2009_.CLK a_3983_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10719 vssd1 _1133_.C a_18673_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10721 a_19388_22467# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10722 a_24481_14735# a_23947_14741# a_24386_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10723 _1736_.X a_21183_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X10724 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_15568_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X10725 a_22369_25615# _1833_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10726 a_13813_24527# _1819_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10727 _1773_.B a_4035_23957# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10728 a_26417_22895# _1968_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10729 _1221_.B a_3095_9867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X10730 a_10570_19743# a_10402_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X10731 _1091_.C1 a_16863_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10732 a_10344_20495# _0921_.B a_10154_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10733 _1187_.A a_18519_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10734 vssd1 a_8051_4667# a_8009_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10735 a_24547_31274# _1447_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10736 vccd1 _1985_.Q a_23299_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10737 vccd1 a_18539_1403# a_18455_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10738 a_15361_10927# _1088_.B a_15289_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10739 vccd1 _1544_.A_N a_9411_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X10742 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10743 a_10327_3855# a_10147_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10745 vssd1 a_22707_9514# _1926_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10746 vccd1 a_18539_32117# a_18455_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10747 a_26854_14303# a_26686_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10748 vssd1 a_5199_1403# a_5157_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10749 a_19593_7663# _1111_.B a_19521_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10750 a_11023_31274# _1479_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10751 a_14674_24233# _1056_.C1 a_14594_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10752 a_12425_22895# _1853_.Q a_11987_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10754 _1795_.X a_6324_13353# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10755 a_4811_26703# _1764_.B _1769_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10756 vccd1 _1850_.CLK a_6651_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10757 a_12253_24233# _0984_.B1 a_12337_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10758 _1255_.A1 a_2807_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10759 _1590_.X a_20815_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10760 a_16201_24349# a_15667_23983# a_16106_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10761 _0975_.X a_18887_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10762 vssd1 _1291_.A1 _1807_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10763 vccd1 _1764_.A a_10814_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10764 vccd1 a_11731_31867# a_11647_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10765 vccd1 _1530_.B a_19619_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10766 a_9920_25223# _1306_.A2 a_10062_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X10768 vssd1 a_9889_15253# a_9823_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10769 a_16911_32362# _1540_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10770 a_12575_29789# a_11877_29423# a_12318_29535# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10771 vccd1 _1327_.A2_N a_6186_21041# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
R21 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X10772 a_14839_25071# _1897_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10773 a_12153_23145# _1901_.Q a_12069_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10774 a_12035_2986# _1617_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10775 vssd1 a_26175_26427# a_26133_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10776 a_16293_8751# a_16127_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10777 a_10041_24527# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10778 vssd1 a_25842_16885# a_25800_17289# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10780 a_24639_14356# _1722_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10781 a_5871_23658# _1375_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10782 vccd1 _1850_.CLK a_14287_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10783 vccd1 a_8822_2741# a_8749_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10785 vccd1 a_13479_25589# a_13395_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10787 a_2309_3855# a_1775_3861# a_2214_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10788 a_22825_8751# a_22659_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10789 vccd1 _1901_.Q a_8522_24643# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10790 a_22181_2773# a_22015_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10792 a_22195_19087# a_22015_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10793 a_24757_17455# a_24591_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10794 a_4765_24759# _1763_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10795 vccd1 _1133_.C a_14655_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10796 a_13265_21807# _1021_.A a_13183_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10797 a_2214_6031# a_1775_6037# a_2129_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10798 a_12525_10383# _1848_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10800 a_25589_22351# _1879_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10801 vccd1 _1136_.B a_22563_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10802 vssd1 _1823_.Q a_21376_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X10804 vccd1 a_15795_25615# a_15963_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10805 a_16219_22057# _0966_.B1 a_16301_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X10806 vssd1 _1311_.B1 a_2472_19605# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X10807 a_5547_12015# _1218_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10808 a_15377_29423# _1858_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10809 a_3759_21237# _1312_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X10810 vccd1 a_28043_16042# _1976_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10811 _1120_.X a_14287_13353# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X10813 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10814 a_25156_23983# a_24757_23983# a_25030_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10816 vssd1 a_2195_12533# _1223_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X10817 vssd1 a_15795_25615# a_15963_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10818 vssd1 _1830_.Q a_15477_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10819 a_10643_6031# a_9945_6037# a_10386_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10821 vssd1 _0930_.Y _1334_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X10823 a_18808_3145# a_18409_2773# a_18682_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X10824 a_24761_17999# _1976_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10825 a_15483_15823# _1020_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10826 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10827 _1969_.Q a_24703_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10829 _1621_.X a_14283_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10830 vssd1 a_3835_2767# a_4003_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10832 a_21810_30877# a_21537_30511# a_21725_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X10835 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10836 a_17221_13353# _1147_.C1 a_17139_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10837 vssd1 a_23047_26677# a_23005_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10838 _1969_.Q a_24703_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10839 a_4847_25437# a_4149_25071# a_4590_25183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10840 vccd1 _1126_.Y a_4715_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X10841 a_27931_27613# a_27149_27247# a_27847_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10842 vssd1 _1133_.C a_17569_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X10843 a_26785_23983# _1885_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10844 a_3249_19453# _1231_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10845 vssd1 a_4739_7093# a_4697_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10846 a_3063_8751# _1170_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10847 _1872_.Q a_22403_30779# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10848 vssd1 _1861_.Q a_14557_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X10849 vccd1 a_15207_20719# _1484_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10850 _0956_.C a_7571_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X10851 a_23285_8213# a_23119_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10852 temp1.capload\[4\].cap.Y temp1.capload\[4\].cap.A a_23941_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10854 vssd1 a_19487_4564# _1636_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10855 vssd1 _1194_.B2 a_13464_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X10856 a_21136_11177# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10857 a_9128_27023# temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X10858 vccd1 _0918_.A a_10041_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10859 a_8027_18793# _1234_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10860 a_6588_16911# _1301_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10861 vssd1 a_8325_10901# a_8259_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10862 _1226_.A2 _1207_.B1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10863 a_4447_6581# _1159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10864 io_out[5] a_3759_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
X10865 a_20574_20291# _1506_.B a_20492_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10868 a_27590_12127# a_27422_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10869 a_18423_24527# a_18243_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X10870 _1140_.X a_10791_23552# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10871 _2009_.CLK a_2686_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10872 vccd1 a_19275_2741# a_19191_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10873 vccd1 _1189_.B2 a_10546_1385# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X10874 a_14081_31433# a_13091_31061# a_13955_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10877 a_17302_27791# a_16863_27797# a_17217_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
D4 vssd1 _1855_.D sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X10878 vccd1 a_6847_22057# _1328_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10879 a_14471_1501# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10881 vssd1 a_27847_12381# a_28015_12283# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10882 _1218_.B a_2715_13371# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10883 vssd1 a_19567_1679# a_19735_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10884 _2004_.D _1764_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10886 a_22369_24527# _1834_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10887 a_18475_30676# _1425_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10888 _1156_.Y _1156_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10889 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10890 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_18335_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X10891 vccd1 fanout37.A a_16863_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10892 a_22369_1135# _1957_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10893 vccd1 _1113_.C a_19807_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10894 vccd1 a_12743_8181# a_12659_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X10895 _1563_.A a_7980_9411# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10896 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10898 a_17029_1685# a_16863_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10899 a_6829_11587# _1086_.A a_6733_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10901 a_7442_17429# _1762_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3275 ps=1.655 w=1 l=0.15
X10902 a_27215_17130# _1389_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X10904 a_27061_8751# _1720_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10905 vssd1 a_24547_24746# _1880_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10908 a_10399_24527# _0921_.B a_10041_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10910 vssd1 _1230_.A4 a_2769_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X10911 vccd1 _1249_.A2 a_4932_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10912 vccd1 a_24554_14709# a_24481_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10913 _1725_.X a_23299_14557# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10914 a_25030_31965# a_24591_31599# a_24945_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10915 a_20303_29789# a_19439_29423# a_20046_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10916 _1300_.B1 _1232_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10917 vccd1 a_24639_18708# _1971_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10918 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10919 a_13587_29967# a_12889_29973# a_13330_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X10920 a_15189_29423# a_15023_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10921 a_25581_27247# a_24591_27247# a_25455_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X10922 a_12805_10089# _1069_.D a_12723_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X10923 _1130_.D1 a_19807_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X10924 vccd1 _1849_.CLK a_13643_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X10926 _1773_.Y _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10927 vccd1 _0925_.A2 a_4525_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X10928 vssd1 _0921_.A _0925_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X10930 vssd1 _1184_.B1 a_18416_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X10931 a_24547_24746# _1504_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10932 a_19734_15823# _1130_.C1 a_19654_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X10934 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10935 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10936 _1395_.A a_18100_19203# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10937 a_10188_18115# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10938 a_15477_14191# a_15207_14557# a_15387_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10939 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10940 _1587_.X a_21136_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10941 a_23535_23060# _1697_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X10942 vssd1 fanout20.X a_22659_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10944 a_5448_2767# _1807_.Y _1808_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X10945 a_1941_4399# a_1775_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X10946 a_19439_8751# _1152_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X10947 vccd1 _1775_.C1 a_5165_2828# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X10948 a_13306_9001# _1059_.X a_13057_8897# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X10949 vccd1 _1424_.A_N a_12079_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X10950 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10951 a_6713_16189# _1261_.A1 a_6641_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X10952 a_3087_20175# _1257_.B2 a_3281_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X10953 temp1.capload\[11\].cap.Y temp1.capload\[11\].cap.A a_22101_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10954 _1690_.A_N a_23671_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X10955 a_20690_28853# a_20522_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X10956 a_6968_25731# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10957 vccd1 _1047_.C a_14287_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X10958 _1039_.B a_12467_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10959 vssd1 _1242_.A2 a_7737_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X10960 vccd1 a_16274_24095# a_16201_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10962 _1066_.B a_23047_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10963 vccd1 _1896_.Q a_14927_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X10964 a_9644_23671# _1335_.A1 a_9786_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X10966 a_27517_10205# a_26983_9839# a_27422_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10967 a_14557_29245# a_14287_28879# a_14467_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X10968 a_18003_29789# a_17139_29423# a_17746_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X10969 _1542_.A a_13408_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10971 a_25129_3855# _1745_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10972 a_24025_11471# _1966_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X10974 vccd1 _0922_.Y a_2769_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X10975 a_24619_21263# a_23837_21269# a_24535_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X10976 _1381_.A a_14144_17027# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X10977 _1453_.X a_10419_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X10978 _1292_.C1 a_3799_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X10980 vccd1 _0921_.B a_8399_23492# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X10982 vssd1 a_15538_25589# a_15496_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X10983 a_27146_9117# a_26707_8751# a_27061_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10984 a_25030_9117# a_24591_8751# a_24945_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X10985 vccd1 _1849_.CLK a_19439_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10986 vccd1 _1887_.CLK a_26063_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X10987 vccd1 _1184_.A2 a_19605_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X10989 vccd1 a_21051_24746# _1887_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10990 _1188_.B a_5015_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10991 vssd1 a_16911_5162# _1942_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10992 a_5404_8323# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10993 _1308_.B a_9871_24527# a_10399_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10994 vccd1 _1021_.A a_17691_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10995 vssd1 a_10995_19899# a_10953_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X10996 a_17673_29789# a_17139_29423# a_17578_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X10997 vccd1 a_21143_21482# _1892_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X10999 vccd1 _1424_.A_N a_18059_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11000 a_13974_21237# a_13806_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11001 _0981_.B _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11002 _1525_.A a_22195_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11003 vccd1 _1061_.B a_22195_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11005 a_9761_27797# a_9595_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11006 vssd1 _1195_.B2 a_16408_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X11008 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11009 a_2217_13469# a_1683_13103# a_2122_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11010 a_27149_3311# a_26983_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11012 a_22199_14557# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11013 _1132_.C a_10865_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X11014 vccd1 _1150_.A2 a_17262_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X11015 a_2340_6409# a_1941_6037# a_2214_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11016 a_2009_21263# _1259_.X a_1643_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11018 vssd1 _1261_.X a_9135_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X11019 a_5271_14191# _1217_.A2 a_5177_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X11020 _1723_.B a_27279_14459# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11021 vssd1 _1941_.CLK a_18243_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11022 a_7550_2589# a_7277_2223# a_7465_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11023 vssd1 a_2807_3829# _1304_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11025 a_17888_29257# a_17489_28885# a_17762_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11026 _1240_.B1 a_2603_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11027 a_24389_15829# a_24223_15829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11030 _1104_.X a_15115_14851# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X11031 a_6467_9001# _1122_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11032 vccd1 _0984_.A2 a_12337_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X11033 vccd1 _1876_.CLK a_22291_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11034 a_26785_17455# _1525_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11035 a_2214_4943# a_1775_4949# a_2129_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11037 vccd1 _0930_.A a_9961_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X11038 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11039 _1074_.C a_9195_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11041 a_27245_10927# _1586_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11044 vssd1 a_24075_16911# a_24243_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11045 _1974_.Q a_25255_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11046 a_22438_29535# a_22270_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11047 a_21150_23007# a_20982_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11048 a_23523_22173# a_22825_21807# a_23266_21919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11049 _0921_.B a_3983_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11050 vccd1 _1775_.A2 a_1975_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X11051 a_21176_16143# _1970_.Q a_20601_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X11053 a_9013_6397# _1188_.B a_8941_6397# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11055 vssd1 _1269_.A1 _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X11056 _1318_.X a_5487_5281# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11057 vssd1 a_22063_11092# _1966_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11058 vssd1 _1242_.A2 a_6817_27023# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X11059 a_7015_19881# _1325_.B1 a_6797_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X11060 a_5301_23983# _1337_.S a_5203_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X11061 _1883_.Q a_26267_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11063 vccd1 _1032_.C a_18887_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11064 _0911_.A a_2623_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11065 vccd1 _1338_.A a_27811_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11067 vccd1 a_27831_15547# a_27747_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11068 _1043_.B a_16607_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11069 vccd1 _1873_.CLK a_25235_26709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11070 vccd1 a_22751_22895# _1882_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11071 vssd1 a_9894_17429# _0981_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11073 _1727_.X a_23483_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11074 vccd1 a_13599_7828# _1749_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11076 _1314_.X a_6559_15936# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11077 a_12199_20495# a_11907_20175# a_12113_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X11078 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11079 a_22285_4221# a_22015_3855# a_22195_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11080 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11081 a_13671_29967# a_12889_29973# a_13587_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11082 vssd1 _1033_.A2 a_20337_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X11083 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_10699_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11085 vccd1 _2005_.Q a_6927_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X11087 vssd1 _2005_.Q a_9195_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X11088 a_16573_4399# a_16396_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11090 vccd1 _0958_.B a_16495_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11091 a_23745_23439# a_23211_23445# a_23650_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11092 a_5545_22057# _1775_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X11093 vssd1 _1823_.CLK a_26799_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11096 a_17029_27797# a_16863_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11097 vccd1 a_26099_26703# a_26267_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11098 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11099 a_25539_27613# a_24757_27247# a_25455_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11101 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_15943_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11102 vssd1 _1289_.B1 a_5692_15253# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X11105 _1310_.Y _1308_.Y a_5813_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X11106 _1057_.B a_24151_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11107 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_16955_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11108 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11109 vccd1 _1273_.A1 a_7479_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X11110 a_1828_14709# _1230_.B1 a_2220_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X11112 a_25639_3855# a_24941_3861# a_25382_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11113 a_7619_2986# _1660_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11114 vccd1 _1183_.A2 a_22563_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11115 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_5639_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11116 a_9284_21781# _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X11117 vccd1 temp1.capload\[10\].cap.A temp1.capload\[10\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11118 vssd1 a_27498_11039# a_27456_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11119 a_10862_27613# a_10589_27247# a_10777_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11120 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X11121 _0922_.Y _0918_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11122 a_25559_21482# _1699_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11123 a_9937_4917# _1293_.A1 a_10190_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X11125 vssd1 _1138_.X a_14655_18115# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11126 vssd1 a_27222_16479# a_27180_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11128 vssd1 a_12467_25339# a_12425_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11129 vssd1 a_11391_23060# _1841_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11130 a_11689_31599# a_10699_31599# a_11563_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11132 a_20072_18543# _1885_.Q a_19497_18689# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X11133 a_19651_17999# a_18869_18005# a_19567_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11136 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13544_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11138 a_18239_27613# a_18059_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11139 a_7843_26703# _1261_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11141 vssd1 _1032_.C a_20421_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11142 vccd1 a_20046_29535# a_19973_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11143 vccd1 _1353_.Y a_7479_28887# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11148 vssd1 a_13183_20719# _0964_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11149 a_24823_28010# _1551_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11151 a_8937_29967# a_8760_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11152 a_16657_23983# a_15667_23983# a_16531_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11153 a_15151_16733# a_14287_16367# a_14894_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11154 a_16911_32362# _1540_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11155 a_14931_27791# _0965_.B1 a_15013_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11157 _1308_.Y _0909_.A a_23849_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11158 vccd1 a_16921_14709# _1091_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X11159 vssd1 _1086_.Y _1289_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11161 vssd1 _1020_.A2 a_16208_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X11162 vccd1 a_25639_16733# a_25807_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11163 a_22454_1501# a_22015_1135# a_22369_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11164 vccd1 _1907_.CLK a_11895_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11165 a_1955_14441# _1223_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11166 a_4627_13967# _1217_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11168 a_19701_31055# _1473_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11170 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11171 a_20709_2223# a_20543_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11172 a_22825_2223# a_22659_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11173 a_17831_11092# _1583_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11174 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11175 a_25313_21807# _1877_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11176 a_13517_14709# _1107_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X11177 vccd1 _1202_.Y a_6559_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X11178 a_7749_9839# _1158_.X a_7531_9813# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X11179 vssd1 _1086_.Y a_6731_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11180 vssd1 _1896_.CLK a_20083_28885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11181 _1474_.A_N a_8215_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X11182 a_19562_15529# _1537_.B a_19480_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11183 a_25030_6941# a_24757_6575# a_24945_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11184 a_10386_6005# a_10218_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11185 a_11842_10089# _1438_.B a_11685_9813# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11186 vccd1 _0963_.B a_16159_20747# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X11188 vccd1 _1486_.B a_13455_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11189 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8392_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11190 vssd1 _1855_.CLK a_9779_29973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11191 a_17470_29941# a_17302_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11192 vccd1 a_17746_29535# a_17673_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11193 vccd1 a_1643_21781# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11194 _1141_.C a_10667_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11195 vccd1 _1590_.A_N a_20267_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11196 a_20690_27765# a_20522_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11197 vccd1 _1775_.A2 _1781_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11198 a_25156_8751# a_24757_8751# a_25030_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11200 a_7479_28585# _1242_.B1 _1274_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X11201 vssd1 a_25455_27613# a_25623_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11202 a_27272_8751# a_26873_8751# a_27146_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11203 vssd1 a_17139_9839# _1293_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X11204 vssd1 _1882_.CLK a_24959_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11205 vccd1 _0911_.A a_3548_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X11206 a_26996_13103# a_26597_13103# a_26870_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11207 vssd1 _1941_.CLK a_20543_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11210 vccd1 _1208_.A1 a_1775_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11211 a_27031_29588# _1352_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11212 vssd1 _0921_.Y _0922_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11213 a_3345_19131# _1231_.B2 a_2836_19319# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X11214 a_17443_31965# a_16661_31599# a_17359_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11215 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11217 a_25455_1501# a_24757_1135# a_25198_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11219 _1760_.B temp1.inv2_2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11220 vssd1 _1764_.B a_4441_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11221 vccd1 a_12759_15645# a_12927_15547# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11222 a_2217_8029# a_1683_7663# a_2122_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11223 a_22553_20175# _1822_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11224 vssd1 _1459_.A a_12815_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X11225 a_21150_7775# a_20982_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11226 a_22162_31711# a_21994_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11227 vssd1 _1270_.A a_2787_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11228 _0930_.B _0921_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11229 fanout33.A a_16863_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X11231 _1775_.A2 a_2327_20183# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11232 _1080_.B a_25623_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11234 vssd1 _2005_.Q a_11711_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X11235 a_9921_16911# _1764_.A a_10279_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11237 a_4256_14191# _1231_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X11238 a_19142_1679# a_18703_1685# a_19057_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11239 a_17736_5263# _0963_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X11240 a_26099_26703# a_25235_26709# a_25842_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11242 vssd1 a_25566_21919# a_25524_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11243 a_27747_22173# a_26965_21807# a_27663_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11244 _1226_.A1 a_1775_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11245 vccd1 a_22567_25071# _1873_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X11246 a_15163_4564# _1621_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11248 a_24903_19087# a_24205_19093# a_24646_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11249 _1254_.A2 a_2143_17705# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X11250 a_5629_7663# _1172_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X11251 vssd1 fanout24.A a_26983_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11252 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11253 _1412_.A a_20171_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11254 vccd1 _1187_.A a_15549_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X11255 _1623_.X a_12488_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11256 a_22063_5162# _1672_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11258 a_27479_16733# a_26615_16367# a_27222_16479# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11259 vccd1 a_20701_14709# _0953_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X11260 a_7019_1679# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11261 vccd1 a_12575_1501# a_12743_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11262 a_2340_5321# a_1941_4949# a_2214_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11263 vssd1 _0963_.B a_17017_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11264 a_14537_9001# _1193_.X a_14465_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11265 vccd1 a_5231_22869# _1307_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X11266 vssd1 _0965_.B1 a_15656_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X11267 vssd1 _1075_.C a_18397_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11268 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_6559_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11269 _1863_.Q a_18355_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11270 a_23316_22729# a_22917_22357# a_23190_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11271 a_13809_1679# a_13275_1685# a_13714_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11273 _1818_.Q a_10627_27765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11274 vssd1 _1974_.Q a_27713_11837# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11275 a_12349_23983# _1902_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11276 a_6651_23439# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11277 a_13408_3561# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11279 a_24278_10357# a_24110_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11280 a_8548_23413# a_8399_23492# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X11281 vccd1 _1459_.A a_11711_16919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11282 vccd1 temp1.capload\[9\].cap.A temp1.capload\[9\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11283 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11284 vccd1 _1489_.A_N a_20819_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11286 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11287 vccd1 a_5031_1501# a_5199_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11288 a_27973_19631# a_26983_19631# a_27847_19997# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11291 a_24757_28335# a_24591_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11292 vssd1 a_2455_2589# a_2623_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11293 vccd1 _1451_.B a_7567_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11297 a_27149_16733# a_26615_16367# a_27054_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11298 _1706_.X a_22931_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11300 a_3063_14191# _1249_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11301 a_4606_1501# a_4333_1135# a_4521_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11302 _1150_.A2 a_24887_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11303 vccd1 a_23818_23413# a_23745_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11304 _1555_.A a_7935_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11305 a_26091_3677# a_25309_3311# a_26007_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11307 vccd1 a_18187_28879# a_18355_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11308 a_14361_7125# a_14195_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11311 a_11693_17821# _2006_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X11312 vccd1 _1046_.B a_23299_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11313 vccd1 a_15725_7809# _1050_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X11314 _1404_.A a_19619_19997# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11317 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_10140_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11318 a_21978_30623# a_21810_30877# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11319 vccd1 a_25750_26271# a_25677_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11320 a_10279_16911# _1764_.A a_9921_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11321 vssd1 a_3111_5652# _0916_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11324 _1329_.S a_8548_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11325 vssd1 a_8143_2491# a_8101_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11327 a_4069_5737# _1281_.A1 _1804_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11328 a_10769_8585# a_9779_8213# a_10643_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11329 vssd1 a_25198_17567# a_25156_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11330 _1611_.X a_9360_3971# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X11332 _1065_.X a_15299_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11333 a_22369_26703# _1839_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11334 a_4127_22869# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X11335 a_11760_23671# _1306_.A2 a_11902_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X11336 a_25129_16367# _1985_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11337 a_21143_23658# _1406_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11338 _1586_.A a_19480_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11339 a_10951_24233# a_10423_23983# _1270_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11340 a_26628_22895# a_26229_22895# a_26502_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11341 vccd1 _1823_.CLK a_26799_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11342 a_12237_19453# _2004_.Q a_12165_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X11343 a_20758_10499# _1577_.B a_20676_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11344 a_4989_16367# a_4719_16733# a_4899_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11347 vccd1 _1055_.C a_13367_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11348 a_24205_11471# a_23671_11477# a_24110_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11349 a_9547_22895# _1306_.A2 a_9184_23047# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X11350 a_1775_12265# _1250_.A1 a_1857_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X11351 vccd1 a_2594_31055# clkbuf_0_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X11352 vccd1 _1277_.B a_3063_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11354 vssd1 _1476_.B a_12625_32509# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11355 vccd1 a_12743_29691# a_12659_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11356 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_11619_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11357 a_12907_7232# _1039_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11358 a_20850_15823# _1081_.D1 a_20601_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X11359 vccd1 a_25439_2741# a_25355_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11360 vssd1 _0958_.B a_18121_12925# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11361 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11362 vssd1 _1830_.CLK a_22050_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11363 a_12679_31764# _1473_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11364 vccd1 _1153_.A a_20267_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11365 vccd1 clkbuf_1_1__f__0380_.A a_2686_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11366 vssd1 _1850_.CLK a_6651_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11368 a_14195_13647# _1050_.B a_14449_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11369 _1660_.X a_12351_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11370 vssd1 a_10883_21271# _1132_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X11371 a_22580_1135# a_22181_1135# a_22454_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11373 a_20666_20969# _1506_.B a_20584_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11374 vssd1 _0958_.B a_20421_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11375 a_20414_32117# a_20246_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11376 a_6607_30186# _1555_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11377 a_14743_29967# a_14563_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11378 a_23358_22325# a_23190_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11380 a_19609_29967# a_19432_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11383 a_22879_2767# a_22015_2773# a_22622_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11384 a_27713_11837# a_27443_11471# a_27623_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11385 vccd1 fanout28.A a_16311_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X11386 a_7657_16617# _1234_.A2 _1291_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X11387 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_13367_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11388 vssd1 a_26007_3677# a_26175_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11389 a_1849_13103# a_1683_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11390 a_16991_9117# a_16127_8751# a_16734_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11391 vccd1 _1313_.A a_2327_20183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11392 vccd1 _1544_.A_N a_7663_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11393 _1156_.D a_16863_11177# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X11395 a_26517_31375# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11396 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11397 vssd1 _0921_.A a_8548_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11400 vssd1 _1850_.CLK a_14287_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11402 vccd1 _1074_.C a_18519_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11403 a_11023_5652# _1355_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11404 _2007_.Q a_5015_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11405 a_20709_22895# a_20543_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11406 a_11685_9813# _0952_.A1 a_11938_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X11407 vssd1 _1074_.C a_15361_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11408 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11409 a_20522_27791# a_20083_27797# a_20437_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11410 vccd1 _1053_.A a_15299_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X11412 vssd1 _1975_.Q a_27897_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11413 vssd1 a_25198_8863# a_25156_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11414 a_20246_32143# a_19973_32149# a_20161_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11415 vssd1 a_27314_8863# a_27272_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11416 vssd1 _1347_.Y a_8767_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11417 a_4433_17999# _1267_.B1 a_4517_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11418 vssd1 _1788_.X a_7008_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
R22 vssd1 temp1.capload\[8\].cap_53.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11419 a_10543_27791# a_9761_27797# a_10459_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11420 _1103_.A1 a_25807_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11421 vssd1 _1140_.C a_11957_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11422 a_22195_10383# a_22015_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11423 a_27337_5487# _1728_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11427 a_18468_5737# _1607_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11428 vssd1 a_2623_6843# a_2581_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11429 vssd1 _1873_.CLK a_21555_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11430 vssd1 a_7803_6740# _1753_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11431 a_6981_12559# _1255_.A1 a_6559_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11433 vccd1 a_21039_4765# a_21207_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11434 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE a_8951_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X11435 a_7479_17277# _2004_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X11436 vssd1 _1878_.Q a_20169_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11437 vccd1 _1882_.CLK a_24959_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11438 vssd1 a_22622_2741# a_22580_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11439 a_22622_1653# a_22454_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11440 _1504_.A a_21827_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11442 _1393_.A a_18560_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11443 a_23119_13647# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11444 vccd1 _1088_.B a_14283_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11445 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11449 a_18187_28879# a_17323_28885# a_17930_28853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11450 a_25455_2589# a_24591_2223# a_25198_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11451 vccd1 a_11759_32362# _1467_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11453 a_6073_25045# _1305_.B a_6230_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X11454 vssd1 _1277_.B a_4983_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X11455 a_27789_15279# a_26799_15279# a_27663_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11456 a_27571_2589# a_26707_2223# a_27314_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11457 vssd1 a_18371_31055# a_18539_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11458 a_25455_17821# a_24591_17455# a_25198_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11459 vccd1 a_18059_9839# _1153_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11460 a_20249_28885# a_20083_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11461 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11462 a_27364_20719# a_26965_20719# a_27238_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11463 a_19268_2057# a_18869_1685# a_19142_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11464 vccd1 a_26267_20149# a_26183_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11465 a_17946_32143# a_17673_32149# a_17861_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11466 vssd1 _1338_.A a_27811_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11467 _1844_.Q a_20655_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11469 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_8307_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X11471 a_22898_27765# a_22730_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11472 _0987_.Y _0961_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11473 a_12625_32509# a_12355_32143# a_12535_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11474 a_2915_24349# a_2051_23983# a_2658_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11477 vccd1 _2004_.Q a_12061_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X11478 vccd1 a_25198_6687# a_25125_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11479 a_25858_18909# a_25419_18543# a_25773_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11480 a_11527_4765# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11481 vssd1 a_15151_10205# a_15319_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R23 vssd1 temp1.capload\[5\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11482 _2003_.D _1762_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11483 a_13337_21807# _1857_.Q a_13265_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11484 a_22063_18218# _1527_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11485 _1175_.B2 _0930_.A a_10515_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11486 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X11487 vccd1 a_14335_25834# _1431_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11488 vccd1 a_17647_23658# _1839_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11489 a_1823_19796# _1776_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11490 a_20083_3855# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11492 a_23450_29941# a_23282_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11493 _1140_.C a_7442_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11494 a_16170_5487# _1195_.A2 a_16080_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X11495 a_9742_7093# a_9574_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11496 a_20897_7663# _1996_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11497 a_2585_24349# a_2051_23983# a_2490_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11498 _1631_.X a_17227_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11499 a_14921_10499# _1007_.X a_14839_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11500 a_2326_32509# _1337_.A1 a_1827_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11501 a_10459_29789# a_9595_29423# a_10202_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11503 _1418_.A a_16904_22467# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11505 _1394_.A a_23323_18811# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11506 a_5692_15253# _1325_.A2 a_6084_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X11507 a_22879_1679# a_22181_1685# a_22622_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11508 vssd1 _1965_.Q a_22837_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11509 a_12886_25615# a_12613_25621# a_12801_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11510 a_17647_23658# _1418_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11511 vccd1 a_19310_14709# a_19237_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11512 _1730_.X a_23759_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11513 vssd1 _1887_.CLK a_25235_20181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11514 _1081_.B1 a_21463_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11515 a_22143_26525# a_21445_26159# a_21886_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11516 vssd1 fanout21.X a_24407_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11517 vccd1 _1685_.A_N a_22567_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11518 a_23282_29967# a_23009_29973# a_23197_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11519 a_12752_22351# _0983_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X11520 vssd1 a_9999_7119# a_10167_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11521 vccd1 _1448_.A a_11711_15831# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X11522 a_14345_15425# _1095_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11523 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11524 vccd1 _1047_.C a_15391_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11527 a_27897_15101# a_27627_14735# a_27807_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11528 _1195_.B2 a_23967_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11529 a_16734_8863# a_16566_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11530 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11531 vssd1 a_15081_12533# _1104_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X11532 a_13625_24533# a_13459_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11533 _1068_.A1 a_15503_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11534 _1083_.A a_7867_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11535 vssd1 _1762_.A _0951_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11536 a_17323_12015# _1098_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11537 a_9828_26935# _1328_.A1 a_9970_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X11538 vssd1 a_24887_1653# a_24845_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11540 a_19961_10749# _1129_.B a_19889_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X11541 vccd1 _1887_.Q a_20574_20291# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X11542 a_4517_25437# a_3983_25071# a_4422_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11543 _1941_.CLK a_13643_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X11545 vccd1 _1313_.X _1786_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11546 a_18869_1685# a_18703_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11547 vccd1 a_24278_11445# a_24205_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11548 a_20246_32143# a_19807_32149# a_20161_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11549 a_20169_19453# a_19899_19087# a_20079_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11550 vssd1 _0987_.B _0987_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11551 _1080_.B a_25623_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11552 vccd1 _0921_.B a_10423_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11553 vssd1 _1246_.A2 a_1791_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X11554 _1293_.A1 a_17139_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X11555 _1165_.C _1123_.X a_6835_7439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11557 vssd1 _1079_.B a_21733_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11558 vccd1 a_11759_1898# _1956_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11560 vccd1 a_15319_10107# a_15235_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11561 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11562 a_27337_9839# _1926_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11563 a_8522_10499# _1782_.A a_8440_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11564 a_25731_11293# a_24867_10927# a_25474_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11566 a_5980_29673# a_5731_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X11568 a_6828_31375# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11570 vssd1 _1390_.B a_22285_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11571 _1025_.B a_15227_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11572 a_9999_7119# a_9301_7125# a_9742_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11574 vssd1 a_7442_17429# _1140_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.212875 pd=1.305 as=0.08775 ps=0.92 w=0.65 l=0.15
X11575 vccd1 a_12759_4943# a_12927_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11576 vssd1 _1155_.C a_16863_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11577 _1250_.B2 _1311_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X11578 _1020_.A2 a_19471_16395# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X11579 _1775_.X a_1735_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11580 _1313_.X a_5455_20541# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X11581 a_17473_15797# _1028_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X11582 a_4859_5162# _1364_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11583 vccd1 a_18751_5162# _1923_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11584 a_18371_31055# a_17507_31061# a_18114_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11585 a_3881_16911# _0925_.A2 a_3799_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11586 vccd1 _1132_.A a_17139_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11587 _1373_.A a_7015_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11588 a_2932_18517# _1325_.B1 a_3324_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X11589 a_4713_12015# _1222_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11590 vccd1 a_1643_23413# io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11591 a_27153_21807# _1878_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11592 _1328_.S a_6847_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X11593 vccd1 a_7883_4765# a_8051_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11594 vccd1 _1090_.C a_17323_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11595 a_17946_32143# a_17507_32149# a_17861_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11596 a_23005_25993# a_22015_25621# a_22879_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11597 vssd1 a_27463_17723# a_27421_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11598 _1569_.A a_10511_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11599 vssd1 _1459_.A a_21187_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X11600 _1154_.A1 a_23691_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11601 a_25030_15645# a_24591_15279# a_24945_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11602 a_19605_20969# _1883_.Q a_19521_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11603 a_24205_19093# a_24039_19093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11604 vssd1 a_18291_2388# _1628_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11605 a_2037_13103# _1810_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11606 a_10147_26409# _0983_.B1 a_10229_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11607 a_18041_31055# a_17507_31061# a_17946_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11608 vccd1 _0911_.A a_6559_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11609 a_15285_32143# _1868_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11610 a_8213_25335# _0909_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X11611 vssd1 a_27590_27359# a_27548_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11612 vssd1 a_22659_17455# _1823_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11615 a_11789_25071# _1852_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11616 vssd1 _1313_.X a_6713_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11617 a_10154_20495# _0921_.B a_10344_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11618 vssd1 _1145_.A1 a_8669_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X11620 _1720_.A a_22195_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11621 vssd1 a_17470_27765# a_17428_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11622 a_4863_23413# _2009_.CLK a_5145_23759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X11623 a_16904_20291# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11624 _1058_.B a_7683_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11625 a_8031_17999# _1764_.A a_8449_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11626 _1965_.Q a_26267_12533# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11627 a_25765_16367# a_24775_16367# a_25639_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11629 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11630 a_15512_12559# _0997_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X11631 a_22745_29199# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11632 a_24895_28879# a_24113_28885# a_24811_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11633 a_10287_26742# _1328_.A1 a_9828_26935# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X11634 a_8355_11254# _1124_.X a_7896_11079# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X11636 vssd1 _1852_.Q a_9268_24233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X11637 a_16760_14191# _1394_.A a_16185_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X11638 a_25125_6941# a_24591_6575# a_25030_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11639 a_17831_11092# _1583_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11640 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11641 a_21177_13103# _0939_.A a_21095_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11642 a_3325_2767# _1951_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11643 vccd1 _1849_.CLK a_20543_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11644 vccd1 _1127_.A a_14379_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11645 _1965_.Q a_26267_12533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11646 vccd1 a_16623_2589# a_16791_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11647 vccd1 _1277_.A a_4897_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X11648 vccd1 _1144_.B a_6739_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11649 vssd1 a_10811_1653# a_10769_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11650 vccd1 a_25842_23413# a_25769_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11651 vccd1 a_6705_16341# _1789_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X11653 a_5509_17973# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X11655 a_7360_15095# _1218_.B a_7288_15095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11656 a_17415_13760# _1023_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11657 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5908_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X11658 a_14921_26409# _0966_.B1 a_15005_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11659 _1097_.X a_13551_15936# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11660 _1547_.A a_11476_20969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11662 a_12069_23145# _1186_.C1 a_11987_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11663 vccd1 a_27571_9117# a_27739_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11664 vssd1 a_25559_21482# _1699_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11666 a_22285_17277# a_22015_16911# a_22195_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11667 a_17221_17277# _1132_.A a_17139_17024# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11668 a_25198_13215# a_25030_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11669 a_26651_4765# a_25787_4399# a_26394_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11670 a_2692_19631# _1311_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X11671 a_4669_9839# _1298_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X11673 a_3977_17231# _1291_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11674 a_24945_31599# _1873_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11675 vssd1 _1325_.X a_4404_18517# vssd1 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X11676 a_16863_11177# _1154_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11677 a_25708_26159# a_25309_26159# a_25582_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11678 a_4525_20175# _1273_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X11679 _1329_.A0 a_1674_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11681 vccd1 a_3759_21237# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X11682 a_27973_9839# a_26983_9839# a_27847_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11684 vccd1 a_2658_24095# a_2585_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11685 a_12885_15279# a_11895_15279# a_12759_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11686 vccd1 _1234_.A2 a_4517_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X11687 a_6671_17231# _0930_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X11689 _2023_.CLK a_2686_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11690 a_17565_24129# _1134_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11691 a_26283_18909# a_25419_18543# a_26026_18655# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11692 vccd1 _1291_.A1 a_5547_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11693 a_14643_13647# _1049_.X _1050_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11694 _1222_.A1 a_5303_9633# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X11695 a_6641_24893# _0911_.A a_6559_24640# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11696 vssd1 a_5271_20719# _1353_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X11697 a_18545_13131# _1110_.A a_18459_13131# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11698 _1876_.CLK a_21831_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X11699 vssd1 a_23783_22325# a_23741_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11700 a_12723_10089# _1069_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X11702 vssd1 a_16382_25071# a_16488_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11703 _1103_.D1 a_15943_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
R24 vccd1 temp1.capload\[6\].cap_51.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X11704 a_9163_2767# a_8381_2773# a_9079_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11705 a_10125_5487# a_9135_5487# a_9999_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11706 a_11287_3677# a_10589_3311# a_11030_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11707 vccd1 _1020_.X a_15483_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11708 vssd1 a_3635_24501# a_3593_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11710 _1832_.Q a_23323_24251# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11711 vccd1 _0985_.A a_15825_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X11712 vssd1 _2005_.Q a_11711_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11713 a_20709_4765# a_20175_4399# a_20614_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11714 _1609_.X a_16307_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X11715 a_5908_5737# _1797_.Y _1798_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X11716 _1797_.Y _1234_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11717 vccd1 a_4774_1247# a_4701_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11718 a_10413_11177# _1051_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11719 a_1898_11587# _1781_.Y a_1816_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11720 a_12985_2767# _1955_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11721 vssd1 _1198_.A2 a_8955_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X11723 a_1849_7663# a_1683_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11724 a_20860_19881# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11725 vssd1 a_21039_4765# a_21207_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11726 a_25589_16911# _1527_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11727 a_6829_3133# a_6559_2767# a_6739_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11728 a_2030_1501# a_1757_1135# a_1945_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11730 a_16304_30511# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11731 a_27847_27613# a_26983_27247# a_27590_27359# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11732 vccd1 _1139_.C a_10731_17483# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X11733 vssd1 a_10195_13268# _1906_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11734 a_17117_8751# a_16127_8751# a_16991_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11735 a_27422_3677# a_27149_3311# a_27337_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11736 a_26601_14191# _1984_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11737 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11738 a_10041_24527# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11739 _2004_.D _1775_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11741 vssd1 fanout21.X a_22659_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11742 a_17853_30345# a_16863_29973# a_17727_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11744 vccd1 a_19487_26922# _1875_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11745 vssd1 _2009_.CLK a_1959_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11747 a_19793_1135# _1945_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11748 _1132_.X a_14839_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11749 vccd1 _2023_.CLK a_1591_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11750 a_3961_3145# a_2971_2773# a_3835_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11751 vssd1 a_20046_29535# a_20004_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11752 vssd1 a_20471_26427# a_20429_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11753 a_12843_4943# a_12061_4949# a_12759_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11754 vccd1 _1140_.C a_9687_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11755 a_12535_32143# a_12355_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11756 a_10585_28169# a_9595_27797# a_10459_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11757 a_2787_20719# _1269_.B1 a_2965_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X11758 a_7704_3561# _1448_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11759 _0906_.X a_8213_25335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11760 a_2382_4511# a_2214_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11761 a_20303_5853# a_19605_5487# a_20046_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11762 a_13721_21263# _1851_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11763 _1011_.A1 a_10811_6005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11764 vssd1 _1532_.A a_5731_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11766 vssd1 a_20775_27412# _1874_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11767 a_19487_26922# _1494_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11768 a_26183_12559# a_25401_12565# a_26099_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X11769 vssd1 a_12743_13621# a_12701_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11770 a_14465_13353# _1116_.X a_14369_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X11771 vccd1 a_13551_17999# _0958_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X11772 a_28135_13866# _1703_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11773 _1189_.C1 a_8859_6144# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X11774 vssd1 a_11777_9269# _1192_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X11775 vccd1 a_23691_22075# a_23607_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11776 a_17305_13353# _1528_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X11777 a_10643_6031# a_9779_6037# a_10386_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11778 a_2594_31055# clkbuf_0_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11779 a_14453_8207# _1149_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X11780 a_21886_26271# a_21718_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11781 a_22238_13647# _1032_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X11783 vccd1 a_18114_31029# a_18041_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11784 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11785 a_21073_11849# a_20083_11477# a_20947_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11786 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X11787 a_10041_24527# _0921_.B a_10399_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11789 a_11711_7663# _1148_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X11790 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11791 vssd1 a_2566_25183# a_2524_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11792 a_26597_23983# a_26431_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11794 vssd1 a_17746_29535# a_17704_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11795 vccd1 a_26670_23007# a_26597_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11797 temp1.capload\[12\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11798 _1802_.X a_4116_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X11799 vccd1 _1816_.CLK a_7939_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11800 a_10218_6031# a_9779_6037# a_10133_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11802 vssd1 a_25623_24251# a_25581_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11804 a_9574_5853# a_9301_5487# a_9489_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11805 vssd1 a_25071_19061# a_25029_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11808 a_7566_28335# _1242_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X11809 _1639_.X a_12815_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X11811 vssd1 a_14345_15425# _1095_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X11812 vssd1 a_11759_32362# _1467_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11813 vccd1 _1074_.C a_13275_17024# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11815 vssd1 _0935_.X a_13551_8215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11816 a_26007_29789# a_25143_29423# a_25750_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11819 _1696_.B a_26451_18811# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11821 a_2413_12559# _1222_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X11822 vccd1 a_13587_29967# a_13755_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11824 vccd1 _1179_.B2 a_19562_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X11825 vssd1 a_3945_4917# _2020_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X11826 a_8480_12879# _1034_.Y a_8177_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X11829 a_25413_30287# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11830 vssd1 _1133_.C a_17625_22923# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X11833 vccd1 a_22063_8426# _1916_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11834 a_8395_12559# _1050_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11835 a_22825_24349# a_22291_23983# a_22730_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11839 a_21183_2767# a_21003_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11840 a_27422_27613# a_27149_27247# a_27337_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11841 _1079_.B a_25899_11195# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11842 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X11843 a_25677_29789# a_25143_29423# a_25582_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11844 _1646_.X a_13455_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X11846 a_21494_20969# _1506_.B a_21412_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11847 a_7573_11791# _1156_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X11848 a_12189_23737# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X11854 vccd1 _1568_.B a_10511_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11855 vssd1 a_12679_31764# _1473_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11856 vssd1 a_22546_6031# a_22652_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11857 vssd1 _1873_.CLK a_21831_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11858 a_3993_27497# _1764_.Y a_4248_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11859 vssd1 fanout37.A a_20543_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11860 vccd1 a_25623_2491# a_25539_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11863 a_25401_6037# a_25235_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11864 a_23649_10927# a_22659_10927# a_23523_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X11867 a_24945_5487# _1593_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11869 a_4213_30663# _1337_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X11870 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X11871 _1270_.Y _1270_.A a_24677_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11872 vssd1 _1070_.A2 a_17485_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X11873 a_12893_12559# _1911_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X11874 vccd1 a_17895_27765# a_17811_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X11875 a_14829_19631# _0964_.A a_14747_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11876 vccd1 a_19567_17999# a_19735_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11878 a_27061_8751# _1720_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11880 vssd1 _0963_.B a_16189_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11881 _1773_.Y _1773_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11882 a_20171_24349# a_19991_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11883 vccd1 a_25842_22325# a_25769_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11884 io_out[0] a_1643_21781# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11885 a_25198_2335# a_25030_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11886 vssd1 a_7883_4765# a_8051_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11887 _1257_.B1 _1254_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11888 vssd1 a_20046_1247# a_20004_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11889 a_24757_28335# a_24591_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11890 a_4213_30663# _1337_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X11891 vssd1 _1855_.CLK a_9595_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11892 a_22457_27797# a_22291_27797# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11894 a_4701_1501# a_4167_1135# a_4606_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11895 vssd1 _0981_.B a_13245_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11896 a_26026_18655# a_25858_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11897 a_22369_2767# _1993_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11898 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11900 vccd1 _1145_.B2 a_11707_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11901 a_13445_31055# _1856_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11902 a_6559_26703# _1286_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11903 a_24301_28879# _1895_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X11904 a_25401_24533# a_25235_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11906 vccd1 a_27111_14557# a_27279_14459# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11907 vssd1 a_5031_1501# a_5199_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11908 vccd1 _1896_.CLK a_19439_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11909 vccd1 _1835_.Q a_20171_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11910 _0958_.A a_13551_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X11911 a_13104_12937# a_12705_12565# a_12978_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11912 vccd1 _1544_.A_N a_7847_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X11913 a_15795_31055# a_14931_31061# a_15538_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11914 vccd1 a_26026_18655# a_25953_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11915 vccd1 _1907_.CLK a_14195_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11917 a_18642_7913# _1577_.B a_18560_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X11918 a_5301_23983# _1294_.B2 a_5392_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11920 a_7933_8573# a_7663_8207# a_7843_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X11921 vccd1 _1139_.C a_14747_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11922 a_6646_27023# _1242_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X11923 vssd1 a_14802_7093# a_14760_7497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11924 vccd1 _0939_.A a_18151_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11925 vssd1 _1999_.CLK a_9595_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11926 _1532_.A a_2327_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X11927 vssd1 a_2807_6005# a_2765_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X11929 _1807_.Y _1321_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11931 a_14905_18115# _1134_.X a_14833_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X11933 _1141_.C _1269_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11934 a_15462_29789# a_15023_29423# a_15377_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11935 a_20947_28879# a_20249_28885# a_20690_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X11937 a_15465_31055# a_14931_31061# a_15370_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11938 vccd1 _1139_.C a_10055_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X11939 vssd1 _1924_.CLK a_24591_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X11940 vssd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11941 a_10506_30511# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11942 vccd1 a_13875_23658# _1840_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11943 a_2836_19319# a_2966_19131# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X11944 _1764_.A a_6927_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11945 a_10971_13469# a_10791_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11947 vccd1 _1855_.CLK a_10699_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11948 vssd1 a_26099_26703# a_26267_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11949 io_out[6] a_21371_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X11950 vccd1 _1849_.CLK a_16113_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11952 a_27295_13469# a_26431_13103# a_27038_13215# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11953 vssd1 a_17102_31711# a_17060_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11954 temp1.inv2_2.A a_2686_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11955 _1882_.CLK a_22751_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X11956 vccd1 _1823_.CLK a_22291_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11957 vccd1 a_22622_24501# a_22549_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11958 _1075_.X a_17691_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X11959 a_4899_16733# a_4719_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X11960 a_22751_15645# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11961 _1272_.B1 a_1779_22453# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X11962 a_1925_21807# _1242_.A2 a_1841_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11965 a_13587_29967# a_12723_29973# a_13330_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X11966 vccd1 a_26479_11690# _1716_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X11967 vccd1 _1242_.A2 a_7479_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X11968 vssd1 _1769_.B1 _1769_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X11969 _1316_.X a_6870_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X11970 a_27590_9951# a_27422_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11971 _1485_.A a_19204_28995# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X11972 a_12532_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X11973 vccd1 _1969_.Q a_23667_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X11974 _1979_.Q a_24979_14709# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11975 a_20073_13353# _1006_.X a_19991_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11976 a_26870_24349# a_26431_23983# a_26785_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X11977 vccd1 _1126_.Y _1170_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11978 a_5573_5281# _1255_.A1 a_5487_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X11979 a_2339_32143# _1337_.A0 a_1827_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X11980 a_23726_8181# a_23558_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X11981 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_10948_28585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X11982 a_23224_10927# a_22825_10927# a_23098_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11983 _0966_.X a_14839_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11984 vssd1 a_9644_23671# _1336_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X11987 a_2616_23983# a_2217_23983# a_2490_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X11988 a_5455_20541# _1313_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X11989 vssd1 a_17565_24129# _1134_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X11992 _1111_.B a_23691_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11993 a_13257_29967# a_12723_29973# a_13162_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11994 _1337_.A0 clkbuf_1_1__f_net57.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X11995 vssd1 a_22983_21482# _1885_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11996 a_18059_27613# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11997 a_8675_22351# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X11998 a_10957_3677# a_10423_3311# a_10862_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X11999 vccd1 _1218_.B a_4351_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X12000 a_21143_8916# _1604_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12001 vccd1 a_11287_27613# a_11455_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12002 a_4903_19631# _1233_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X12003 vccd1 _1999_.CLK a_14471_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12005 a_10202_22325# a_10034_22351# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12006 a_2199_21583# _1242_.A2 a_2009_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12007 a_19567_17999# a_18703_18005# a_19310_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12008 vssd1 a_6611_29111# _1259_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12010 a_10344_6409# a_9945_6037# a_10218_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12011 a_11312_16367# a_11269_16600# a_11240_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X12012 _2009_.CLK a_2686_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12013 vccd1 a_2198_1247# a_2125_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12014 _1279_.A1 _1158_.X a_7573_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12015 a_12000_25071# a_11601_25071# a_11874_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12016 a_5278_22390# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X12017 _1194_.B2 a_13663_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12018 vssd1 a_14066_24501# a_14024_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12020 _1397_.A a_16904_20291# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12022 vssd1 a_28043_16042# _1976_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12024 vssd1 _1855_.CLK a_12723_29973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12025 a_23849_26159# _1308_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12026 vccd1 a_22898_24095# a_22825_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12027 a_17139_11584# _1977_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12029 vccd1 _1885_.Q a_20666_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12031 a_15737_15823# _1029_.X a_15931_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12032 a_9945_8213# a_9779_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12033 a_10727_29967# a_9945_29973# a_10643_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12034 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X12035 vssd1 _1217_.A3 a_4627_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12036 a_12334_4943# a_11895_4949# a_12249_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12037 vccd1 a_20775_30186# _1871_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12038 a_15969_13131# _0935_.X a_15883_13131# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12039 a_2639_3677# a_1941_3311# a_2382_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12041 a_19237_17999# a_18703_18005# a_19142_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12042 _1886_.Q a_27923_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12043 a_10034_22351# a_9761_22357# a_9949_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
R25 vccd1 temp1.capload\[14\].cap_44.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12044 clkbuf_0_net57.X a_2594_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12045 a_21617_18543# _1879_.Q a_21545_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12048 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_8109_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X12050 vssd1 _1192_.A2 a_9773_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12051 a_11934_9295# _1139_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X12053 _1107_.X a_13091_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12054 a_7295_6031# _1171_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12055 a_20613_28335# a_19623_28335# a_20487_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12056 a_8301_15055# a_8109_14796# _1793_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X12057 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_6559_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R26 temp1.capload\[12\].cap.A vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12058 a_4876_27791# a_4627_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12059 _2004_.D _1242_.A1 a_4441_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12060 vccd1 a_28015_26427# a_27931_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12061 vssd1 a_10257_27001# a_10191_27069# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X12063 vccd1 fanout24.A a_23671_10389# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12064 a_10839_10602# _1436_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12065 a_4213_24135# _1763_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X12066 _1775_.C1 a_7387_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12069 a_4163_4943# _1780_.B1 a_3945_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X12070 _1197_.D a_14287_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X12071 vccd1 _1855_.CLK a_13091_31061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12072 vccd1 temp1.capload\[8\].cap_53.LO temp1.capload\[8\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12073 vccd1 _1021_.A a_13183_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12074 a_7939_13647# _1175_.B2 _1175_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12076 a_17359_31965# a_16495_31599# a_17102_31711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12077 a_12383_25437# a_11601_25071# a_12299_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12078 a_15696_21263# _1074_.X a_15594_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X12079 a_12610_10383# a_12171_10389# a_12525_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12080 a_11711_12672# _1092_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12082 vccd1 a_3210_24501# a_3137_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12083 a_20629_6575# a_20359_6941# a_20539_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12084 vccd1 a_16911_31274# _1896_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12085 vssd1 _1081_.C1 a_20601_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X12087 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_4811_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12088 vccd1 a_21511_28500# _1870_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12089 _1291_.A1 a_2623_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12090 vccd1 a_7531_9813# _1159_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X12091 a_20429_13103# _1007_.A1 a_19991_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12092 vccd1 a_21051_4074# _1743_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12093 vccd1 a_24535_10383# a_24703_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12094 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12098 _1136_.B a_25531_9269# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12100 _1502_.A a_20079_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12101 a_23481_16367# a_23211_16733# a_23391_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12104 vccd1 _1780_.B1 a_7189_13408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X12105 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X12106 a_4337_25071# _2007_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12107 a_9489_7119# _1812_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12108 a_13432_26703# a_13183_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12110 a_27215_17130# _1389_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12111 _1194_.A2 a_17895_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12112 a_25731_11293# a_25033_10927# a_25474_11039# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12114 a_25125_21085# a_24591_20719# a_25030_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12115 a_25842_20149# a_25674_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12117 vssd1 a_2836_19319# _1233_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12119 a_10034_2589# a_9595_2223# a_9949_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12120 vssd1 _1234_.A2 a_4903_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12121 a_9037_19087# _1234_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X12122 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12123 vssd1 a_10202_22325# a_10160_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12124 vccd1 a_15538_31029# a_15465_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12125 vccd1 _1125_.X a_4519_9991# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X12126 _2007_.D _1771_.B a_1591_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12127 vssd1 a_20690_27765# a_20648_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12128 vccd1 _1139_.C a_11711_12672# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12129 vssd1 a_11023_18218# _1820_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12130 a_7366_15279# a_7189_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12131 vccd1 _1104_.X a_9779_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12132 vssd1 a_18187_28879# a_18355_28853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12133 a_14604_27497# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12135 a_25309_26159# a_25143_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12137 _1179_.B2 a_21115_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12138 vccd1 a_10459_27791# a_10627_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12139 a_13521_22895# _1868_.Q a_13449_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12140 vccd1 a_7387_15823# _1775_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12142 a_17710_7119# _1062_.X a_17630_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12143 vccd1 a_15319_30779# a_15235_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12144 a_25674_20175# a_25401_20181# a_25589_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12145 temp1.capload\[9\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12146 a_5271_26409# _1353_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12147 a_9613_16600# _1269_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12149 a_24945_2223# _1743_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12150 vssd1 _1110_.A a_18059_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12151 a_24462_1653# a_24294_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12152 a_19977_28335# _1429_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12153 a_10202_27765# a_10034_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12154 vccd1 a_27590_3423# a_27517_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12155 vccd1 _1242_.B1 _0909_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12156 vccd1 a_17831_30676# _1471_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12158 a_21051_24746# _1519_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12160 a_14287_8207# _0991_.X a_14465_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X12161 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12163 vccd1 a_27038_13215# a_26965_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12164 a_22963_1501# a_22181_1135# a_22879_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12166 a_27146_9117# a_26873_8751# a_27061_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12168 a_25030_1501# a_24591_1135# a_24945_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12171 vccd1 a_17013_19777# _1024_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X12172 _1207_.B1_N a_4015_8779# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X12173 vccd1 _1893_.Q a_17630_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12174 a_9921_16911# _1764_.A a_10279_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12175 vccd1 a_13047_12180# _1911_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12176 a_10543_2589# a_9761_2223# a_10459_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12177 a_18475_30676# _1425_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12178 vccd1 _1764_.B a_4248_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12180 vssd1 _1171_.Y a_7295_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12181 _1594_.X a_17456_7913# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12182 a_2125_1501# a_1591_1135# a_2030_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12185 a_5047_21237# _1292_.C1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X12186 a_13698_31029# a_13530_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12187 a_2122_9839# a_1945_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12188 a_2726_11587# _1221_.B a_2644_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12189 vccd1 io_in[0] a_2962_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12190 vccd1 _1051_.A1 a_8522_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12193 vccd1 a_10811_6005# a_10727_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12194 _1429_.A a_18239_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12196 a_15453_8751# _1059_.B a_15381_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12198 a_7013_28157# a_6743_27791# a_6923_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12199 _1270_.A a_10423_23983# a_10951_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12200 a_13047_12180# _1569_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12201 a_22396_29423# a_21997_29423# a_22270_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12202 a_21108_22895# a_20709_22895# a_20982_23261# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12203 _1750_.X a_9683_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X12204 vssd1 a_23903_24746# _1881_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12205 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_6808_29673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12206 a_22181_25621# a_22015_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12207 vssd1 _0929_.A a_3983_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X12208 vccd1 a_6610_13879# _1263_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X12209 a_11425_8751# _1010_.A a_11343_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12210 _1842_.Q a_22587_31867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12211 _1481_.A a_14604_27497# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12212 vssd1 a_24639_18708# _1971_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12213 _1398_.X a_15479_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12214 a_1945_9295# _1780_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12215 a_13452_26159# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12216 vccd1 a_21787_8916# _1591_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12217 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12218 a_24535_10383# a_23671_10389# a_24278_10357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12219 vccd1 _0935_.X a_17967_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12221 _1191_.B1 a_19103_13985# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X12222 vccd1 a_9742_5599# a_9669_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12223 vccd1 _1304_.B _1794_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12224 vccd1 a_9135_25071# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12225 vccd1 a_15078_2741# a_15005_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12226 a_14449_13647# _1050_.B a_14195_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12228 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12230 a_9142_14774# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X12231 a_11777_9269# _0991_.X a_11934_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12232 _1551_.A a_8440_24643# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12234 vccd1 _0987_.Y a_10681_6825# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X12235 a_12460_5321# a_12061_4949# a_12334_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12236 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4876_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12237 a_23745_16911# a_23211_16917# a_23650_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12238 a_16577_12015# _1010_.A a_16495_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12240 _1572_.B a_15319_10107# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12241 vssd1 clkbuf_0_temp1.i_precharge_n.X a_5354_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12242 a_24757_20719# a_24591_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12243 vccd1 a_2455_6941# a_2623_6843# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12244 temp1.capload\[7\].cap.Y temp1.capload\[7\].cap.A a_24769_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12245 a_25566_21919# a_25398_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12246 _1723_.A_N a_22015_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X12247 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12248 vccd1 a_28015_19899# a_27931_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12249 vccd1 _1123_.X a_6717_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X12250 vccd1 _1067_.B a_7199_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12251 _1113_.C a_11693_17821# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X12252 a_1791_13647# _1301_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X12253 a_2673_7663# a_1683_7663# a_2547_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12254 a_2953_20969# _1269_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X12255 a_5547_7913# _1210_.B a_5629_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12256 a_1644_18517# _1311_.A1 a_1864_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12258 a_26597_13103# a_26431_13103# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12259 a_2639_4765# a_1775_4399# a_2382_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12260 a_21031_11471# a_20249_11477# a_20947_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12261 a_2999_27613# a_2217_27247# a_2915_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12262 a_21718_26525# a_21445_26159# a_21633_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12263 vccd1 a_20690_28853# a_20617_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12265 a_8785_20473# _1232_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X12266 a_25674_20175# a_25235_20181# a_25589_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12267 vssd1 a_10459_2589# a_10627_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12268 vccd1 fanout21.X a_23565_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X12269 vccd1 a_11023_7338# _1649_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12270 a_18601_16911# _1179_.B1 a_18685_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12271 temp1.capload\[6\].cap.B a_15750_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12272 a_10459_27791# a_9595_27797# a_10202_27765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12273 a_4517_17999# _1267_.B2 a_4433_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12274 a_8381_2773# a_8215_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12275 a_13057_8897# _1057_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X12276 a_22504_12559# _1151_.X a_22402_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X12278 vccd1 a_10257_27001# a_10287_26742# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12279 a_4441_26159# _1764_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X12280 _1858_.Q a_16055_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12282 a_21249_13103# _1079_.B a_21177_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12283 a_3605_8207# _0930_.B _1289_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X12284 a_11053_31599# _1855_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12285 vccd1 a_2287_16885# _1231_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12286 vssd1 a_10627_27765# a_10585_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12287 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13432_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12288 vssd1 a_21235_7338# _1924_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12289 a_7637_8751# _1162_.X a_7553_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X12290 a_1779_22453# _1242_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X12291 vccd1 a_25198_20831# a_25125_21085# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12293 vssd1 a_10167_5755# a_10125_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12295 vccd1 fanout21.X a_24591_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12296 _1086_.B _1084_.C1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12297 a_9841_6575# _1144_.B a_9769_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12298 a_25213_16201# a_24223_15829# a_25087_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12299 vssd1 a_15299_18543# _0961_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12300 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X12301 vssd1 a_10202_29535# a_10160_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12302 a_17415_20719# _1876_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12303 vccd1 a_13783_5162# _1610_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12304 a_23523_9117# a_22659_8751# a_23266_8863# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12305 vccd1 _1861_.Q a_14467_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12306 vssd1 a_8307_16367# _0935_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12307 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_4811_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12308 a_17293_17277# _1822_.Q a_17221_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12309 _1175_.Y _0930_.A a_8387_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12310 vccd1 a_5455_14735# _1231_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12312 vssd1 a_20487_28701# a_20655_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12313 a_25030_7119# a_24757_7125# a_24945_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12314 a_10103_23478# _1335_.A1 a_9644_23671# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X12315 a_17727_27791# a_17029_27797# a_17470_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12316 vssd1 a_17159_9019# a_17117_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12317 vssd1 _1768_.A a_9687_12919# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X12319 vssd1 _1074_.C a_17017_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12320 a_14641_30511# _1447_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12321 _1242_.B1 a_7479_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12323 vssd1 _0930_.A _0930_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12324 a_24945_15279# _1975_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12325 a_10160_2223# a_9761_2223# a_10034_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12326 a_25589_6031# _1591_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12327 _1168_.X a_6867_8545# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X12328 a_17041_12879# _1830_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X12330 vssd1 _1038_.C1 a_12873_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X12331 a_24110_10383# a_23837_10389# a_24025_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12332 a_7289_2045# a_7019_1679# a_7199_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12333 _1530_.B a_24243_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12334 a_2582_1679# a_2309_1685# a_2497_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12337 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12338 a_5565_22649# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X12339 _1391_.A a_22195_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12340 a_25283_14356# _1706_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12341 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12342 a_23408_30345# a_23009_29973# a_23282_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12343 _1544_.A_N a_8307_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X12344 a_9683_8029# a_9503_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12345 vccd1 a_10643_29967# a_10811_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12346 _1836_.Q a_28015_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12347 _1530_.B a_24243_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12348 a_25125_31965# a_24591_31599# a_25030_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12350 _1604_.X a_20447_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X12351 _1038_.D1 a_16035_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12352 vccd1 a_14839_11471# _1127_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12353 a_25674_4943# a_25401_4949# a_25589_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12354 a_3181_9867# _1177_.B a_3095_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12355 vssd1 _1830_.CLK a_22935_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12356 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_4903_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12357 _1098_.B a_23691_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12358 _1719_.B a_26819_7931# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12359 _1052_.B1 _1198_.A2 a_10413_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X12361 _1484_.B a_15207_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X12363 vccd1 _1234_.A2 a_3965_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X12364 a_24577_15823# _1701_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12365 temp1.dcdc.A a_5354_28335# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12366 vccd1 _1763_.A2 a_5099_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X12368 a_23542_3829# a_23374_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12369 a_1945_8207# _1786_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12370 a_7442_3829# a_7274_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12371 vssd1 a_13599_7828# _1749_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12372 _1680_.A a_22563_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12373 a_18087_29789# a_17305_29423# a_18003_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12374 vssd1 a_2382_28447# a_2340_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12376 a_14549_7119# _1759_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12377 vssd1 a_7571_14191# _1374_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X12378 vccd1 _1924_.CLK a_24591_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12379 _1056_.C1 a_15851_22895# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12382 a_25156_1135# a_24757_1135# a_25030_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12383 vssd1 a_25198_28447# a_25156_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12384 _0951_.B _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12385 _1677_.X a_21827_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X12387 vssd1 a_7111_25071# _1242_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X12388 vssd1 a_1737_14165# _1277_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12389 a_23013_3311# _1989_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12390 vccd1 _0952_.A1 a_18979_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12393 a_8387_13647# _1766_.A0 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X12394 a_26229_22895# a_26063_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12395 _1786_.A1 _1313_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12397 a_8177_21781# _1270_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X12398 vssd1 _1261_.A1 a_5183_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X12399 a_27038_24095# a_26870_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12400 a_27847_26525# a_27149_26159# a_27590_26271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12401 a_10399_24527# a_9871_24527# _1308_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12405 a_12189_23737# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X12406 vssd1 _1252_.A a_5731_12567# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12407 a_21235_31274# _1486_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12409 a_22580_31433# a_22181_31061# a_22454_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12410 vssd1 _1448_.A a_8215_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12412 a_22645_23983# _1832_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12413 a_14802_7093# a_14634_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12414 a_22334_15055# _1973_.Q a_22244_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X12415 a_14537_13353# _1120_.B a_14465_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12416 vssd1 a_27831_20987# a_27789_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12417 a_16439_3677# a_15741_3311# a_16182_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12418 vssd1 _0917_.A a_2971_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X12419 vssd1 _1999_.CLK a_9779_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12420 a_1775_12265# _1250_.A1 a_1857_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12421 a_21695_19796# _1393_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12422 a_20349_17455# _1127_.A a_20267_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12423 _1566_.X a_8579_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12424 a_16159_9867# _0939_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12425 a_9000_14967# _1772_.A0 a_9142_14774# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X12426 _1156_.Y _1071_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12427 a_2198_8181# a_2030_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12428 vccd1 a_23818_16885# a_23745_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12429 a_14453_30511# a_14287_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12431 a_23266_8863# a_23098_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12432 a_26007_3677# a_25143_3311# a_25750_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12433 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_9595_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12434 vccd1 _1744_.A_N a_20359_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12436 a_13360_28335# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12438 vssd1 _0999_.C1 a_16863_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X12439 vccd1 _1039_.B a_7786_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12440 a_4847_1679# a_3983_1685# a_4590_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12442 _1027_.X a_17139_17024# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12443 vssd1 a_7975_2589# a_8143_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12444 a_24462_25589# a_24294_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12445 vssd1 _1055_.C a_14563_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12447 a_22063_5162# _1672_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12448 vssd1 _1530_.B a_19709_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12449 a_2686_23439# clkbuf_1_1__f__0380_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12450 a_19746_23555# _1506_.B a_19664_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12451 a_17017_10749# _1089_.B a_16945_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12453 a_10229_26409# _1818_.Q a_10147_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12454 a_26996_17455# a_26597_17455# a_26870_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12455 vssd1 a_10814_14709# _0951_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12456 _2021_.D a_5349_3616# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X12457 temp1.capload\[6\].cap.Y temp1.capload\[6\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12458 a_20387_1501# a_19605_1135# a_20303_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12459 vccd1 _0951_.B a_15299_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12460 vccd1 a_10021_9985# _1012_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X12461 a_6151_22869# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X12462 a_23542_3829# a_23374_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12463 a_18329_6575# a_18059_6941# a_18239_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12464 vssd1 a_20046_31711# a_20004_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12465 vssd1 a_5048_14165# _1249_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X12466 _0994_.B2 a_18539_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12467 a_7442_3829# a_7274_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12469 a_21143_8916# _1604_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12470 vssd1 a_7625_26677# _1261_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12471 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X12472 a_25455_5853# a_24757_5487# a_25198_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12473 a_19562_25321# _1484_.B a_19480_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12474 a_27973_12015# a_26983_12015# a_27847_12381# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12475 a_27931_12381# a_27149_12015# a_27847_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12476 a_24757_20719# a_24591_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12477 a_24159_23439# a_23377_23445# a_24075_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12478 a_22195_21263# a_22015_21263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12479 a_24294_25615# a_24021_25621# a_24209_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12480 _1490_.A a_18607_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12481 vccd1 _1074_.C a_13367_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12482 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_7606_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12483 vssd1 a_21115_28853# a_21073_29257# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12485 vssd1 _1886_.Q a_21181_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12486 a_8449_17999# _1764_.A a_8031_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12487 vccd1 a_26099_12559# a_26267_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12488 a_25539_13469# a_24757_13103# a_25455_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12489 vssd1 a_4590_1653# a_4548_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12491 vssd1 _1896_.Q a_15017_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12492 vssd1 _1205_.A1 a_4167_8527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X12494 a_26091_26525# a_25309_26159# a_26007_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12497 vccd1 _1010_.A a_12907_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12498 vccd1 a_20690_27765# a_20617_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12499 vssd1 _1147_.X a_16863_11177# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X12500 a_2639_28701# a_1775_28335# a_2382_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12502 vccd1 a_20315_26922# _1895_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12503 vccd1 _1884_.Q a_21494_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12504 vccd1 _0958_.A a_21463_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12505 a_3133_2057# a_2143_1685# a_3007_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12506 a_11759_7338# _1657_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12507 vssd1 _1143_.X _1156_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X12508 vssd1 a_26099_12559# a_26267_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12509 _0985_.X a_15575_19881# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X12510 vccd1 a_10167_4667# a_10083_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12511 vccd1 _1286_.A1 a_6457_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X12512 a_23266_27359# a_23098_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12513 vssd1 _0984_.A2 a_12425_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X12514 vccd1 _1860_.CLK a_11711_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12515 a_25455_28701# a_24591_28335# a_25198_28447# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12516 a_19405_15797# _1130_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X12517 vssd1 a_25991_22075# a_25949_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12518 vccd1 a_24087_13866# _1967_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12519 vccd1 _1127_.A a_17415_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12520 a_9937_4917# _0988_.X a_10094_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X12521 vssd1 _1353_.A _1347_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12523 a_14369_9001# _1196_.D a_14287_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X12524 a_3299_22325# _1337_.S a_3730_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X12525 _1020_.B1 a_13919_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12527 a_8395_22057# _0922_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12528 vssd1 _1141_.C a_15269_9661# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12529 a_1828_14709# _1277_.A a_2048_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12530 vccd1 fanout20.X a_24591_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12532 vccd1 _1544_.A_N a_14287_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12533 a_12321_22325# _1142_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X12534 a_22063_29098# _1490_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12535 a_18785_27791# _1872_.Q a_18703_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12536 vccd1 a_4220_21959# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X12537 a_24087_13866# _1686_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12538 a_1757_8213# a_1591_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12540 vccd1 a_25198_31711# a_25125_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12541 a_4428_14441# _1278_.X a_4173_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X12542 a_2290_7775# a_2122_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12543 vssd1 a_5693_16341# _1267_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X12544 vccd1 _1075_.C a_17999_16395# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X12545 a_12065_11471# _1847_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12546 a_18703_27791# _0965_.B1 a_18785_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X12547 _1024_.A2 a_17541_15307# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X12548 _1265_.A1 _1231_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12549 vssd1 a_2455_6941# a_2623_6843# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12551 vssd1 _1072_.X a_14379_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X12553 vssd1 _1033_.A1 a_19112_9411# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12554 _1057_.B a_24151_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12555 a_17302_29967# a_16863_29973# a_17217_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12557 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_5639_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12558 _1050_.Y _1049_.X a_14643_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12559 vccd1 _1277_.B a_1965_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12560 vssd1 a_17381_7093# _1069_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X12561 a_19709_24893# a_19439_24527# a_19619_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12563 _1353_.A a_5271_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X12564 a_2685_22057# _0925_.Y a_2769_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12565 a_4598_21807# _1242_.B1 a_4220_21959# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X12566 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_16304_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X12567 _1034_.Y _1034_.D a_15931_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12569 a_22622_26677# a_22454_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12570 vccd1 a_20839_32117# a_20755_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12572 a_23983_8207# a_23119_8213# a_23726_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12573 a_6073_25045# _1242_.A1 a_6326_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X12574 a_13551_11471# _1071_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12575 a_14441_17455# _1852_.Q a_14369_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12576 _1222_.B1 a_2644_11587# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12577 _1843_.Q a_23875_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12578 _1447_.A a_9268_24233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X12580 a_26225_22729# a_25235_22357# a_26099_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12582 vssd1 _0999_.X a_14839_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X12583 _1896_.CLK a_18830_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12584 vssd1 _1829_.Q a_15569_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12585 vccd1 a_27314_8863# a_27241_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12586 a_27153_15279# _1389_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12587 a_9601_13353# _1198_.A2 a_9186_13255# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X12588 vssd1 a_10839_10602# _1848_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12589 vssd1 _1817_.Q a_7105_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12590 vccd1 a_20499_23658# _1835_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12591 a_10731_17483# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12592 a_20303_31965# a_19439_31599# a_20046_31711# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12593 a_22015_15823# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12594 a_20539_3677# a_20359_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12595 vssd1 a_25198_1247# a_25156_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12596 a_12989_7485# _1010_.A a_12907_7232# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12597 _1057_.X a_15115_9408# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12598 _1326_.A3 _1231_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12599 vccd1 a_25198_7093# a_25125_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12600 vccd1 a_12771_21482# _1901_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12601 a_17342_19881# _1022_.X a_17262_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12602 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_15483_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12603 _1094_.X a_12907_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12605 a_2214_28701# a_1941_28335# a_2129_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12606 vccd1 a_13551_17999# _0958_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12607 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5888_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X12608 a_5520_10933# _0916_.A a_5448_10933# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X12609 a_2594_31055# clkbuf_0_net57.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X12611 a_11874_2589# a_11601_2223# a_11789_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12612 a_5115_1501# a_4333_1135# a_5031_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12613 _1033_.A2 a_18551_11809# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X12614 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12615 a_27755_28701# a_27057_28335# a_27498_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12616 a_14024_24905# a_13625_24533# a_13898_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12617 vccd1 _1267_.A1 a_4069_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X12618 a_25125_8213# a_24959_8213# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12620 a_17047_4765# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12621 a_26099_12559# a_25235_12565# a_25842_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12622 _1764_.B a_1766_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12623 a_6651_5853# _1782_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12624 a_18100_19203# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12625 vssd1 a_2382_4917# a_2340_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12626 a_14287_5487# _1066_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12627 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X12628 a_20954_15055# _0952_.A2 a_20864_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X12629 a_7381_13103# a_7189_13408# _1791_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X12631 vssd1 a_17749_9269# _1120_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X12632 vssd1 _1020_.A2 a_21176_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X12633 vssd1 a_25750_29535# a_25708_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12634 a_7843_26703# _1242_.B1 a_7625_26677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X12635 a_14335_25834# _1431_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12636 _1306_.A2 _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12639 a_6559_15936# _1261_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12641 vccd1 _1873_.Q a_18607_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12642 vccd1 a_23323_27765# a_23239_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12643 vccd1 _1132_.C a_16711_22923# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X12645 vssd1 a_13035_10383# a_13203_10357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12646 a_16064_19087# _1020_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X12647 _1889_.Q a_23691_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12649 a_9183_12180# _1570_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12650 vssd1 a_9275_24746# _1900_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12651 a_20131_21972# _1523_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12652 a_23098_4943# a_22825_4949# a_23013_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12653 io_out[3] a_4863_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12654 vccd1 a_21150_23007# a_21077_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12655 vssd1 a_2198_8181# a_2156_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12656 vccd1 _1250_.A1 a_1775_10496# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12658 a_4314_7093# a_4146_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12659 _1719_.B a_26819_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12660 vccd1 a_23875_29941# a_23791_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12661 vccd1 a_27847_3677# a_28015_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12662 a_12901_10089# _1069_.C a_12805_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X12663 vssd1 _1053_.A a_10883_21271# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12664 vccd1 a_9460_15431# _1199_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X12665 vssd1 _1532_.A a_9135_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12666 a_5701_12015# _1218_.B a_5629_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12668 _1216_.A2 _1246_.B2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12669 vssd1 a_23395_17455# _1887_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12670 a_24639_12180# _1709_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12672 a_2962_14735# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X12673 a_2132_16367# _1249_.A1 a_1829_16341# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X12674 a_27931_5853# a_27149_5487# a_27847_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12675 a_11023_5652# _1355_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12676 vccd1 a_11711_25615# _1855_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12677 a_5437_2223# a_5271_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12678 a_6736_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12679 a_27238_22173# a_26799_21807# a_27153_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X12680 vccd1 a_2807_4667# a_2723_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12681 vssd1 a_21787_8916# _1591_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12682 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE a_7790_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X12683 vssd1 a_2971_16367# _0921_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X12686 vccd1 a_21235_25236# _1883_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12687 vssd1 _1887_.CLK a_25419_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12688 _1090_.X a_16219_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12689 vssd1 _1247_.B1 a_1828_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X12690 _1888_.Q a_26267_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12691 vssd1 _1032_.C a_21617_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12692 _1074_.C _1768_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12693 a_15569_17455# a_15299_17821# a_15479_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12694 a_26651_8029# a_25953_7663# a_26394_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12695 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_12355_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12696 a_7105_22717# a_6835_22351# a_7015_22351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12697 vssd1 _1170_.B2 a_2148_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X12698 _1274_.A _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X12699 _0965_.X a_18703_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X12700 a_3993_27497# _1775_.C1 _2004_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12701 _1888_.Q a_26267_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12702 vccd1 a_9644_20871# _1335_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X12703 vccd1 _1941_.CLK a_18243_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12704 a_10938_16341# _2006_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X12705 a_23391_16733# a_23211_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12706 vccd1 _1208_.A1 a_7002_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X12707 a_13441_1685# a_13275_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12708 a_12150_1501# a_11877_1135# a_12065_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12709 vccd1 a_23047_1653# a_22963_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12710 a_8399_4943# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12711 vssd1 _1184_.B1 a_20072_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X12713 a_17415_24640# _1873_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12714 a_16219_22057# _0966_.B1 a_16301_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12716 vssd1 _1254_.A2 a_4247_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X12717 _1179_.B1 a_18459_13131# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X12718 a_17405_12015# _1110_.A a_17323_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12719 a_24757_31599# a_24591_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12721 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12723 _1047_.C a_8454_15797# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X12724 a_24757_8751# a_24591_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12725 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_8477_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X12726 _1150_.A2 a_24887_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12727 a_26873_8751# a_26707_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12728 a_25309_26159# a_25143_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12729 vccd1 _1823_.Q a_23391_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12731 vccd1 a_23691_9019# a_23607_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12732 vccd1 a_22015_11471# _1723_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12733 vssd1 _1337_.S a_4534_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X12734 a_24677_25071# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12735 a_13367_22895# _1868_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12736 a_4571_7119# a_3873_7125# a_4314_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X12737 a_21279_14191# _1975_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X12739 a_27222_16479# a_27054_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12740 _1602_.X a_20676_10499# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12741 vssd1 fanout33.A a_14287_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12742 vssd1 _1282_.A2 a_4253_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X12743 vssd1 a_27755_11293# a_27923_11195# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12744 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12745 vccd1 _0921_.A _0921_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12746 a_17497_20719# _1021_.A a_17415_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12747 vssd1 _1238_.X a_4351_22359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12748 a_22825_18909# a_22291_18543# a_22730_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12749 a_22549_1501# a_22015_1135# a_22454_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12750 vccd1 _1337_.S a_4547_30833# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X12751 vssd1 a_25198_20831# a_25156_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12752 _1849_.CLK a_15794_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X12753 _1059_.X a_15299_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12754 vccd1 fanout24.A a_24499_9301# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12755 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X12756 _1145_.A1 a_8971_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12757 a_12123_24893# _1306_.A2 a_11760_24759# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X12758 a_4859_5162# _1364_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12759 _1112_.B1 a_15391_8320# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12760 a_25800_14025# a_25401_13653# a_25674_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12761 vccd1 a_2750_1653# a_2677_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12762 vssd1 a_18751_5162# _1923_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12763 vccd1 _1033_.A1 a_19194_9411# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12764 a_27241_9117# a_26707_8751# a_27146_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12765 a_1823_19796# _1776_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12766 vccd1 fanout12.A a_7606_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X12767 vssd1 _1873_.CLK a_25235_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12768 a_19053_20175# _1884_.Q a_18969_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12769 vccd1 _0956_.C a_10667_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X12770 a_24201_23817# a_23211_23445# a_24075_23439# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12771 vssd1 a_27038_13215# a_26996_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12774 _1068_.C1 a_14287_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12775 a_17029_29973# a_16863_29973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12777 a_23579_5853# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12778 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12779 _1838_.Q a_22311_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12782 a_25125_7119# a_24591_7125# a_25030_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12783 vccd1 a_25842_4917# a_25769_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12784 _1907_.CLK a_8307_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X12785 a_10506_30511# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12786 vccd1 a_25842_16885# a_25769_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12789 _1665_.A a_15387_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12790 vssd1 a_9282_16341# _1090_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12791 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5639_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12792 vssd1 _0911_.A a_3276_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12794 vssd1 _1055_.C a_13521_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12795 a_2566_25183# a_2398_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12797 a_20437_11471# _1573_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12798 vccd1 _1685_.A_N a_21647_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12799 a_22181_26709# a_22015_26709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12800 a_8392_26159# _1344_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12801 a_10593_22057# _0921_.B a_10951_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12802 vssd1 a_15411_4917# a_15369_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12806 vccd1 a_25106_9269# a_25033_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12807 vccd1 _1723_.A_N a_27167_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12808 vssd1 a_5692_15253# _1291_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X12809 _1979_.Q a_24979_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12810 vssd1 fanout20.X a_25787_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12812 vssd1 _1775_.C1 _1769_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12813 a_4719_16733# _1249_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12814 vccd1 a_23443_9514# _1965_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12815 _1287_.A _1242_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X12816 vccd1 a_20046_31711# a_19973_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12817 a_15795_25615# a_14931_25621# a_15538_25589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12818 vssd1 a_15081_22325# _1116_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
R27 temp1.capload\[13\].cap_43.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X12819 a_2290_13215# a_2122_13469# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X12820 a_10822_25731# _1422_.B a_10740_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12821 a_2639_3855# a_1775_3861# a_2382_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12823 vccd1 _1284_.B1 a_4127_22869# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X12825 vssd1 _1459_.A a_18611_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12826 a_15929_3311# _1610_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12827 vccd1 a_2807_4667# _0913_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12828 vssd1 _1762_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12829 _1073_.X a_16219_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X12830 _1672_.A a_20999_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X12831 a_26183_23439# a_25401_23445# a_26099_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12832 vccd1 fanout20.X a_22015_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12833 vssd1 a_2639_4943# a_2807_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12834 vssd1 a_4035_10901# _1246_.A3 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X12835 vccd1 a_6607_6250# _1783_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12836 vccd1 a_24811_14735# a_24979_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12838 a_12268_9615# _0991_.X a_11777_9269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12839 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_5731_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12840 vccd1 _1221_.A a_2726_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X12841 a_15465_25615# a_14931_25621# a_15370_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12842 vssd1 a_17139_9839# _1293_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12843 a_5416_21781# _1242_.A1 a_5545_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X12844 vccd1 _1744_.B a_17812_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X12845 vssd1 _1153_.A a_19439_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12847 a_19388_8323# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12848 _1125_.X a_6651_11587# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X12849 vssd1 _1269_.A1 a_11403_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X12850 vccd1 a_27215_1300# _1951_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12851 a_16127_6941# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12852 vccd1 a_24039_12559# _1985_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12854 _1137_.X a_18519_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X12855 vssd1 _1047_.C a_17017_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12856 a_4252_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X12857 a_13122_23555# _1422_.B a_13040_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12858 vccd1 a_14563_21807# _0958_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12859 a_24945_7119# _1599_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12860 vccd1 _1975_.Q a_27807_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12862 vccd1 a_4259_13103# _1780_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12863 vssd1 fanout28.A a_9779_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12864 vssd1 a_2382_3829# a_2340_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12865 _1636_.A a_18147_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X12867 vssd1 _1941_.CLK a_22015_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12869 vssd1 _1119_.A1 a_18697_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12870 a_2957_24527# _1769_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12871 vssd1 a_11760_24759# _1352_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X12872 vssd1 a_10073_23737# a_10007_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X12874 vccd1 a_2686_23439# _1763_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12875 a_4709_13647# _1217_.B1 a_5241_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12876 _1128_.B a_25991_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12877 a_25750_3423# a_25582_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12878 a_9779_11791# _1121_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12879 vccd1 a_10167_31029# a_10083_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X12880 vssd1 a_14894_16479# a_14852_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12882 _1102_.B a_22771_5755# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12883 a_16209_16617# _1889_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X12884 a_5428_13109# _0917_.A a_5356_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X12885 a_6743_10703# _1086_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.19825 ps=1.26 w=0.65 l=0.15
X12886 vssd1 a_8822_2741# a_8780_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X12887 a_16649_12015# _1685_.B a_16577_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X12888 a_10873_23805# _0958_.A a_10791_23552# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12889 a_18642_22467# _1484_.B a_18560_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X12890 a_10350_10089# _1008_.X a_10270_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12891 a_5817_10089# _1291_.A1 a_5721_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X12892 a_26203_10602# _1727_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X12893 a_25401_22357# a_25235_22357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12894 a_7828_6351# _1173_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X12896 vssd1 _1084_.C1 a_6559_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X12897 vccd1 _1086_.A a_7019_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12898 a_22361_30511# a_21371_30511# a_22235_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12899 a_3168_24905# a_2769_24533# a_3042_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12900 vccd1 _1053_.A a_13183_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X12901 a_5817_19087# _1234_.A2 _1280_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X12902 vssd1 a_10811_6005# a_10769_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X12903 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12904 vccd1 _0956_.C a_10699_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12905 _1448_.A a_5731_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X12906 _1155_.B a_14287_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X12907 a_6808_31849# a_6559_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X12908 _1879_.Q a_26267_22325# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12910 vccd1 _1148_.B a_6831_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X12911 vssd1 _1907_.CLK a_9135_7125# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12912 a_6564_25071# _1305_.B a_6073_25045# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X12913 a_10765_19407# _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12915 a_25198_17567# a_25030_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12916 vccd1 _0918_.A _1232_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12918 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_6651_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X12919 vssd1 _1763_.A2 a_4534_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X12920 vccd1 _1448_.A a_7387_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12921 a_5354_28335# clkbuf_0_temp1.i_precharge_n.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X12922 a_15512_22351# _0965_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X12923 a_23649_21807# a_22659_21807# a_23523_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X12924 a_26597_17455# a_26431_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12925 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12927 vssd1 a_19487_26922# _1875_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X12928 vccd1 a_22898_18655# a_22825_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12929 a_12282_11177# _1045_.C1 a_12202_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X12930 a_17443_26525# a_16661_26159# a_17359_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X12931 _1879_.Q a_26267_22325# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12932 _1519_.A a_21091_24349# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12933 _1887_.Q a_28015_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12934 a_12299_25437# a_11435_25071# a_12042_25183# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X12935 _1738_.X a_20539_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X12936 a_14545_4949# a_14379_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12937 vccd1 _1139_.C a_9595_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12938 a_15693_12043# _0958_.A a_15607_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X12940 _1521_.A a_20492_20291# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12941 a_4337_1679# _1649_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X12942 vccd1 a_7711_5652# _1565_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12944 _1344_.Y _1344_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12945 a_19487_26922# _1494_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12946 a_2965_20719# _1268_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X12947 vssd1 _1089_.B a_17409_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X12948 vccd1 a_26387_9514# _1678_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12950 vccd1 _1306_.A2 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12951 vssd1 _1141_.C a_17293_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X12952 a_7005_1135# _1755_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12953 vccd1 _1830_.CLK a_20083_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12955 a_27330_28701# a_27057_28335# a_27245_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12956 vccd1 a_10073_23737# a_10103_23478# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X12957 _1776_.X a_6968_21379# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X12958 vccd1 _1544_.A_N a_9043_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12959 vccd1 _1113_.C a_17691_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X12960 a_25033_9295# a_24499_9301# a_24938_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X12961 a_18697_10927# a_18427_11293# a_18607_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X12963 _1250_.A1 _1199_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12964 vssd1 _1833_.Q a_18560_23145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X12965 a_23667_10205# a_23487_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X12966 vccd1 _1474_.A_N a_13275_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12967 a_15377_29423# _1858_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12968 vccd1 _1110_.A a_18243_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12969 _1025_.B a_15227_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12970 vccd1 a_20947_11471# a_21115_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12972 a_19878_1501# a_19605_1135# a_19793_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X12973 fanout28.A a_1591_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X12974 _0973_.B a_27463_6843# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12975 a_9186_13255# _1198_.B2 a_9400_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X12976 vccd1 _1924_.CLK a_22659_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X12977 vccd1 _1768_.A a_9503_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12978 vccd1 a_20407_2986# _1989_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12979 a_6549_9001# _1086_.B a_6467_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X12980 a_4601_12879# _1218_.B _1277_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X12981 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12982 _1834_.Q a_23047_24501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12983 _1031_.X a_14747_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X12984 a_12061_4949# a_11895_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12985 vccd1 _1374_.A_N a_8675_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X12986 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12987 a_13257_20495# _1781_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12988 a_19793_5487# _1942_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12989 vssd1 a_20947_11471# a_21115_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12990 a_25800_24905# a_25401_24533# a_25674_24527# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X12991 a_14733_3855# _1622_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X12992 _1767_.Y _1767_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12993 vssd1 _1907_.CLK a_6283_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X12994 _1834_.Q a_23047_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12995 a_8828_16189# a_8785_15974# a_8756_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X12998 vccd1 _1353_.A a_5271_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12999 vccd1 _1265_.A1 a_5911_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X13000 a_25125_15645# a_24591_15279# a_25030_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13001 a_27295_24349# a_26431_23983# a_27038_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13002 vccd1 a_22311_26427# a_22227_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13003 a_13806_21263# a_13367_21269# a_13721_21263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13004 _1619_.X a_14328_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13005 vssd1 _1828_.Q a_16904_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13008 vccd1 _1242_.A1 a_4248_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13010 a_13621_3145# a_12631_2773# a_13495_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13011 vssd1 a_15411_3829# a_15369_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13012 a_8385_30511# a_8208_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X13013 vccd1 a_17727_29967# a_17895_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13014 vccd1 a_15538_25589# a_15465_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13015 a_9945_6037# a_9779_6037# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13016 a_12705_10383# a_12171_10389# a_12610_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13017 a_8178_12015# _1084_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X13018 a_14441_5487# _1066_.B a_14369_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13019 vccd1 _1141_.C a_15115_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13020 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_17132_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13022 a_2217_23983# a_2051_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13023 a_23224_21807# a_22825_21807# a_23098_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13024 _1265_.A2 _1249_.A1 a_5081_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13025 _1165_.C _1086_.B a_6917_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X13026 a_19912_31433# a_19513_31061# a_19786_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13027 vssd1 a_2991_25339# a_2949_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13030 vccd1 a_2807_3579# _1234_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13031 vccd1 _1066_.B a_17227_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13032 a_8395_7119# a_8215_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13033 a_10593_24233# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13034 a_14829_12015# _1010_.A a_14747_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13035 a_26183_22351# a_25401_22357# a_26099_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13038 _0966_.B1 a_16711_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X13040 _1821_.Q a_19735_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13041 vccd1 _1448_.A a_4259_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X13042 a_21533_2223# a_20543_2223# a_21407_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13044 _1110_.A a_14103_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13045 a_20161_32143# _1896_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13046 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13047 _1068_.D1 a_11711_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X13048 vccd1 a_20959_26922# _1903_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13049 vccd1 _1053_.A a_14655_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13050 _1771_.B a_2471_22869# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13051 a_9503_16911# _1269_.A1 a_9921_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13052 vccd1 _1859_.Q a_7383_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13053 vssd1 _1876_.CLK a_22015_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13054 vccd1 _1843_.Q a_17996_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X13055 a_19521_8751# _1153_.A a_19439_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13056 a_11601_25071# a_11435_25071# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13057 vssd1 a_22419_31965# a_22587_31867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13058 temp1.inv2_2.A a_2686_26703# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13059 a_1769_20719# _1282_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X13060 vccd1 a_23266_4917# a_23193_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13061 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13062 vssd1 a_9613_22869# a_9547_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X13063 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X13064 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_7387_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13065 a_5271_26409# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13067 vssd1 _0953_.C1 a_19807_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13068 vssd1 a_11030_3423# a_10988_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13069 vssd1 _1184_.C1 a_19439_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13070 _1108_.C1 a_11711_14848# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X13071 _1794_.Y _1316_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13072 vccd1 fanout20.X a_25235_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13073 vccd1 _1074_.C a_14319_7691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13074 a_5639_26703# _1764_.B _1762_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13076 _1752_.X a_7659_8029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X13077 a_22764_20553# a_22365_20181# a_22638_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13079 a_9999_4765# a_9301_4399# a_9742_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13080 vssd1 _1141_.C a_12049_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13081 a_13875_23658# _1421_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13082 vssd1 a_20315_25834# _1893_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13083 a_17861_32143# _1841_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13084 vssd1 _1113_.C a_19593_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13085 vccd1 a_15151_10205# a_15319_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13086 vccd1 _1132_.C a_14839_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13087 a_20758_12265# _1577_.B a_20676_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13088 a_24769_30287# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13089 vssd1 a_11711_27791# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13091 vccd1 a_17159_9019# a_17075_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13092 vssd1 a_26267_22325# a_26225_22729# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13093 vssd1 _1008_.A a_14839_10499# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X13095 vccd1 a_1641_13879# _1230_.A4 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X13097 _1534_.A a_17548_25321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13098 a_25029_19465# a_24039_19093# a_24903_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13099 vssd1 fanout20.X a_24591_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13100 vccd1 _2023_.CLK a_1775_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13101 _1760_.A_N a_2807_28603# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13102 vccd1 _1875_.Q a_19562_25321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X13104 vssd1 a_2807_4667# _0913_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13105 a_25769_26703# a_25235_26709# a_25674_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13106 a_4441_26159# _1273_.A1 _1769_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13107 vccd1 _1882_.CLK a_23671_21269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13108 _1020_.D1 a_15483_13760# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X13109 vccd1 a_20131_6250# _1745_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13111 a_16156_7913# _1071_.B1 a_16054_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X13112 vccd1 a_11858_17973# _1133_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X13114 a_27238_21085# a_26965_20719# a_27153_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13116 vccd1 _1685_.A_N a_22015_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13117 a_25198_6687# a_25030_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13118 vssd1 a_20046_5599# a_20004_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13119 a_12042_25183# a_11874_25437# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13120 _1549_.A a_9223_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X13121 a_25566_8181# a_25398_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13122 a_18072_32521# a_17673_32149# a_17946_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13124 _1700_.X a_28083_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13125 a_19268_15113# a_18869_14741# a_19142_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13126 a_15657_19881# _0984_.X a_15575_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X13127 a_6808_30761# a_6559_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X13128 vccd1 a_24535_21263# a_24703_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13129 a_9200_26703# a_8951_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X13130 a_12801_25615# _1901_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13131 a_2198_8181# a_2030_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13132 a_7564_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13133 vssd1 _1841_.CLK a_15023_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13134 vssd1 _2023_.CLK a_1775_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13135 vssd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_15750_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13139 _1180_.X a_14931_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13141 vssd1 a_24535_21263# a_24703_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13142 _1861_.Q a_15963_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13144 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_13183_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13145 vssd1 _1231_.B2 a_3249_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13146 vssd1 a_22235_30877# a_22403_30779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13147 vssd1 a_22863_29691# a_22821_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13148 _1761_.X a_27167_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13149 vssd1 a_21575_23163# a_21533_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13150 _0961_.A a_15299_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13151 a_16623_2589# a_15759_2223# a_16366_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13152 a_14545_3861# a_14379_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13153 vssd1 _1438_.B a_12349_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13154 a_23941_31375# temp1.capload\[6\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13155 vccd1 _1316_.X a_7189_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X13156 vccd1 _1021_.A a_17415_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13158 a_25539_1501# a_24757_1135# a_25455_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13159 vssd1 _1065_.B a_22285_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13160 _1861_.Q a_15963_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13161 a_25455_27613# a_24757_27247# a_25198_27359# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13162 vssd1 a_12587_14954# _1850_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13163 _1607_.X a_18468_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13164 a_13725_22717# _0964_.A a_13643_22464# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13165 vssd1 _1344_.B a_5271_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13166 _1427_.A a_18239_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X13167 _1102_.B a_22771_5755# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13168 vccd1 a_2686_10383# _2023_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13171 vssd1 _2023_.CLK a_1591_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13172 _1070_.A2 a_16711_15307# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X13173 _1801_.Y _1267_.A1 a_13821_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13174 a_6829_29199# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13175 vssd1 _1882_.CLK a_26431_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13176 vccd1 a_10627_22325# a_10543_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13177 a_5061_23439# _1308_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13179 a_25474_11039# a_25306_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13180 a_1828_19061# _1270_.A a_2220_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X13181 a_11269_16600# _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X13182 vccd1 a_25198_15391# a_25125_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13183 a_25198_31711# a_25030_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13184 a_9258_19881# _1422_.B a_9176_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13185 a_12587_14954# _1441_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13186 _1040_.X a_17691_8320# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X13187 a_27590_27359# a_27422_27613# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13189 vssd1 _1024_.A2 a_16760_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X13190 vssd1 a_6607_6250# _1783_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13193 a_18850_3829# a_18682_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13194 a_16064_11471# _1071_.B1 a_15962_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X13195 a_8955_11791# _1120_.X a_8818_11703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X13196 vccd1 a_26175_10107# a_26091_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13197 _1486_.B a_20563_30779# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13199 a_6261_2223# a_5271_2223# a_6135_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13200 a_20782_4511# a_20614_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13201 a_10969_18543# a_10699_18543# a_10865_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13202 vssd1 a_27847_27613# a_28015_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13203 a_22603_5853# a_21905_5487# a_22346_5599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13204 _1523_.A a_19388_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13205 vssd1 _1762_.A a_7360_15095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X13206 vccd1 a_12778_10357# a_12705_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13208 a_2547_8029# a_1683_7663# a_2290_7775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13209 _1857_.Q a_13755_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13210 a_24853_9295# _1678_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13211 a_11115_7828# _1614_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13212 vssd1 a_7111_25071# _1242_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13213 vccd1 a_27038_24095# a_26965_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13214 _1764_.B a_1766_26159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13216 vccd1 _1198_.A1 a_9601_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X13217 _1007_.X a_19991_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X13218 a_20982_2589# a_20709_2223# a_20897_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13219 vccd1 a_2807_3829# a_2723_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13220 vccd1 _1763_.A2 a_2408_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13221 vccd1 _0964_.A a_11711_14848# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13222 vccd1 a_4495_11989# _1217_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X13223 _1374_.A_N a_7571_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13224 vccd1 _1075_.C a_21127_12897# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13225 _1642_.X a_14328_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13227 a_23193_4943# a_22659_4949# a_23098_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13228 a_24109_8585# a_23119_8213# a_23983_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13229 vccd1 _1459_.A a_15207_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X13230 vssd1 _1857_.Q a_10740_25731# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13231 a_25581_13103# a_24591_13103# a_25455_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13232 vccd1 a_17727_1679# a_17895_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13233 a_3983_28585# _1764_.B _1764_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13237 vssd1 _1177_.Y a_2121_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X13240 _1607_.B a_9135_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X13242 vssd1 a_23691_4917# a_23649_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13244 vssd1 _1448_.A a_4259_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13247 vccd1 _1098_.B a_16307_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13248 vssd1 a_17470_29941# a_17428_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13249 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13360_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13250 vssd1 _1210_.B a_5389_9633# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X13251 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13252 a_1757_2223# a_1591_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13253 a_4061_7119# _2020_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13254 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_16955_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13255 a_6682_7913# _1809_.B a_6600_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13256 vccd1 _1207_.B1_N a_2696_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X13257 _1156_.Y _1156_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13259 _1616_.A a_9683_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13260 a_20138_30623# a_19970_30877# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13261 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.LO a_17139_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13262 a_1857_12265# _1219_.A2 a_1775_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13263 a_24535_21263# a_23671_21269# a_24278_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13264 a_7015_19881# _1325_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13265 vssd1 _1195_.B2 a_20629_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13266 a_14453_8207# _1440_.B a_14369_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13267 vccd1 _1123_.X a_6901_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X13268 vccd1 a_12631_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X13270 _0966_.A2 a_18367_25099# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X13271 _0973_.B a_27463_6843# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13272 a_5731_20541# _1242_.A1 a_5625_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X13273 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13276 a_11159_14191# _1846_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13277 a_4333_1135# a_4167_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13279 vccd1 _1855_.CLK a_14287_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13281 a_2686_23439# clkbuf_1_1__f__0380_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X13282 _1116_.B1 a_17231_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X13284 vccd1 a_23155_18909# a_23323_18811# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13285 a_18850_3829# a_18682_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13286 a_11793_6031# _0988_.X a_11877_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13287 a_5639_21807# _0911_.A a_5545_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X13288 vccd1 a_3578_2741# a_3505_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13289 a_20819_4943# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X13290 a_15479_17821# a_15299_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13292 a_7295_6031# _1173_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13293 _0903_.C a_5639_10089# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X13294 a_10643_29967# a_9945_29973# a_10386_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13295 a_21235_25834# _1513_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13298 vccd1 _1801_.Y a_4163_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X13299 a_23487_10205# _1723_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X13300 a_22645_18543# _1393_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13301 a_14821_10205# a_14287_9839# a_14726_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13302 a_17857_28879# a_17323_28885# a_17762_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13303 a_12973_10089# _1069_.B a_12901_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13304 vssd1 _1321_.C a_5701_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13305 _1749_.A a_17319_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13306 a_1814_11177# _1263_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X13307 vssd1 a_10506_30511# temp1.capload\[15\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13309 vccd1 a_26387_1898# _1651_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13310 vssd1 a_13882_1653# a_13840_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13312 a_5080_29423# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13313 vccd1 a_24639_4564# _1959_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13314 a_18597_2767# _1938_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13315 _1842_.Q a_22587_31867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13317 vssd1 _1685_.B a_23849_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13319 vssd1 a_13755_29941# a_13713_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13320 a_22730_27791# a_22457_27797# a_22645_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13321 _1054_.C a_12061_19087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X13322 vccd1 a_16083_17130# _1822_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13323 a_22063_9514# _1577_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13324 a_5086_24893# _1261_.A1 a_4587_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X13327 a_27847_12381# a_26983_12015# a_27590_12127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13328 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI a_9200_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X13329 vccd1 _1317_.X a_5908_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X13331 vccd1 a_19487_11690# _1586_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13332 vccd1 a_27859_30676# _1450_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13333 a_8569_2767# _1614_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13334 a_23266_2335# a_23098_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13335 _0989_.A2 a_3175_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13336 vssd1 a_19275_2741# a_19233_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13337 vccd1 a_8177_12533# _1123_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X13338 a_1857_12265# _1208_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X13339 _2004_.Q a_3635_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13340 a_17485_18543# _1832_.Q a_17139_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X13341 vssd1 _1762_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13342 vccd1 _1199_.X a_12927_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X13343 vccd1 _1924_.CLK a_24959_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13344 vccd1 a_2696_11177# _1219_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13345 a_18637_11809# _1127_.A a_18551_11809# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13346 vssd1 a_21511_28500# _1870_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13347 vccd1 a_16531_24349# a_16699_24251# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13348 a_22645_23983# _1832_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13349 a_17477_12015# _1098_.B a_17405_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13350 a_19470_22467# _1405_.B a_19388_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13351 a_12149_6351# _1145_.A1 a_11711_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13353 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13354 vssd1 a_21187_9295# _1685_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13355 a_19487_11690# _1586_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13357 vssd1 _1353_.A _1342_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13358 a_22269_26159# a_21279_26159# a_22143_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13359 _1652_.X a_3748_3971# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13360 a_25309_3311# a_25143_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13363 a_22195_15823# a_22015_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13364 a_12701_11849# a_11711_11477# a_12575_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13365 _1880_.Q a_26175_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13366 _1509_.A a_20308_21379# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13368 vssd1 _2023_.CLK a_1775_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13369 a_17569_20719# _1876_.Q a_17497_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13370 a_5710_2589# a_5437_2223# a_5625_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13372 vssd1 a_16911_31274# _1896_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13373 a_11138_31965# a_10699_31599# a_11053_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13375 vccd1 _1464_.B a_9775_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13376 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_7479_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13378 a_16301_21807# _1898_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X13379 a_24110_21263# a_23837_21269# a_24025_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13380 vccd1 a_26099_6031# a_26267_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13381 vccd1 a_1828_14709# _1311_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X13382 _1084_.B1 a_9176_10089# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13383 vssd1 a_18003_29789# a_18171_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13384 vccd1 _1823_.CLK a_26983_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13385 a_24945_6575# _1605_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13388 a_7809_18517# _0925_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X13389 a_11940_9615# _1139_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X13390 a_16106_24349# a_15667_23983# a_16021_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13391 a_12318_8181# a_12150_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13392 vssd1 fanout33.A a_16863_27797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13393 _1267_.B2 _1234_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13394 vssd1 a_2382_3423# a_2340_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13395 a_11907_20175# _2004_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X13396 vssd1 _1149_.C1 a_14287_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13397 vssd1 a_20407_24746# _1837_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13398 vssd1 _1890_.Q a_19480_17705# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13399 vssd1 fanout20.X a_22015_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13400 vccd1 a_18751_21972# _1877_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13401 vccd1 a_22063_18218# _1527_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13403 a_6953_8545# _1165_.A a_6867_8545# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13404 a_2769_22057# _1237_.B2 a_2685_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13406 a_27149_9839# a_26983_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13407 a_25030_5853# a_24591_5487# a_24945_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13408 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13409 vccd1 _1685_.A_N a_21463_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13410 a_14726_30877# a_14287_30511# a_14641_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13411 _1074_.C a_9195_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13412 a_20341_4399# a_20175_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13413 a_15081_12533# _1103_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X13414 a_19954_31029# a_19786_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13415 vssd1 a_17831_30676# _1471_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13417 vccd1 a_2455_8207# a_2623_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13419 vssd1 a_23707_29967# a_23875_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13421 a_10386_1653# a_10218_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13422 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13423 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_15483_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13425 a_24209_25615# _1837_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13426 vccd1 _0913_.A1 a_5455_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X13428 a_23377_16917# a_23211_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13429 _1355_.X a_5404_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13430 a_4519_9991# _1298_.A1 a_4753_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X13431 a_27422_12381# a_27149_12015# a_27337_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13432 a_20897_22895# _1829_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13433 vssd1 a_16991_9117# a_17159_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13434 vccd1 _1818_.Q a_8855_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13435 a_14453_9839# a_14287_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13437 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X13438 vccd1 _0909_.A a_6559_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13439 a_17946_1501# a_17507_1135# a_17861_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13440 vssd1 a_13047_12180# _1911_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13441 a_23649_3311# a_22659_3311# a_23523_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13443 vccd1 _1857_.Q a_10822_25731# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X13444 vssd1 a_8447_20884# _1433_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
R28 temp1.capload\[8\].cap_53.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X13446 a_14825_2767# _1934_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13447 vccd1 a_8447_7828# _1751_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13448 _1403_.B a_24243_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13449 a_23799_3855# a_23101_3861# a_23542_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13450 a_3505_2767# a_2971_2773# a_3410_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13451 a_16623_2589# a_15925_2223# a_16366_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13452 vccd1 _1110_.A a_15391_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13453 a_12150_13647# a_11711_13653# a_12065_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13454 _1675_.X a_22563_8029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13455 a_15496_32521# a_15097_32149# a_15370_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13458 a_21032_15823# _1020_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X13459 a_7699_3855# a_7001_3861# a_7442_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13460 a_13047_12180# _1569_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13462 a_8447_20884# _1433_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13463 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13464 a_16159_20747# _1053_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13465 a_2765_6409# a_1775_6037# a_2639_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13466 a_4988_32463# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13467 a_18409_2773# a_18243_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13468 _1598_.X a_19112_9411# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13469 vccd1 _1304_.B a_6277_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X13471 a_7975_2589# a_7111_2223# a_7718_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13472 vssd1 a_20131_6250# _1745_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13474 _1893_.Q a_23691_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13475 vccd1 _1844_.Q a_13122_23555# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X13476 _1247_.B1 _1246_.B2 a_3329_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.105 ps=1.21 w=1 l=0.15
X13477 vssd1 a_25807_3829# a_25765_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13479 a_5878_2335# a_5710_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13480 vssd1 a_13783_5162# _1610_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13481 vccd1 a_14894_9951# a_14821_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13482 vssd1 fanout12.A a_8307_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13484 a_9284_21781# a_9135_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13485 a_26601_14191# _1984_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13486 vccd1 _1073_.A2 a_17305_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X13489 a_16711_22923# _0961_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13490 _1321_.C a_3707_6144# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X13491 a_22730_27791# a_22291_27797# a_22645_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13492 vccd1 _1972_.Q a_16064_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X13493 a_10643_1679# a_9945_1685# a_10386_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13494 vssd1 _1882_.Q a_20768_22057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13495 vccd1 _1974_.Q a_22238_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X13496 _1197_.B a_10515_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X13497 a_17538_7913# _1577_.B a_17456_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13498 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_8158_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X13499 vccd1 a_10349_25045# a_10379_25398# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13500 a_14467_14557# a_14287_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13501 vssd1 a_21575_2491# a_21533_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13503 a_11877_8213# a_11711_8213# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13504 a_26597_17455# a_26431_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13505 vssd1 a_25455_13469# a_25623_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13506 vssd1 fanout21.X a_26707_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13507 a_8945_8573# a_8675_8207# a_8855_8207# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
R29 temp1.capload\[5\].cap_50.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X13508 a_17017_21629# _1838_.Q a_16945_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13509 a_20867_8426# _1598_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13510 a_2581_9673# a_1591_9301# a_2455_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13511 a_25030_27613# a_24757_27247# a_24945_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13512 a_20584_20969# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13513 _1662_.X a_12535_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13514 a_5487_5281# _1255_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13515 _0965_.B1 a_17539_22923# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X13516 a_27847_19997# a_27149_19631# a_27590_19743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13517 a_10945_23805# _1855_.Q a_10873_23805# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13518 vccd1 _1132_.A a_15483_23552# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13519 a_11934_9295# _1436_.B a_11777_9269# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13520 vccd1 a_11023_31274# _1868_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13521 a_24972_18377# a_24573_18005# a_24846_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13522 a_5889_10089# _1281_.A1 a_5817_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13524 _1855_.CLK a_11711_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13526 vccd1 _0918_.A a_9135_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X13527 vccd1 _0964_.A a_17231_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13528 a_7469_8751# _1279_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13529 a_27498_11039# a_27330_11293# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13531 a_17102_31711# a_16934_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13532 a_4627_13967# _1217_.A2 a_4877_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13533 vccd1 a_26099_23439# a_26267_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13534 _1645_.A a_14651_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13535 a_21235_1898# _1738_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13536 a_3748_3971# _1448_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13537 a_25539_24349# a_24757_23983# a_25455_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13538 _1873_.CLK a_22567_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X13541 vssd1 _1768_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13542 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_8215_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13543 a_13122_14441# _1038_.D1 a_12873_14337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X13544 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_8477_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13545 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13546 a_22155_23658# _1691_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13547 vccd1 _1896_.CLK a_19439_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13549 a_25953_18909# a_25419_18543# a_25858_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13550 vssd1 a_26099_23439# a_26267_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13551 a_19069_12879# _1090_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X13552 vccd1 a_3210_27765# a_3137_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X13553 vssd1 _1243_.A a_6564_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X13554 vssd1 a_4220_21959# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X13555 a_9779_11471# _1120_.X _1122_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13556 a_4252_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13557 _1270_.A _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13559 vssd1 a_12978_27791# a_13084_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13560 a_15473_8573# _1110_.A a_15391_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13561 vssd1 a_28015_10107# a_27973_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13563 vccd1 a_12321_22325# _1142_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X13567 vccd1 _1132_.A a_17415_24640# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13568 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13570 a_12532_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13571 _1181_.X a_15667_24527# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X13572 vssd1 _0913_.Y temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13573 a_21463_15279# _1976_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13574 a_19973_1501# a_19439_1135# a_19878_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13576 a_26141_7663# _1982_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13577 vssd1 _0913_.A1 a_5731_20541# vssd1 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X13578 a_10589_3311# a_10423_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13579 vssd1 _1840_.Q a_12488_26409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13581 a_25589_22351# _1879_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13582 a_10218_8207# a_9945_8213# a_10133_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13583 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13584 vccd1 a_10471_7828# _1813_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13585 a_3873_11791# _1177_.B a_3789_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X13587 vccd1 a_16791_2491# a_16707_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13588 a_17302_1679# a_16863_1685# a_17217_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13589 vssd1 _1274_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X13590 vccd1 _0961_.A a_13367_22895# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13591 a_15933_22895# _1053_.A a_15851_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13593 vccd1 a_26479_1300# _1616_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13594 a_1941_7125# a_1775_7125# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13595 vccd1 _1277_.A a_3063_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13596 _1999_.CLK a_6283_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X13598 vssd1 _1325_.A2 a_5720_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X13599 a_8209_15529# _1313_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X13600 _1198_.A2 a_9779_12015# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X13601 vccd1 fanout37.A a_18703_18005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13602 a_24830_15797# a_24662_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13603 a_9142_15101# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X13604 vccd1 a_24639_14356# _1984_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13605 _1517_.A a_20584_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13606 vssd1 _1768_.A a_8307_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13607 vssd1 _1032_.C a_21433_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X13608 a_8546_1653# a_8378_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13609 vssd1 _2023_.CLK a_1683_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13610 vssd1 a_12502_4917# a_12460_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13611 vssd1 fanout24.A a_25143_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13613 a_24159_16911# a_23377_16917# a_24075_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13614 vccd1 a_16290_4399# a_16396_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X13615 vccd1 a_3299_22325# _1240_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X13617 a_2129_4943# _2021_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13618 a_17113_11177# _1155_.B a_17041_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X13619 vssd1 _1999_.CLK a_10423_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13622 a_4035_23957# _1304_.B a_4262_24305# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X13623 a_11711_21263# _0984_.B1 a_11793_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13624 a_6463_14441# _1810_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13625 vssd1 _0918_.A a_9135_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X13626 a_17841_17601# _1049_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13627 a_23443_31764# _1474_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13628 a_25283_14356# _1706_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13629 a_8392_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13630 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z _1243_.Y a_8392_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13631 _1768_.A a_6835_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13633 vccd1 a_24887_25589# a_24803_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13634 vccd1 _1032_.C a_21463_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13635 _1405_.B a_17047_17455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X13636 a_25156_5487# a_24757_5487# a_25030_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13637 a_25455_6941# a_24591_6575# a_25198_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13639 vccd1 a_2715_7931# a_2631_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13640 a_17313_19453# _0964_.A a_17231_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13641 a_3152_18543# _1300_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X13643 vssd1 a_12318_8181# a_12276_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13644 a_2769_24533# a_2603_24533# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13645 a_24941_3861# a_24775_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13646 a_4338_20969# _1282_.A2 a_4035_20693# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X13647 vssd1 _0987_.B _1071_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13648 vssd1 _1146_.B a_14328_3561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13649 a_3276_20495# _1282_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13650 a_7002_5263# _1202_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13651 a_26226_8029# a_25787_7663# a_26141_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13652 vssd1 _1242_.B1 a_6099_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13653 a_17853_18377# a_16863_18005# a_17727_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13654 a_3091_1679# a_2309_1685# a_3007_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13655 vssd1 _1876_.CLK a_22015_26709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13656 a_10951_22057# _0921_.B a_10593_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13657 a_23098_11293# a_22825_10927# a_23013_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13658 vccd1 _1143_.A a_14905_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X13659 vccd1 a_9275_10602# _1561_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13661 a_27697_8751# a_26707_8751# a_27571_9117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13662 vccd1 _1941_.CLK a_19439_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13663 a_15512_12559# _1100_.X a_15410_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X13664 a_7561_17277# _1768_.A a_7479_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X13666 vssd1 a_17102_26271# a_17060_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13667 vssd1 _1301_.A1 a_3247_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X13668 a_15496_25993# a_15097_25621# a_15370_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13669 vssd1 a_11759_1898# _1956_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13670 a_17497_24893# _1132_.A a_17415_24640# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13671 vccd1 _1328_.S a_5047_21237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X13672 vccd1 _1690_.A_N a_21923_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13673 a_26183_4943# a_25401_4949# a_26099_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13674 vssd1 _1907_.CLK a_9779_6037# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13675 vssd1 a_23167_14954# _1985_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13676 vssd1 a_7683_1403# a_7641_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13677 a_2198_1247# a_2030_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13678 a_15185_7497# a_14195_7125# a_15059_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13679 vccd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13680 _1074_.C _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X13682 a_2649_23047# _1763_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X13683 a_1643_21781# _1775_.A2 a_1925_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X13684 a_23903_24746# _1507_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13685 a_26099_23439# a_25235_23445# a_25842_23413# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13686 vccd1 _1878_.Q a_20079_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13687 vccd1 a_7479_17277# _1139_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X13688 vccd1 a_14345_15425# _1095_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X13689 vccd1 _1744_.A_N a_22015_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13690 a_4146_7119# a_3707_7125# a_4061_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13691 vssd1 a_20315_26922# _1895_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13692 a_10279_16911# a_10667_16885# _1141_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13693 a_27238_15645# a_26799_15279# a_27153_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13694 vccd1 _1242_.B1 a_4526_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X13696 vssd1 _1813_.Q a_8215_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13697 a_9681_10927# a_9411_11293# a_9591_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X13698 a_15207_1679# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X13699 a_11877_13653# a_11711_13653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13700 vssd1 a_9284_21781# _1282_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X13701 a_21695_19796# _1393_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13702 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13703 a_23167_14954# _1723_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13704 vssd1 a_6056_20871# _1328_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13707 _1985_.CLK a_24039_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13708 _1368_.X a_5588_6825# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13709 a_8464_28879# a_8215_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X13710 vccd1 _0952_.A1 a_9687_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13712 a_20387_5853# a_19605_5487# a_20303_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13713 a_21235_31274# _1486_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13714 vssd1 _1208_.A1 a_6644_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13715 a_2765_5321# a_1775_4949# a_2639_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13717 io_out[1] a_1643_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13718 a_25566_8181# a_25398_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13719 vccd1 a_23047_26677# a_22963_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13720 _1824_.Q a_27647_16635# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13722 a_14345_15425# _1094_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X13723 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13724 a_24757_23983# a_24591_23983# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13726 a_11138_31965# a_10865_31599# a_11053_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13727 a_18272_17705# _1184_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X13728 vccd1 a_23691_27515# a_23607_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13730 vccd1 a_9828_26935# _1329_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X13731 a_12907_18543# _1845_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13732 vssd1 _2005_.Q a_11969_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X13733 a_24205_19093# a_24039_19093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13735 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13736 _2003_.Q a_3083_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13737 a_5231_22869# _1306_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X13738 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_12263_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X13739 vssd1 a_5354_28335# temp1.dcdc.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X13741 a_1643_21781# _1240_.X a_1841_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X13745 vccd1 _1882_.CLK a_25235_22357# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13746 a_16665_25071# a_16488_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X13747 vccd1 _1032_.C a_20267_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13750 _1195_.B2 a_23967_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13751 a_9742_5599# a_9574_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13753 _1068_.A1 a_15503_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13755 _1083_.A a_7867_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13756 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13757 vccd1 _0965_.A2 a_15013_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13758 a_23565_23439# _1892_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13759 a_24201_17289# a_23211_16917# a_24075_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13760 vccd1 a_8654_29967# a_8760_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X13761 vccd1 a_26099_22351# a_26267_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13762 a_8669_5309# a_8399_4943# a_8579_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X13763 _1853_.Q a_15319_30779# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13765 _0930_.A a_6559_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X13766 a_10777_27247# _1555_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13768 vssd1 a_4035_30485# _1330_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X13769 vccd1 a_12771_3476# _1624_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13770 vccd1 _1843_.Q a_18239_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13772 a_17359_26525# a_16495_26159# a_17102_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13773 vccd1 _1685_.A_N a_22383_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13774 a_12065_29423# _1902_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13775 vssd1 a_26099_22351# a_26267_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13778 a_5912_15279# _1289_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X13779 vssd1 a_16182_3423# a_16140_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13780 vssd1 a_3801_28981# _0909_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X13781 vssd1 a_1643_21237# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13782 a_25401_16917# a_25235_16917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13783 _0909_.B a_6600_24233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13784 _1139_.C a_7479_17277# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X13785 a_17428_2057# a_17029_1685# a_17302_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13786 _1149_.A1 a_23047_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13787 a_23009_29973# a_22843_29973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13788 _1081_.D1 a_18151_10496# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X13789 a_9442_3971# _1607_.B a_9360_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13790 vssd1 a_12759_4943# a_12927_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13791 vccd1 a_10938_16341# _1075_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X13792 a_2581_2223# a_1591_2223# a_2455_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13795 _1122_.A1 _1198_.A2 a_10227_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X13797 vssd1 _1033_.A2 a_20429_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X13798 a_10094_4943# _0989_.B2 a_9937_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X13800 _1385_.A a_20860_19203# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13801 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13802 vssd1 _1855_.CLK a_13459_24533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13804 _1528_.A a_26267_16885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13805 a_26965_13469# a_26431_13103# a_26870_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13806 _1171_.Y _1162_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13807 a_22879_25615# a_22181_25621# a_22622_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13808 a_21327_1300# _1734_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13809 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_3063_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X13810 _1364_.X a_8855_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13811 vssd1 a_22622_31029# a_22580_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13812 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13813 a_13797_22717# _1899_.Q a_13725_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X13815 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13817 a_22454_25615# a_22015_25621# a_22369_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13818 a_23005_1135# a_22015_1135# a_22879_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13819 a_15614_6031# _0952_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X13822 _0939_.A a_16863_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X13823 a_14323_24527# a_13459_24533# a_14066_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13826 vccd1 a_27755_28701# a_27923_28603# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13827 a_15633_19061# _1020_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X13828 vssd1 _1011_.A1 a_7933_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13830 vssd1 a_17573_4917# _1155_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X13831 a_23849_5487# a_23579_5853# a_23759_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X13832 a_19562_11177# _1577_.B a_19480_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13833 a_10515_19407# _0929_.A _0930_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13834 vssd1 a_25198_5599# a_25156_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X13835 _1878_.Q a_27831_22075# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13836 a_9503_16911# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13838 a_14471_6575# _1063_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13839 a_14894_30623# a_14726_30877# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13840 vccd1 a_2991_25339# a_2907_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13841 vccd1 _1424_.A_N a_19439_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13842 a_25198_15391# a_25030_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13843 _1019_.B a_21575_7931# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13844 vccd1 a_22879_24527# a_23047_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13845 _1140_.C a_7442_17429# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13846 _1324_.A _1034_.Y a_8118_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X13847 vccd1 temp1.capload\[6\].cap_51.LO temp1.capload\[6\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13848 vccd1 a_12575_29789# a_12743_29691# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13849 vssd1 a_12689_6721# _1069_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X13850 a_26352_7663# a_25953_7663# a_26226_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13852 a_13367_16367# _1840_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X13853 a_7185_4399# a_7019_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13854 a_9301_4399# a_9135_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13856 a_25639_16733# a_24941_16367# a_25382_16479# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13857 a_7883_4765# a_7019_4399# a_7626_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13858 a_4337_25071# _2007_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13859 a_13490_3561# _1607_.B a_13408_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X13860 vssd1 a_22879_24527# a_23047_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13862 vssd1 a_3983_3311# _1816_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13864 a_25214_16733# a_24775_16367# a_25129_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13866 a_6559_12559# _1255_.A1 a_6981_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13867 a_9912_13763# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13868 a_22081_13621# _0952_.A1 a_22334_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X13870 a_14986_3829# a_14818_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13871 a_8447_6740# _1359_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13872 a_17029_1685# a_16863_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13873 a_19803_7119# a_19623_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X13874 a_14641_9839# _1571_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13875 a_4333_1135# a_4167_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13876 vccd1 _1841_.CLK a_19623_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13878 vccd1 a_23523_11293# a_23691_11195# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X13879 vccd1 clkbuf_0_temp1.i_precharge_n.X a_5354_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13880 _1838_.Q a_22311_26427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13881 vccd1 _1690_.A_N a_22935_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13882 vccd1 a_11299_11092# _1439_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13883 a_9700_31433# a_9301_31061# a_9574_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13884 a_24823_28010# _1551_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13885 vccd1 _1140_.C a_14379_20719# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13886 a_3240_32463# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13887 _1658_.X a_10327_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X13888 vssd1 _1063_.B a_14741_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X13889 a_25582_10205# a_25309_9839# a_25497_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13890 _1538_.A a_15800_26819# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X13891 vccd1 _1188_.B a_4531_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13892 a_4272_7497# a_3873_7125# a_4146_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13893 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_8464_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X13894 a_17565_24129# _1133_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X13895 vccd1 _1132_.C a_15883_13131# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13896 _1744_.B a_25623_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13897 a_2214_4765# a_1941_4399# a_2129_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13898 a_10202_29535# a_10034_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13899 _1459_.A a_12815_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X13901 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13902 a_14821_30877# a_14287_30511# a_14726_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13903 vccd1 a_20591_1898# _1940_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13904 _1261_.A2 a_8615_25953# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X13906 vccd1 _0918_.A a_10593_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13907 _1148_.B a_10167_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13908 vccd1 _1041_.A1 a_16156_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X13909 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13910 a_26099_22351# a_25235_22357# a_25842_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13911 a_12759_15645# a_12061_15279# a_12502_15391# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13912 a_17923_26922# _1461_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13914 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13915 a_12973_5461# _1293_.A1 a_13226_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X13916 a_12613_25621# a_12447_25621# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13917 a_12334_15645# a_11895_15279# a_12249_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X13918 vssd1 _1982_.CLK a_26983_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13919 vccd1 _1177_.B a_3979_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X13920 _1035_.X a_13367_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X13921 a_12383_2589# a_11601_2223# a_12299_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13922 a_9183_12180# _1570_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13923 vssd1 _1855_.CLK a_11435_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13924 a_11023_16042# _1371_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13925 a_7718_2335# a_7550_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13926 vccd1 a_16175_9514# input3.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X13928 vssd1 _1304_.B a_6324_13353# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X13929 a_19057_1679# _1643_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X13930 a_9669_7119# a_9135_7125# a_9574_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13931 a_2970_22895# _1286_.A1 a_2471_22869# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X13932 vccd1 _1390_.B a_22195_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X13933 vssd1 _2023_.CLK a_1775_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X13934 vccd1 _1882_.CLK a_23211_23445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X13935 a_25271_17999# a_24407_18005# a_25014_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X13936 a_1757_6575# a_1591_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13937 a_4248_26409# _1769_.B1 a_3993_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13938 a_12253_24233# _0983_.X a_12171_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13939 a_2248_13103# a_1849_13103# a_2122_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X13941 _1976_.Q a_25439_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13942 vccd1 a_9135_3311# _1607_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13943 a_13599_1300# _1645_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X13944 vccd1 a_5354_28335# temp1.dcdc.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13945 a_24895_14735# a_24113_14741# a_24811_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13946 a_1945_1135# _1808_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X13947 a_24639_12180# _1709_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13948 vssd1 a_25467_28010# _1856_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13950 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13951 a_26183_16911# a_25401_16917# a_26099_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13952 vccd1 _1202_.Y a_7002_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13953 _0991_.X a_15607_12043# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X13954 a_8113_25117# _0911_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X13957 a_5816_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X13959 vccd1 _1801_.B a_3707_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X13960 vssd1 a_2594_31055# clkbuf_0_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13961 vssd1 a_21235_25236# _1883_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X13962 vssd1 a_12500_15797# _1071_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X13963 a_25857_10927# a_24867_10927# a_25731_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X13964 a_13901_21263# a_13367_21269# a_13806_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X13966 vccd1 _1141_.C a_18459_13131# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X13967 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_6736_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13968 vccd1 a_2309_29789# _1760_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X13969 vccd1 a_15750_28335# temp1.capload\[6\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13970 a_2382_28447# a_2214_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13971 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_11711_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X13976 a_25467_28010# _1453_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X13977 a_4149_25071# a_3983_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13978 a_17539_22923# _0964_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X13979 a_3873_7125# a_3707_7125# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13981 a_17727_29967# a_17029_29973# a_17470_29941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13982 vssd1 a_2639_28701# a_2807_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13983 a_25198_28447# a_25030_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13984 vssd1 a_4035_23957# _1773_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X13985 a_9301_5487# a_9135_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13986 vccd1 a_3083_27515# a_2999_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X13987 _1483_.A a_16904_25731# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X13988 vccd1 _0922_.Y a_2953_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X13989 a_16945_12559# _1070_.A2 a_17029_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13990 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7564_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X13991 _1232_.Y a_9963_20175# a_10344_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13992 vccd1 a_1591_5487# fanout28.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13994 _1133_.C a_11858_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X13995 vccd1 _1231_.B1 a_2225_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X13996 vccd1 _1639_.X a_14471_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X13997 a_16615_24349# a_15833_23983# a_16531_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13998 vssd1 a_26451_18811# a_26409_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X13999 vssd1 _1873_.CLK a_24591_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14000 a_10459_27791# a_9761_27797# a_10202_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14001 vccd1 _1192_.A2 a_11934_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X14002 a_21412_20969# _1506_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14003 a_15948_6351# _0993_.X a_15457_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X14004 a_15299_6575# _1065_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14005 a_9384_32143# a_9135_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14006 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_18335_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X14007 a_12650_22351# _1140_.X a_12570_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X14008 a_19877_20719# _1835_.Q a_19439_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14009 vssd1 _1696_.B a_23205_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14010 vccd1 a_19326_29967# a_19432_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X14011 a_10034_27791# a_9595_27797# a_9949_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14012 a_22707_18218# _1500_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14013 vccd1 a_10386_8181# a_10313_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14014 vssd1 _1071_.X a_8178_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X14016 a_3730_22671# _1240_.B1 a_3435_22671# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X14017 vccd1 a_27031_29588# _1353_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14019 _1425_.A a_15939_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14020 a_15568_27247# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X14021 vccd1 _1834_.Q a_19470_22467# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X14022 a_4525_20495# _1327_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X14023 a_4253_10927# _1226_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14024 vssd1 _1090_.C a_17477_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14025 a_10257_27001# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X14026 vccd1 a_27590_26271# a_27517_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14027 vccd1 _1374_.A_N a_23303_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14029 a_7742_6031# _1171_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14030 vssd1 a_22622_24501# a_22580_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14031 vssd1 a_27038_17567# a_26996_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14032 a_19439_24527# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14033 vssd1 a_12299_2589# a_12467_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14035 a_6644_5263# _1208_.A1 a_6559_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14038 a_3249_19453# a_2966_19131# a_2836_19319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14039 a_27238_15645# a_26965_15279# a_27153_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14041 a_12069_23145# _0984_.B1 a_12153_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14042 a_5545_21807# _0913_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X14043 a_20997_6397# a_20727_6031# a_20907_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14045 vccd1 a_15630_29535# a_15557_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14046 vccd1 a_8177_21781# _1294_.B2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X14047 a_5080_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X14048 a_6369_22895# _1328_.S a_6151_22869# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X14049 a_2129_7119# _1791_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14050 a_12604_27497# a_12355_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14051 a_4497_7637# _1168_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X14052 a_5888_28879# a_5639_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14054 a_17470_17973# a_17302_17999# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14055 vssd1 a_23691_3579# a_23649_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14056 a_13360_29199# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X14057 a_17139_5853# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14058 vccd1 _0929_.A a_5269_13367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X14059 a_20635_10205# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14061 vccd1 a_14066_24501# a_13993_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14063 vssd1 _0918_.A a_7667_22901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14065 vccd1 a_25623_6843# a_25539_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14066 a_11868_26409# a_11619_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14067 a_11902_24893# _1287_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X14068 a_8859_6144# _1188_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14069 vccd1 _1985_.CLK a_24591_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14071 _1900_.Q a_15963_25589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14073 a_2073_30287# _1775_.A2 a_1975_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X14075 a_12249_4943# _1751_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14076 vccd1 a_15243_3855# a_15411_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14078 vssd1 a_26394_7775# a_26352_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14079 a_7573_11791# _1164_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14081 vccd1 a_5687_4564# _2001_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14082 a_15917_5461# _1293_.A1 a_16170_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X14083 vccd1 _0913_.A1 a_2408_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14084 _1515_.A a_21412_20969# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X14086 _1900_.Q a_15963_25589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14088 a_15737_15823# _1024_.X a_15483_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14089 vssd1 _1084_.C1 a_1945_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14090 a_19973_32149# a_19807_32149# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14091 _1278_.A1 a_3063_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X14092 a_4422_1679# a_4149_1685# a_4337_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14093 a_16209_16367# _1829_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X14094 vssd1 a_19671_25834# _1876_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14095 a_2198_2335# a_2030_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14096 vccd1 a_14894_30623# a_14821_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14098 a_15565_14013# _1127_.A a_15483_13760# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14099 a_17305_13353# _1403_.B a_17221_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14100 a_26295_2986# _1318_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14101 a_18121_8751# _1719_.B a_18049_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14102 vssd1 a_9779_12015# _1198_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14103 vssd1 _1195_.A2 a_16904_3971# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14104 a_12351_3855# a_12171_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14105 a_12065_8207# _1561_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14106 vssd1 a_8286_27247# a_8392_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14107 vssd1 _1270_.A a_2603_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14108 vccd1 _1590_.A_N a_14103_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
R30 vccd1 temp1.capload\[12\].cap_42.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X14109 vccd1 _0922_.Y a_1757_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X14111 a_23205_19453# a_22935_19087# a_23115_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14112 a_15974_7913# _1040_.X a_15725_7809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X14113 a_12219_24566# _1305_.B a_11760_24759# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X14116 a_2382_7093# a_2214_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14117 vccd1 _1782_.A a_8767_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14118 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14119 a_14674_15529# _1095_.C1 a_14594_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X14120 vssd1 a_23443_9514# _1965_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14121 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_14370_31599# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14122 vssd1 a_23443_31764# _1475_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14123 a_18795_7232# _1061_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14124 vccd1 a_27923_28603# a_27839_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14125 a_22622_1247# a_22454_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14128 vssd1 a_27215_1300# _1951_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14129 a_1643_23413# _1272_.B1 a_1841_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X14130 a_20429_1135# a_19439_1135# a_20303_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14131 a_23443_7338# _1675_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14133 a_12318_8181# a_12150_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14134 vssd1 _1907_.CLK a_11895_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14137 _1293_.A1 a_17139_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14138 a_9363_15101# _1772_.A0 a_9000_14967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X14139 vssd1 _1156_.C _1156_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14140 a_4116_4649# _1801_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14141 a_27295_17821# a_26431_17455# a_27038_17567# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14142 vccd1 _1108_.X a_14537_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X14143 vssd1 a_3210_24501# a_3168_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14144 a_18243_24527# _1424_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14146 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_12631_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X14147 a_7828_6351# _1171_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X14148 vccd1 a_25559_10602# _1720_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14149 a_20131_30186# _1481_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14150 a_15299_17821# _1374_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14151 a_25581_7497# a_24591_7125# a_25455_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14152 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5080_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14153 vccd1 a_13974_21237# a_13901_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14154 vccd1 _1764_.A a_7442_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X14155 vccd1 a_25014_17973# a_24941_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14156 vssd1 _1841_.Q a_16029_29245# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14157 vccd1 a_5455_17455# _1234_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X14158 a_12160_18365# a_11711_17999# a_11858_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14159 a_25589_13647# _1986_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14161 a_25769_6031# a_25235_6037# a_25674_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14163 vccd1 a_23523_2589# a_23691_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14164 vssd1 _1907_.CLK a_11711_8213# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14165 vccd1 a_14123_31029# a_14039_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14166 a_20387_29789# a_19605_29423# a_20303_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14167 a_24547_5162# _1730_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14168 a_22178_5853# a_21739_5487# a_22093_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14169 vccd1 a_23351_32362# _1477_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14170 _1820_.Q a_17895_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14171 vccd1 a_23063_20175# a_23231_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14172 clkbuf_1_1__f_io_in[0].A a_2962_14735# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14173 _1150_.B2 a_23047_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14175 vssd1 _1775_.C1 _1773_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14176 vssd1 a_25842_13621# a_25800_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14177 a_10313_8207# a_9779_8213# a_10218_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14178 vssd1 _0929_.A a_5520_10933# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X14179 vccd1 _1132_.A a_10055_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14181 _1028_.X a_18427_15279# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X14182 a_14986_4917# a_14818_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14183 _1145_.A1 a_8971_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14184 a_2455_1501# a_1591_1135# a_2198_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14185 a_2639_7119# a_1941_7125# a_2382_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14186 a_9292_28879# a_9043_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14187 vccd1 _1474_.A_N a_6743_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14188 vssd1 a_20046_26271# a_20004_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14189 a_12065_13647# _1906_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14190 vccd1 _0992_.A2 a_7659_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14191 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_9384_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14193 vccd1 _1690_.A_N a_27443_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14194 vssd1 a_23063_20175# a_23231_20149# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14195 vccd1 a_22419_31965# a_22587_31867# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14196 vccd1 _1353_.B a_12482_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X14199 vccd1 clkbuf_0_temp1.i_precharge_n.X a_1674_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14200 a_27111_14557# a_26413_14191# a_26854_14303# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14201 vssd1 _1226_.A1 _1246_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14202 vccd1 _0951_.B a_18551_11809# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X14203 a_8803_1679# a_7939_1685# a_8546_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14204 a_15630_29535# a_15462_29789# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14205 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_10699_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X14206 vssd1 _1242_.B1 _1287_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X14209 vssd1 a_12318_13621# a_12276_14025# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14211 _0909_.A _1234_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14212 vccd1 _1140_.C a_11803_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X14213 vccd1 a_27590_19743# a_27517_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14214 vccd1 a_1674_28879# _1329_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14215 a_15289_10927# _1110_.A a_15207_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14216 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_6559_30511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X14217 vssd1 a_21051_4074# _1743_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14218 vssd1 fanout24.A a_23671_10389# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14220 a_24301_14735# _1979_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14221 _1808_.Y a_5165_2828# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X14222 _1148_.B a_10167_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14223 vssd1 a_3467_27791# a_3635_27765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14224 _1074_.C _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14225 a_9773_7663# a_9503_8029# a_9683_8029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14226 vssd1 _1855_.CLK a_13091_31061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14227 a_1757_20969# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14229 a_22572_13967# _1190_.B1 a_22081_13621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X14230 _1637_.X a_16904_3971# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14231 vssd1 a_7711_5652# _1565_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14232 vccd1 fanout12.A a_8307_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X14233 vssd1 a_22898_27765# a_22856_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14234 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12604_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14235 a_25750_29535# a_25582_29789# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14236 _1342_.Y _1342_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14238 vssd1 a_25198_24095# a_25156_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14240 vccd1 _1113_.C a_18519_21376# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X14242 a_21165_4399# a_20175_4399# a_21039_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14243 _1293_.A1 a_17139_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X14245 a_15833_24527# _1474_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14246 vssd1 a_8546_1653# a_8504_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14247 vccd1 _1291_.A1 a_18969_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14248 a_17691_22464# _1870_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14249 a_19878_5853# a_19605_5487# a_19793_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14250 vssd1 a_26007_29789# a_26175_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14251 vccd1 _1119_.A1 a_18607_11293# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14253 vssd1 a_25623_9019# a_25581_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14254 vssd1 _1941_.CLK a_19439_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14255 vssd1 a_27739_9019# a_27697_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14256 vccd1 _1073_.A2 a_17029_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X14257 vssd1 a_20959_26922# _1903_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14258 _1269_.A1 a_6927_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14259 _1007_.A1 a_23691_9019# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14260 a_1841_21807# _1308_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14261 _1438_.B a_13203_10357# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14262 _1762_.A a_7755_21263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14264 a_23105_22351# _1828_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14265 a_4248_26409# _1764_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14266 vccd1 _1261_.A2 a_7111_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X14267 a_9999_5853# a_9135_5487# a_9742_5599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14268 _1375_.A a_8855_22351# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14269 a_12334_15645# a_12061_15279# a_12249_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14270 vssd1 a_26387_9514# _1678_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14271 a_4232_32143# a_3983_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14273 _1048_.X a_18519_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X14274 a_17956_7439# _1744_.B a_17381_7093# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X14275 a_14894_9951# a_14726_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14276 temp1.capload\[11\].cap.Y temp1.capload\[15\].cap.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14277 _1310_.B1 a_7481_23555# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X14278 vccd1 _1904_.Q a_8027_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14279 vccd1 _0989_.A2 a_10094_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X14280 a_26870_6941# a_26431_6575# a_26785_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14282 temp1.capload\[15\].cap.B a_10506_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14283 vccd1 _1108_.A1 a_13948_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X14284 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X14285 _1451_.X a_7567_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14286 _1055_.C a_12027_20495# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X14287 a_5595_22390# _1303_.A1 a_5136_22583# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X14288 vssd1 _1858_.Q a_13316_25321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14289 _1497_.X a_18560_22467# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14290 a_22457_23983# a_22291_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14291 a_17385_19453# _1881_.Q a_17313_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14293 a_20077_13967# _1877_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X14295 a_20487_28701# a_19789_28335# a_20230_28447# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14296 vssd1 a_9195_17973# _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14297 a_17428_28169# a_17029_27797# a_17302_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14298 vccd1 _0909_.X a_25695_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14299 a_13070_2767# a_12797_2773# a_12985_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14301 _1747_.A a_20539_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14302 a_9384_26409# a_9135_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14303 vccd1 a_4351_22359# _1337_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X14304 a_17604_6351# _0997_.X a_17113_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X14305 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_7656_31375# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14306 vccd1 a_16175_1898# _1957_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14307 a_5486_8323# _1782_.A a_5404_8323# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14309 vccd1 _0958_.B a_17691_22464# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X14310 _1403_.B a_24243_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14311 _1756_.X a_6555_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14312 a_24945_2223# _1743_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14313 a_15059_7119# a_14195_7125# a_14802_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14314 _1128_.B a_25991_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14315 _0999_.X a_16863_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X14316 a_20303_26525# a_19439_26159# a_20046_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14317 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14318 a_14287_23261# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14319 a_23063_20175# a_22199_20181# a_22806_20149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14321 a_25750_9951# a_25582_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14322 _1764_.A a_6927_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14323 a_27881_10927# a_26891_10927# a_27755_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14324 vccd1 _1243_.A _1243_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14325 a_25823_8207# a_24959_8213# a_25566_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14326 vccd1 a_1766_26159# _1764_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14327 a_17569_24893# _1873_.Q a_17497_24893# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14328 a_12892_15823# _1071_.B1 a_12637_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X14329 a_17381_14337# _1033_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X14330 vccd1 a_6135_2589# a_6303_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14331 vccd1 a_11759_7338# _1657_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14332 a_14979_17130# _1381_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14333 a_27605_16367# a_26615_16367# a_27479_16733# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14334 vssd1 _1941_.CLK a_15575_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14335 vccd1 a_2382_4511# a_2309_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14336 a_10643_29967# a_9779_29973# a_10386_29941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14338 vssd1 _1308_.B a_2009_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14340 a_25156_31599# a_24757_31599# a_25030_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14342 vccd1 a_9184_23047# _1341_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X14343 a_17861_1135# _1956_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14344 a_6808_32143# a_6559_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14347 vccd1 a_11953_11073# _1050_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14348 a_27973_5487# a_26983_5487# a_27847_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14350 a_20073_13353# _1191_.B1 a_20157_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14352 a_26965_20719# a_26799_20719# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14354 a_2957_27791# _2004_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14355 vccd1 _1999_.CLK a_12631_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14356 vssd1 a_11299_11092# _1439_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14357 vccd1 a_27038_17567# a_26965_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14358 a_27038_13215# a_26870_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14359 _1703_.A a_27623_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14360 a_15285_32143# _1868_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14361 vccd1 _1075_.C a_17967_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X14363 a_21827_22173# a_21647_22173# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14364 _1226_.B1 a_6644_5263# a_7002_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14366 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_9292_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14367 vssd1 _1860_.CLK a_11711_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X14368 vssd1 _2008_.Q _1772_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14369 vccd1 a_10195_13268# _1906_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14370 fanout24.A a_22935_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X14371 vssd1 _1924_.CLK a_24591_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14372 vccd1 _1242_.A1 a_6454_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X14373 _1142_.D1 a_11895_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X14374 a_22603_6941# a_21739_6575# a_22346_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14376 a_2199_21583# _0923_.Y a_1643_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14377 a_22304_5487# a_21905_5487# a_22178_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14378 a_22622_26677# a_22454_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14379 _1763_.A2 a_2686_23439# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14380 vccd1 _1896_.CLK a_19149_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X14381 vssd1 _1448_.A a_8307_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14382 vssd1 _1914_.Q a_20676_12265# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14383 a_13119_10383# a_12337_10389# a_13035_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14384 vccd1 a_19107_2767# a_19275_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14385 vccd1 a_27215_4074# _1367_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14387 a_15235_16733# a_14453_16367# a_15151_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14388 a_15335_2767# a_14471_2773# a_15078_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
D5 vssd1 _1900_.Q sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X14389 vccd1 _1287_.A fanout12.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14390 a_4877_13967# _1217_.A2 a_4627_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14392 a_1674_30511# clkbuf_0_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14393 a_20096_30511# a_19697_30511# a_19970_30877# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14394 vssd1 a_1674_28879# _1329_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14395 a_20249_28885# a_20083_28885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14396 a_22454_26703# a_22181_26709# a_22369_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14397 vssd1 _1436_.B a_11061_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14398 vccd1 a_12575_8207# a_12743_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14399 _1685_.B a_24703_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14400 a_12604_28879# a_12355_28879# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14401 vccd1 a_8215_23983# _1474_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14402 a_19746_18793# _1137_.X a_19497_18689# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X14403 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X14404 temp1.dcdc.A a_5354_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14405 a_2680_22895# a_2649_23047# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X14406 a_25129_16367# _1985_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14407 vssd1 _0921_.A _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14408 a_25539_5853# a_24757_5487# a_25455_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14410 _0913_.Y _0913_.A1 a_5542_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X14411 vssd1 a_13054_25589# a_13012_25993# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14413 _1685_.B a_24703_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14414 a_7277_2223# a_7111_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14415 a_9945_29973# a_9779_29973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14416 a_10257_27001# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X14418 vssd1 a_10667_16885# _1141_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14419 a_15017_28335# a_14747_28701# a_14927_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14420 _1835_.Q a_25623_27515# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14421 a_16185_14337# _1099_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X14422 vssd1 _1982_.CLK a_23246_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14424 a_12488_26409# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14425 a_9889_25913# _1329_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X14426 vssd1 a_15078_2741# a_15036_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14427 _1882_.Q a_27095_25339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14428 a_3789_11791# _1177_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14429 a_21725_30511# _1487_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14430 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_11619_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X14431 a_10147_26409# _0983_.B1 a_10229_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X14433 vssd1 _0929_.A a_5428_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X14434 vccd1 _1639_.X a_6559_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14435 vccd1 a_18940_12533# _0975_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X14436 _1511_.A a_20768_22057# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X14437 vssd1 _2004_.Q a_10791_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14438 _1301_.A1 _1218_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X14439 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4232_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14440 vccd1 a_19487_4564# _1636_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14441 vccd1 _0921_.A _0930_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14442 a_2214_3855# a_1941_3861# a_2129_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14443 vccd1 a_2122_9839# a_2228_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X14444 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_8392_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14445 vssd1 a_16055_29691# a_16013_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14447 a_17302_17999# a_16863_18005# a_17217_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14448 a_5261_10973# _0917_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14450 a_22730_24349# a_22291_23983# a_22645_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14451 a_10218_1679# a_9779_1685# a_10133_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14452 a_10769_6409# a_9779_6037# a_10643_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14454 vssd1 a_2327_20183# _1775_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X14455 vssd1 _1132_.C a_13797_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14456 vssd1 a_9742_4511# a_9700_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14457 vssd1 _1841_.CLK a_19623_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14458 a_10279_16911# _1764_.A a_9921_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14459 a_21617_15279# _1976_.Q a_21545_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14460 a_14641_30511# _1447_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14461 vccd1 a_22063_29098# _1873_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14462 vssd1 _1851_.Q a_9176_19881# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14464 a_20850_22057# _1506_.B a_20768_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14465 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z _1243_.Y a_9384_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14466 vssd1 a_2932_18517# _1302_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X14467 _1376_.X a_11983_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14468 a_26996_6575# a_26597_6575# a_26870_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14469 vccd1 _1013_.X a_9779_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X14470 vssd1 a_15151_16733# a_15319_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14471 vccd1 _2006_.Q a_6835_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14472 _1156_.C a_11711_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X14473 _1144_.X a_9687_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X14474 a_4896_29199# _1342_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X14476 vccd1 _0909_.B a_5911_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X14477 a_27847_3677# a_27149_3311# a_27590_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14478 vccd1 _1023_.B a_19562_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X14479 a_24113_28885# a_23947_28885# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14480 vssd1 a_27463_24251# a_27421_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14481 a_25769_12559# a_25235_12565# a_25674_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14482 a_15013_27791# _1841_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X14483 a_1955_14441# _1223_.B1 a_1737_14165# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X14484 a_10931_2986# _1611_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14485 _1443_.A a_9360_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14486 a_11115_7828# _1614_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14487 a_25581_17455# a_24591_17455# a_25455_17821# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14488 vccd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14489 vccd1 a_4590_1653# a_4517_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14490 _1713_.X a_27347_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14491 vssd1 a_2962_29967# clkbuf_0_temp1.i_precharge_n.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14492 _0922_.Y _0921_.Y a_6651_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14494 a_24945_20719# _1699_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14495 a_4146_7119# a_3873_7125# a_4061_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14496 vssd1 a_16083_17130# _1822_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14497 a_9889_15253# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X14498 a_19651_14735# a_18869_14741# a_19567_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14499 a_7090_1501# a_6651_1135# a_7005_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14501 vccd1 a_6611_29111# _1259_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X14502 _1422_.X a_12488_26409# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X14503 a_23903_19796# _1387_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14504 a_10681_6825# _1562_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X14505 vccd1 a_20046_26271# a_19973_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14506 vccd1 fanout20.X a_22015_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14507 vssd1 a_23266_4917# a_23224_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14510 vccd1 _2009_.CLK _0909_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14511 a_1757_6575# a_1591_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14512 a_26141_7663# _1982_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14514 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14515 _1859_.Q a_17527_31867# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14516 a_23098_2589# a_22825_2223# a_23013_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14517 _1863_.Q a_18355_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14519 a_11497_8751# _1042_.B a_11425_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14520 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14521 a_25087_15823# a_24389_15829# a_24830_15797# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14522 vssd1 a_23351_32362# _1477_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14523 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14524 vssd1 _1010_.A _1071_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14525 a_4351_2589# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14526 a_18114_31029# a_17946_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14527 vccd1 _1261_.A1 a_6553_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X14528 _1141_.C a_10667_16885# a_10279_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14529 a_21491_2589# a_20709_2223# a_21407_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14530 a_11793_6031# _1144_.X a_11711_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14532 a_24619_11471# a_23837_11477# a_24535_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14533 vccd1 a_15795_32143# a_15963_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14536 vccd1 _1850_.CLK a_11711_11477# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14537 a_18940_12533# _1293_.A1 a_19163_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X14538 _1775_.X a_1735_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14539 vccd1 _1590_.A_N a_11527_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14541 vssd1 a_4519_9991# _1172_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X14542 a_7531_9813# _1158_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X14543 vccd1 a_23535_23060# _1972_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14544 a_18371_1501# a_17507_1135# a_18114_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14545 a_25953_7663# a_25787_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14546 a_3514_25615# _1761_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14547 vccd1 _1685_.B a_23759_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14548 a_14910_2767# a_14471_2773# a_14825_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14549 vssd1 _1982_.CLK a_22015_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X14550 vssd1 a_15795_32143# a_15963_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14551 a_21647_22173# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14552 a_26965_20719# a_26799_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14553 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_11960_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14554 _1270_.A a_10423_23983# a_10951_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14555 a_4433_17999# _0925_.A2 a_4351_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14557 vccd1 _1111_.B a_21459_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14560 a_10402_19997# a_10129_19631# a_10317_19631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14561 vccd1 _2023_.CLK a_3707_7125# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14563 a_25014_2741# a_24846_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14564 vccd1 a_12575_11471# a_12743_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14566 a_4341_6621# _1210_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14569 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A a_8944_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14571 vssd1 a_27479_16733# a_27647_16635# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14573 a_15285_31055# _1465_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14574 vssd1 a_22346_5599# a_22304_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14575 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.A a_14370_31599# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14576 a_27675_29588# _1463_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14577 vccd1 _1826_.Q a_18642_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X14579 a_15207_10927# _1088_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14580 vssd1 a_12575_11471# a_12743_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14581 a_18427_28701# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14583 _1088_.B a_19275_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14585 vccd1 a_12189_18150# a_11858_17973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X14586 a_6739_2767# a_6559_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14587 vccd1 a_2623_1403# a_2539_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14588 vssd1 _1145_.B2 a_11797_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14589 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_12604_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14590 a_26686_14557# a_26247_14191# a_26601_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14591 _1098_.B a_23691_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14592 a_4163_4943# _1802_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14593 a_18699_26703# a_18519_26703# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14594 vssd1 a_8654_29967# a_8760_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14595 vssd1 _1887_.CLK a_22751_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X14596 a_11527_17821# _2004_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14597 _1231_.B1 a_5455_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X14598 vssd1 _1150_.B2 a_20353_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14599 a_1673_22453# _2009_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14600 vccd1 a_8971_1653# a_8887_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14601 vccd1 _1086_.Y a_3605_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14602 vccd1 a_25743_1898# _1952_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14603 vssd1 a_27859_30676# _1450_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14604 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5908_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14605 vccd1 a_8548_23413# _1329_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14606 vccd1 _0922_.Y a_1965_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14607 a_15882_19087# _1020_.D1 a_15633_19061# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X14608 a_22369_31055# _1874_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14609 a_27590_5599# a_27422_5853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14610 vccd1 a_9871_10391# _1537_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X14612 vccd1 a_5731_12567# _1325_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X14613 a_19954_31029# a_19786_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14614 vccd1 a_6703_26133# _1306_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X14615 vssd1 _1075_.C a_17845_21629# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14616 a_20062_28701# a_19789_28335# a_19977_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14617 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14619 vccd1 _2004_.Q a_6927_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14620 vssd1 a_21407_2589# a_21575_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14621 vccd1 a_15151_30877# a_15319_30779# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14623 vssd1 a_19497_18689# _1138_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X14624 a_22063_9514# _1577_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14625 a_6900_31055# a_6651_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14626 vssd1 a_2686_23439# _1763_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14627 vssd1 a_16863_9295# _0939_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14628 _1528_.A a_26267_16885# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14629 vssd1 _1451_.B a_7657_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14630 vssd1 _1985_.CLK a_24591_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14631 _1149_.C1 a_11711_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X14632 _1062_.X a_17967_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X14633 vssd1 a_3514_25615# clkbuf_1_1__f__0380_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14634 vccd1 a_13019_20495# _1781_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X14635 a_9205_3145# a_8215_2773# a_9079_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14636 a_13545_31599# a_13275_31965# a_13455_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14637 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14639 a_5911_16617# _1325_.A2 a_5693_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X14640 _0909_.X a_3801_28981# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X14643 vccd1 _1823_.CLK a_25235_16917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14644 a_12318_1247# a_12150_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14646 clkbuf_0_temp1.i_precharge_n.X a_2962_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14647 a_3299_22325# _1329_.S a_3517_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X14648 vssd1 _1979_.Q a_27437_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14649 _1697_.A a_23115_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14650 _1862_.Q a_18539_31029# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
D6 vssd1 _1337_.A0 sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X14651 a_22563_13469# a_22383_13469# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14652 vccd1 _1424_.A_N a_15759_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14653 vccd1 a_17565_24129# _1134_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14654 a_2490_27613# a_2217_27247# a_2405_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14655 vssd1 _0956_.C a_10699_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14656 vssd1 a_17113_6005# _0999_.C1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X14657 a_13101_20495# _1781_.B a_13019_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X14658 vssd1 _0981_.B a_16245_9867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X14660 a_10344_2057# a_9945_1685# a_10218_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14661 vccd1 a_25623_27515# a_25539_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14662 _1862_.Q a_18539_31029# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14663 _1132_.A a_10883_21271# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X14664 vccd1 a_26099_16911# a_26267_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14665 vssd1 a_17727_1679# a_17895_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14666 a_16117_10927# _1127_.A a_16035_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14667 a_17029_18005# a_16863_18005# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14668 a_25539_17821# a_24757_17455# a_25455_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14669 _1667_.X a_18239_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14670 a_19325_20495# _1836_.Q a_18887_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14672 vccd1 _1766_.A0 a_8387_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14673 a_13948_14735# _1105_.X a_13846_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X14674 vssd1 _1887_.CLK a_26063_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14675 a_12325_8751# _1043_.B a_12253_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14676 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_15943_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14677 vssd1 _1985_.CLK a_24223_15829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14678 a_10073_23737# _1328_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X14679 _1699_.A a_23023_21085# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X14680 vssd1 _0961_.A _0987_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14681 a_10386_6005# a_10218_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14682 vccd1 a_8307_31599# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X14683 a_14833_30333# a_14563_29967# a_14743_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14684 a_12885_5321# a_11895_4949# a_12759_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14685 vssd1 a_27847_10205# a_28015_10107# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14686 a_2999_24349# a_2217_23983# a_2915_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14688 a_8293_1679# _1565_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14689 a_8914_23439# _0918_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14692 _1043_.B a_16607_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14693 _0930_.B _0929_.A a_10515_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14694 a_28083_16911# a_27903_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14696 a_27847_12381# a_27149_12015# a_27590_12127# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14699 a_27253_27023# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14700 vssd1 a_17895_27765# a_17853_28169# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14701 a_23098_22173# a_22825_21807# a_23013_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14702 vssd1 a_7442_17429# _1140_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14705 vssd1 a_20471_1403# a_20429_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14706 a_11793_7663# _1153_.A a_11711_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14707 a_12575_11471# a_11711_11477# a_12318_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14708 a_2225_17705# _1250_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X14709 vccd1 a_3983_17455# _0921_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14711 vccd1 a_15227_7093# a_15143_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14712 _1577_.B a_12539_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X14713 a_4547_24305# _1772_.A0 a_4035_23957# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X14714 a_15081_22325# _1116_.D1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X14715 vccd1 _2007_.Q _1053_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14716 vccd1 _1021_.A a_13367_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14717 vccd1 _1448_.A a_7571_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X14718 a_9503_1501# _1590_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14720 vssd1 _0984_.B1 a_13448_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X14721 vssd1 a_9920_25223# _1349_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X14722 _1813_.Q a_10811_8181# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14723 vccd1 _1903_.Q a_7935_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14724 a_27399_16042# _1700_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14725 a_7216_1135# a_6817_1135# a_7090_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14726 a_5169_13149# _0916_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14727 vccd1 a_25991_8181# a_25907_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14728 vccd1 _1330_.X a_21371_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14729 vssd1 a_26670_23007# a_26628_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14730 vssd1 a_7803_20884# _1852_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14731 a_5060_32143# a_4811_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14732 vccd1 _1374_.A_N a_15207_14557# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14733 vssd1 a_16185_14337# _1104_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X14734 a_22383_8029# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14735 a_2121_12015# _1208_.A1 a_1775_12265# vssd1 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X14736 a_15637_14013# _1019_.B a_15565_14013# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X14739 vssd1 a_1766_26159# _1764_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14740 vssd1 a_8447_7828# _1751_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14741 vssd1 a_3635_27765# _2004_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14742 a_12245_11471# a_11711_11477# a_12150_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14743 a_15277_26159# _1476_.B a_14839_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14744 a_15299_20291# _1181_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X14745 vccd1 a_27847_19997# a_28015_19899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14746 a_17573_4917# _0952_.A1 a_17826_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X14748 a_7657_31599# a_7387_31965# a_7567_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14751 _0951_.B a_10814_14709# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14752 a_11858_17973# _2004_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X14753 a_24945_31599# _1873_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14754 vccd1 a_25255_15797# a_25171_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14757 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14758 vssd1 _1816_.CLK a_7939_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14759 _1007_.A1 a_23691_9019# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14760 _1597_.A a_19619_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14761 vccd1 a_26007_10205# a_26175_10107# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14762 vssd1 a_25455_17821# a_25623_17723# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14764 a_15243_4943# a_14379_4949# a_14986_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14765 vssd1 _0925_.A2 a_2695_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X14766 a_25455_7119# a_24591_7125# a_25198_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14767 a_23565_16911# _1831_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14768 a_27153_20719# _1823_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14769 vccd1 _1153_.A a_16863_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14770 vccd1 _1007_.A1 a_20815_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14771 a_8120_27791# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14772 _1769_.Y _1775_.C1 a_3993_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14773 vccd1 a_11760_23671# _1346_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X14774 a_4035_30485# _1353_.A a_4244_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X14775 a_22695_29789# a_21831_29423# a_22438_29535# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14776 a_4932_16911# _1249_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14777 a_10585_2223# a_9595_2223# a_10459_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14778 vssd1 _0923_.Y a_6968_21379# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14779 a_11601_2223# a_11435_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14780 a_27973_27247# a_26983_27247# a_27847_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14781 vssd1 _1855_.CLK a_12447_25621# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14783 a_3007_1679# a_2143_1685# a_2750_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14784 a_22101_30287# temp1.capload\[15\].cap.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14785 vccd1 clkbuf_0_temp1.dcdel_capnode_notouch_.X a_15750_28335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14786 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14787 _1782_.A a_4627_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X14788 _1110_.X a_18519_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X14791 _1112_.A1 a_26819_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14793 vccd1 a_1735_29941# _1775_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X14795 vccd1 a_22771_6843# a_22687_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14796 a_18455_31055# a_17673_31061# a_18371_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14797 a_11969_25437# a_11435_25071# a_11874_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14798 a_3965_16911# _1291_.B2 a_3881_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14799 a_17139_17024# _1822_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X14800 a_20648_28169# a_20249_27797# a_20522_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14801 a_12232_18365# a_12189_18150# a_12160_18365# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X14802 a_10147_3855# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14803 _1246_.B2 _1221_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14804 vssd1 a_6847_22057# _1328_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14805 a_19985_17231# _1914_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X14806 vccd1 _1226_.A1 _1217_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14807 vccd1 a_27831_22075# a_27747_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14809 a_22365_29789# a_21831_29423# a_22270_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14810 a_27011_23261# a_26229_22895# a_26927_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14811 a_26099_22351# a_25401_22357# a_25842_22325# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14812 a_26099_16911# a_25235_16917# a_25842_16885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14813 _1219_.B1 a_7201_14851# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X14816 vccd1 a_15503_2741# a_15419_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X14817 vccd1 a_13403_12559# a_13571_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14818 a_17352_14735# _1091_.B1 a_17250_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X14819 vssd1 a_26099_6031# a_26267_6005# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14820 a_13698_31029# a_13530_31055# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14821 vssd1 a_26267_6005# a_26225_6409# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14822 a_19521_20969# _1184_.B1 a_19605_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14823 a_27111_14557# a_26247_14191# a_26854_14303# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14824 a_23299_14557# a_23119_14557# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14825 vssd1 a_21207_4667# a_21165_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14826 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A a_6900_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14828 a_14144_26819# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14830 a_19973_5853# a_19439_5487# a_19878_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14831 vssd1 a_19326_29967# a_19432_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14832 vssd1 a_2750_1653# a_2708_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14833 a_15163_4564# _1621_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X14834 a_27149_5487# a_26983_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14835 vssd1 a_13403_12559# a_13571_12533# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14836 vssd1 _1282_.A2 a_6469_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X14837 a_5664_24233# _1287_.A a_5203_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X14838 _1824_.Q a_27647_16635# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14840 a_14379_18793# _1073_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X14842 vccd1 a_8723_4074# _1567_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14843 vssd1 a_11023_31274# _1868_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14844 vssd1 a_27406_20831# a_27364_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14845 a_2195_12533# _1301_.A1 a_2626_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X14846 a_13530_31055# a_13257_31061# a_13445_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14847 _1126_.Y _1125_.X a_6743_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X14849 a_5167_19407# _1301_.A1 _1327_.A1_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X14850 a_6743_10383# _1324_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14851 a_27437_12925# a_27167_12559# a_27347_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X14852 a_2122_8029# a_1849_7663# a_2037_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14854 a_19619_24527# a_19439_24527# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14855 vssd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14857 vccd1 a_10287_2986# _1659_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14858 vccd1 a_25271_2767# a_25439_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14859 vssd1 a_10471_7828# _1813_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14860 vssd1 a_2455_8207# a_2623_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14861 a_25984_18543# a_25585_18543# a_25858_18909# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14862 vssd1 _1113_.C a_17257_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X14863 vssd1 a_26479_1300# _1616_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14864 a_2723_4943# a_1941_4949# a_2639_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14865 a_20591_7338# _1747_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X14867 a_15753_19881# _0975_.X a_15657_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X14868 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_5080_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14869 vssd1 _1006_.B2 a_22572_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X14870 vccd1 a_24087_6250# _1674_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14871 vccd1 _1019_.B a_17319_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X14872 a_22825_10927# a_22659_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14873 a_9945_1685# a_9779_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X14874 vccd1 a_2382_3829# a_2309_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14875 a_16945_8573# _1153_.A a_16863_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14876 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14877 vssd1 _0994_.A2 a_15432_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X14878 _1458_.A a_10740_25731# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14879 vssd1 a_24639_14356# _1984_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X14880 a_15614_6031# _0994_.B2 a_15457_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
R31 vssd1 temp1.capload\[15\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X14881 a_26965_24349# a_26431_23983# a_26870_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X14882 vccd1 _1839_.Q a_12478_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X14883 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13360_29199# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X14884 vccd1 a_5871_23658# _1819_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14885 a_15538_31029# a_15370_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14886 a_15243_3855# a_14545_3861# a_14986_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14887 a_27038_6687# a_26870_6941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14888 vssd1 _1347_.Y a_8215_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X14889 a_22898_24095# a_22730_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14890 a_8295_15279# _1261_.A1 _1790_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X14891 vssd1 _1977_.Q a_22653_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X14892 a_13488_9001# _0987_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X14893 a_10862_27613# a_10423_27247# a_10777_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14896 a_23098_3677# a_22659_3311# a_23013_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14901 _1170_.B1 a_5496_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14902 _1903_.Q a_10627_29691# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14903 a_12150_29789# a_11711_29423# a_12065_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14904 a_25030_13469# a_24757_13103# a_24945_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14905 a_22563_12381# a_22383_12381# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X14906 vccd1 _0935_.X a_9595_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14908 vssd1 _1242_.A2 a_8204_28111# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X14909 vssd1 _0922_.Y a_3041_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X14910 vccd1 a_19497_18689# _1138_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X14911 a_1775_26703# _1773_.B _1773_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14912 a_18064_5263# _0997_.X a_17573_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X14913 vssd1 a_2715_13371# a_2673_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14915 vccd1 a_2455_2589# a_2623_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14917 a_7656_11471# _1156_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14918 _1431_.A a_13040_23555# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X14920 a_13714_1679# a_13441_1685# a_13629_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X14923 a_26367_18909# a_25585_18543# a_26283_18909# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14924 a_9167_14219# _1286_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X14925 vccd1 _1321_.C a_5632_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X14926 _1982_.CLK a_22050_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X14929 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_5060_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X14930 vccd1 a_5565_22649# a_5595_22390# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X14931 a_17470_17973# a_17302_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14932 vccd1 _1127_.A a_17691_8320# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14933 a_8286_27247# a_8109_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X14934 vccd1 _1277_.B a_2505_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X14935 vssd1 _1032_.C a_17385_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X14936 a_19899_13647# _1191_.B1 a_20077_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X14937 a_2539_8207# a_1757_8213# a_2455_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14940 a_9489_4399# _1753_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X14941 a_20372_32521# a_19973_32149# a_20246_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14942 a_5829_15529# _0930_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14943 vccd1 a_12318_11445# a_12245_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14944 vccd1 _1273_.A1 a_6559_15936# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14945 a_14818_4943# a_14379_4949# a_14733_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14946 vccd1 a_4314_7093# a_4241_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14947 _1759_.A a_8947_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14948 vssd1 a_7258_1247# a_7216_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X14949 a_5449_6351# _1207_.B1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14951 vccd1 _1489_.A_N a_20911_24349# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X14952 a_27406_21919# a_27238_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X14954 vccd1 a_23523_22173# a_23691_22075# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X14955 _1362_.X a_10603_9117# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X14956 vccd1 _1896_.CLK a_19807_32149# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14957 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14958 vssd1 _1308_.B a_1937_22711# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X14959 a_23607_3677# a_22825_3311# a_23523_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14960 clkbuf_0_net57.X a_2594_31055# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14961 a_15512_22351# _1116_.B1 a_15410_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X14963 a_15750_28335# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14964 vccd1 a_23266_2335# a_23193_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14965 a_8955_11791# _1121_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14966 _1240_.B1 a_2603_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X14967 a_13403_12559# a_12539_12565# a_13146_12533# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14968 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X14969 a_8101_2223# a_7111_2223# a_7975_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X14972 vccd1 _1887_.CLK a_22659_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X14974 a_9844_27497# a_9595_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X14975 a_7561_22941# _0921_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X14976 a_20947_11471# a_20083_11477# a_20690_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X14977 vssd1 _1202_.Y a_6644_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14979 a_4422_25437# a_3983_25071# a_4337_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X14982 a_13955_31055# a_13257_31061# a_13698_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X14983 _2006_.Q a_3635_24501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14984 a_22963_24527# a_22181_24533# a_22879_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X14985 a_5241_13647# _1249_.A2 _1230_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14986 a_15929_3311# _1610_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X14987 vssd1 _1999_.CLK a_14471_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X14988 vccd1 a_18475_30676# _1842_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X14989 _1798_.Y a_5625_5792# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
X14990 a_19889_10749# _1153_.A a_19807_10496# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X14991 a_4035_23957# _1772_.A0 a_4244_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X14993 vccd1 _1321_.C a_5547_12015# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X14996 a_25156_15279# a_24757_15279# a_25030_15645# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X14999 vccd1 a_27215_17130# _1389_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15000 a_13073_12559# a_12539_12565# a_12978_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15001 vccd1 _0935_.X a_15115_9408# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15002 a_11023_26922# _1458_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15003 a_22653_13103# a_22383_13469# a_22563_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15004 _1389_.A a_23483_15823# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15005 _1041_.C1 a_12907_7232# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15006 vccd1 a_22438_29535# a_22365_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15007 a_24075_23439# a_23377_23445# a_23818_23413# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15008 a_13524_26409# a_13275_26159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X15009 a_4709_9295# _1226_.B1 _1246_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X15010 vccd1 a_26007_3677# a_26175_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15011 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_1932_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15012 _1306_.A2 _1305_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15015 vccd1 a_6835_18543# _1768_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15016 a_17773_8573# _1127_.A a_17691_8320# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15017 vssd1 a_23535_23060# _1972_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15018 a_22622_2741# a_22454_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15019 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_6559_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15020 a_19793_29423# _1471_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15021 a_5416_21781# _1775_.A2 a_5639_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X15022 vccd1 clkbuf_0_temp1.i_precharge_n.X a_1674_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15023 a_3237_17705# _1311_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X15024 fanout21.X a_23246_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15025 vccd1 _1780_.B1 a_5625_5792# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X15026 vccd1 temp1.capload\[12\].cap.A temp1.capload\[12\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15027 a_1941_6037# a_1775_6037# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15029 vccd1 a_27739_9019# a_27655_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15031 a_20245_17231# _1968_.Q a_19807_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X15032 _1601_.A a_20308_9001# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15033 a_13162_29967# a_12723_29973# a_13077_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15034 vssd1 a_7479_28887# temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X15035 a_25401_22357# a_25235_22357# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15036 vccd1 _1780_.B1 a_8109_14796# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X15038 _1138_.B1 a_19439_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15041 vssd1 a_12226_16341# _0963_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15042 vccd1 _1690_.A_N a_22751_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15043 a_14927_28701# a_14747_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15044 a_22093_5487# _1923_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
R32 temp1.capload\[4\].cap_49.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X15045 vccd1 _1403_.B a_19619_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15046 vssd1 _1021_.A a_13551_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X15047 a_2581_6575# a_1591_6575# a_2455_6941# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15048 _1127_.A a_14839_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X15049 vssd1 _1234_.A1 _0909_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15050 vccd1 temp1.capload\[2\].cap_47.LO temp1.capload\[2\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15051 vssd1 a_12771_3476# _1624_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15053 a_16035_10927# _1037_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X15054 temp1.capload\[8\].cap.Y temp1.capload\[8\].cap_53.LO a_25413_30287# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15055 vssd1 _1841_.CLK a_16863_29973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15056 a_15833_23983# a_15667_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15057 _1024_.D1 a_17415_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15058 a_10202_2335# a_10034_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15059 vssd1 a_23742_4399# a_23848_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15060 vssd1 a_25750_26271# a_25708_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15061 vccd1 _0983_.A2 a_10229_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X15062 a_17904_15823# _1029_.B1 a_17802_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X15063 a_20522_11471# a_20249_11477# a_20437_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15064 a_22645_18543# _1393_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15066 vssd1 _0965_.A2 a_15840_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X15067 a_14265_2057# a_13275_1685# a_14139_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15068 a_7189_13408# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15069 a_5417_18517# _1234_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X15070 a_14737_18115# _1142_.X a_14655_18115# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X15071 a_11793_15101# _0964_.A a_11711_14848# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15072 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_5448_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X15073 _1269_.A1 a_6927_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X15074 vccd1 _1090_.C a_12171_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X15075 vccd1 _1424_.A_N a_18059_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15077 vccd1 a_9613_16600# a_9282_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X15078 _1045_.B1 a_11343_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
R33 vssd1 temp1.capload\[1\].cap.A sky130_fd_pr__res_generic_po w=0.48 l=0.045
X15079 a_21997_29423# a_21831_29423# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15080 a_3551_24527# a_2769_24533# a_3467_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15081 a_19107_3855# a_18243_3861# a_18850_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15083 a_4248_26409# _1273_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15084 a_15667_24527# _0966_.B1 a_15845_24847# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X15085 a_20709_22895# a_20543_22895# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15086 a_23224_3311# a_22825_3311# a_23098_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15087 _1112_.A1 a_26819_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15088 a_22825_10927# a_22659_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15089 _1308_.B _0921_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X15090 a_17894_24233# _1132_.X a_17814_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X15091 a_7288_15095# a_7101_14735# a_7201_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X15092 a_21327_1300# _1734_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15094 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15095 _1674_.A a_20907_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X15096 a_17923_26922# _1461_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15098 a_3185_20495# _1257_.B2 a_3276_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15099 a_14092_15055# _1108_.A1 a_13517_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X15100 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_4968_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15101 vccd1 a_20039_5162# _1929_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15102 a_4241_7119# a_3707_7125# a_4146_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15104 vccd1 _1941_.CLK a_17507_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15105 vssd1 _1830_.CLK a_20083_11477# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15106 vssd1 a_1643_21781# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15108 a_17302_29967# a_17029_29973# a_17217_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15109 vssd1 fanout20.X a_21739_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15110 vssd1 a_14839_11471# _1127_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15112 vssd1 a_20407_2986# _1989_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15114 a_22622_2741# a_22454_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15115 a_17409_5487# a_17139_5853# a_17319_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15116 vssd1 a_14491_24501# a_14449_24905# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15118 a_11023_16042# _1371_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15120 vssd1 _1032_.C a_21617_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15121 a_17270_6031# _1047_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X15122 a_21077_2589# a_20543_2223# a_20982_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15123 a_26651_4765# a_25953_4399# a_26394_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15124 a_23193_2589# a_22659_2223# a_23098_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15126 vccd1 a_6245_14165# _1810_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15127 a_17485_31599# a_16495_31599# a_17359_31965# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15129 a_13311_25615# a_12613_25621# a_13054_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15130 a_2472_19605# _1310_.B1 a_2864_19881# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X15131 a_20267_15279# _1046_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X15132 a_19605_29423# a_19439_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15133 vccd1 _1267_.A1 a_4198_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X15134 a_15879_31055# a_15097_31061# a_15795_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15135 a_22235_30877# a_21537_30511# a_21978_30623# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15136 a_26417_25071# _1882_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15138 vccd1 clkbuf_1_1__f__0380_.A a_1766_26159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15139 vssd1 _1764_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X15141 a_13316_25321# _1484_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15142 _0958_.B a_14563_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X15143 vccd1 a_2686_15823# _2009_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15144 vccd1 a_9429_15033# a_9459_14774# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15145 a_14944_5321# a_14545_4949# a_14818_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15146 a_2330_31921# a_2281_31751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X15147 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_9844_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15148 vccd1 _0989_.B2 a_9683_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15149 a_22369_1679# _1940_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15151 _1242_.A2 a_7111_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15152 a_1769_23145# _0925_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X15153 vssd1 a_4127_22869# _1285_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X15154 vccd1 a_12973_5461# _1196_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X15155 a_26785_6575# _1676_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15156 vccd1 _0983_.B1 a_12637_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15158 a_8447_6740# _1359_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15160 _1337_.S a_4351_22359# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X15161 _1924_.CLK a_22015_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X15162 vccd1 _1880_.CLK a_16863_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X15163 a_25198_20831# a_25030_21085# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15164 a_18777_2767# a_18243_2773# a_18682_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15165 a_12575_1501# a_11711_1135# a_12318_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15166 a_10769_30345# a_9779_29973# a_10643_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15169 vccd1 _1170_.A2 _1202_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15170 a_23013_8751# _1920_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15171 _1130_.C1 a_18243_12015# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15172 a_7821_23145# _0921_.B a_7749_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X15173 a_17217_17999# _1820_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15174 vccd1 a_18611_15823# _1506_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15175 a_25271_2767# a_24407_2773# a_25014_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15176 a_22687_5853# a_21905_5487# a_22603_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15177 vssd1 _1173_.X a_7828_6351# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X15178 vccd1 a_6927_17999# _1764_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15179 vccd1 a_8785_15974# a_8454_15797# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X15180 a_19480_11177# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15181 vssd1 a_23523_3677# a_23691_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15182 vccd1 a_13146_12533# a_13073_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15183 a_10865_31599# a_10699_31599# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15187 vssd1 a_26267_26677# a_26225_27081# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15188 vssd1 a_17470_17973# a_17428_18377# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15189 a_27379_13469# a_26597_13103# a_27295_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15190 a_21407_8029# a_20709_7663# a_21150_7775# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15192 a_22457_18543# a_22291_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15193 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_13524_26409# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15195 _1851_.Q a_14399_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15196 vccd1 a_15411_4917# a_15327_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15197 a_19651_1679# a_18869_1685# a_19567_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15198 vccd1 a_25623_7093# a_25539_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15199 a_26007_26525# a_25143_26159# a_25750_26271# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15200 vssd1 _1832_.Q a_18836_23555# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15201 vssd1 a_20303_29789# a_20471_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15202 _1100_.X a_14747_19631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15203 _0984_.X a_12171_23983# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X15204 vccd1 _0930_.Y a_2966_19131# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X15205 _1049_.B1 a_20267_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15207 _1851_.Q a_14399_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15208 a_20157_13353# _1878_.Q a_20073_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15209 a_24646_19061# a_24478_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15211 a_17749_9269# _1112_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X15213 vccd1 a_25559_21482# _1699_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15215 a_19107_2767# a_18409_2773# a_18850_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15217 vccd1 a_25842_13621# a_25769_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15218 vssd1 a_25014_2741# a_24972_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15222 vssd1 _1896_.CLK a_19149_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15224 _1249_.A2 a_2472_15431# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X15226 a_2585_29423# _1775_.A2 a_2485_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X15227 _1461_.A a_13316_25321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X15228 a_25589_24527# _1513_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15229 a_3979_9295# _1177_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15230 a_25677_26525# a_25143_26159# a_25582_26525# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15231 vssd1 a_7366_15279# a_7472_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15232 a_13599_1300# _1645_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15233 a_13183_11177# _1197_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X15234 vssd1 a_24823_28010# _1902_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15235 vccd1 _1789_.A1 a_6923_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X15238 _1237_.B2 _1234_.Y a_4903_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15239 a_24478_19087# a_24205_19093# a_24393_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15240 _1904_.Q a_11455_27515# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15243 a_19977_28335# _1429_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15244 a_10073_23737# _1328_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X15245 a_10951_22057# a_10423_21807# _0925_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15247 a_1643_21237# _0923_.Y a_2199_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15248 _1045_.C1 a_12171_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15249 vssd1 a_16175_9514# input3.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15250 vccd1 a_19567_14735# a_19735_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15251 vssd1 a_24087_6250# _1674_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15252 vccd1 _1084_.C1 a_1945_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X15254 vccd1 a_17831_11092# _1584_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15255 a_1674_30511# clkbuf_0_net57.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15256 _1902_.Q a_12743_29691# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15258 vssd1 io_in[4] a_1626_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15259 a_20676_12265# _1577_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15260 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_12482_27791# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15261 vccd1 _0984_.A2 a_11793_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X15262 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE _1306_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15263 _1586_.A a_19480_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X15264 a_12889_29973# a_12723_29973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15265 a_2129_28335# _1775_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15267 a_17102_26271# a_16934_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15268 a_18682_3855# a_18243_3861# a_18597_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15269 a_13455_31965# a_13275_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15270 vccd1 _1267_.A1 a_5889_10089# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X15271 a_2706_21583# _1260_.B1 a_1643_21237# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.08775 ps=0.92 w=0.65 l=0.15
X15272 fanout12.A _1287_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15274 vssd1 _1882_.CLK a_23671_21269# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15276 _1086_.Y _1086_.B a_7019_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15277 a_18560_23145# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15278 _1064_.D1 a_14471_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15279 vccd1 _0974_.A2 a_19069_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X15280 vccd1 a_2290_7775# a_2217_8029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15282 vssd1 _0985_.X _1012_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15283 a_24757_5487# a_24591_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15284 vccd1 _1084_.B1 a_7993_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X15285 _1580_.A a_19388_8323# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15286 vssd1 a_27031_29588# _1353_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15287 vccd1 a_2971_16367# _0921_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15290 _1316_.A a_9167_14219# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X15292 a_6559_26703# _1242_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15293 a_2497_1679# _1651_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15294 vssd1 a_5136_22583# _1303_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X15295 a_23837_10389# a_23671_10389# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15296 vccd1 a_7387_15823# _1775_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15297 vssd1 a_25623_31867# a_25581_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15298 a_13599_29588# _1469_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15299 a_19395_5162# _1667_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15300 a_24639_7828# _1717_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15301 a_13257_31061# a_13091_31061# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15304 a_13183_21807# _1857_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X15306 vssd1 a_23266_3423# a_23224_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15307 vssd1 a_9742_31029# a_9700_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15308 a_20601_15797# _1081_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X15309 _1156_.D a_16863_11177# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X15310 a_20261_23983# a_19991_24349# a_20171_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15312 a_10730_12675# _0987_.B a_10648_12675# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15313 a_11030_27359# a_10862_27613# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15314 vccd1 _1242_.A2 a_2009_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15316 vccd1 _0964_.A a_16219_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15317 a_3217_8751# _1170_.A2 a_3145_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15318 a_4601_12879# _1217_.A2 a_4351_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15319 a_4805_4175# a_4613_3916# _2019_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X15321 vssd1 a_20223_8426# _1582_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15322 vssd1 _0913_.A1 a_13101_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X15323 vssd1 a_13551_17999# _0958_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X15326 vssd1 _1053_.A a_15299_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X15327 a_16189_10927# _1037_.B a_16117_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15328 vssd1 _0935_.X a_16863_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X15329 clkbuf_1_1__f__0380_.A a_3514_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X15330 a_14315_21263# a_13533_21269# a_14231_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15331 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15332 a_19826_18793# _1138_.C1 a_19746_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X15333 a_11858_17973# a_11711_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X15335 a_15588_29423# a_15189_29423# a_15462_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15337 vssd1 _1033_.A2 a_17956_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X15338 vssd1 _2009_.CLK a_2051_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15339 vccd1 a_13882_1653# a_13809_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15341 _1018_.X a_14379_20719# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15342 vssd1 a_16921_14709# _1091_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X15343 a_24846_2767# a_24407_2773# a_24761_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15344 vssd1 clkbuf_0_temp1.i_precharge_n.A a_2962_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15345 vccd1 _0994_.A2 a_15614_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X15346 a_9176_19881# _1422_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15348 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A a_5908_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X15349 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15350 vssd1 a_1779_22453# _1272_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15351 a_22285_4399# a_22015_4765# a_22195_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15352 a_24462_25589# a_24294_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15353 a_14920_23983# _1862_.Q a_14345_24129# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X15356 a_2198_6687# a_2030_6941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15358 _1504_.A a_21827_22173# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15360 a_20614_4765# a_20341_4399# a_20529_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15361 vccd1 _1084_.C1 _1052_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X15362 vssd1 _1572_.B a_14557_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15363 a_24547_5162# _1730_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15364 vccd1 _1165_.C _1210_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15365 a_10601_9661# a_10331_9295# a_10511_9295# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15366 vssd1 _1347_.Y a_9043_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15367 vssd1 _1132_.C a_14993_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15368 a_27053_25071# a_26063_25071# a_26927_25437# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15369 vccd1 _1140_.C a_13183_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X15370 a_24478_19087# a_24039_19093# a_24393_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15372 a_9779_11471# _1104_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15373 a_7567_31965# a_7387_31965# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15375 vccd1 a_25807_16635# a_25723_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15376 vssd1 clkbuf_1_1__f_io_in[0].A a_2686_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15377 vssd1 _1868_.Q a_14604_27497# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15378 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15380 a_26996_23983# a_26597_23983# a_26870_24349# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15381 vssd1 _1250_.A1 a_1929_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15382 vssd1 a_10627_2491# a_10585_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15383 vssd1 a_27571_9117# a_27739_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15384 vssd1 a_25455_9117# a_25623_9019# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15385 vssd1 a_23266_11039# a_23224_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15387 a_8392_14735# _1793_.A2 _1793_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X15388 vssd1 _1941_.CLK a_15759_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15389 a_11053_31599# _1855_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15390 vssd1 a_20563_30779# a_20521_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15391 vccd1 _1880_.CLK a_22567_25071# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X15392 vssd1 a_2658_24095# a_2616_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15393 vssd1 a_2472_15431# _1249_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X15394 a_23299_13647# a_23119_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15395 a_14287_13353# _1120_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X15396 a_20429_5487# a_19439_5487# a_20303_5853# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15397 a_19567_14735# a_18703_14741# a_19310_14709# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15398 a_9761_29423# a_9595_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15399 a_27859_30186# _1456_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15400 a_27295_6941# a_26431_6575# a_27038_6687# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15402 _0909_.C _2009_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15403 a_7101_14735# _0930_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15404 a_6743_10383# _1086_.Y a_6997_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15406 a_27337_26159# _1887_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15407 vssd1 a_17359_31965# a_17527_31867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15408 vccd1 _1242_.A1 a_5635_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X15410 a_19593_8751# _1152_.B a_19521_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15412 vssd1 a_11711_15831# _1424_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X15414 a_3514_25615# _1761_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15415 a_6921_26159# _1337_.S a_6703_26133# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X15416 vccd1 a_21143_23658# _1833_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15417 _1071_.B1 _1010_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X15418 a_16921_14709# _1090_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X15419 a_19237_14735# a_18703_14741# a_19142_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15422 a_2030_2589# a_1757_2223# a_1945_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15423 vccd1 a_12927_15547# a_12843_15645# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15424 a_24945_15279# _1975_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15425 a_22829_6031# a_22652_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15426 a_24830_15797# a_24662_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15427 a_18182_19203# _1405_.B a_18100_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15428 a_20315_25236# _1416_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15430 a_15921_31433# a_14931_31061# a_15795_31055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15431 vssd1 a_25623_1403# a_25581_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15432 a_13226_5487# _1194_.A2 a_13136_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X15433 a_16293_8751# a_16127_8751# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15434 a_6185_20719# _1327_.A1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X15436 _1138_.C1 a_20267_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15437 vccd1 _1310_.B1 _1310_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X15438 a_9429_15033# _0930_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X15439 vccd1 a_12679_31764# _1473_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15441 vssd1 _1813_.Q a_8945_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15442 vssd1 a_26387_1898# _1651_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15443 a_2309_4943# a_1775_4949# a_2214_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15444 _0921_.A a_2971_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15445 a_23351_7828# _1602_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15446 a_27422_3677# a_26983_3311# a_27337_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15447 _1695_.A a_22103_16733# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15448 vssd1 _1843_.Q a_18329_25981# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15449 clkbuf_0_temp1.i_precharge_n.A a_25695_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15450 a_24662_15823# a_24389_15829# a_24577_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15451 a_20629_3311# a_20359_3677# a_20539_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15452 a_5241_10749# _1234_.A1 a_5169_10749# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15453 vccd1 _1110_.A a_15207_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15454 a_26133_9839# a_25143_9839# a_26007_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15457 a_18969_20175# _0975_.C1 a_18887_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15459 a_14557_10927# a_14287_11293# a_14467_11293# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15460 _1899_.Q a_17895_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15462 vccd1 a_1828_19061# _1260_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X15463 a_3835_2767# a_2971_2773# a_3578_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15464 _1277_.A _1218_.B a_4601_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X15465 a_12736_10761# a_12337_10389# a_12610_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15467 a_18808_4233# a_18409_3861# a_18682_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15468 a_2036_18793# _1311_.B1 a_1781_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X15469 vssd1 _1761_.X a_3514_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15470 vccd1 a_25382_16479# a_25309_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
R34 vccd1 temp1.capload\[7\].cap_52.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X15471 _1732_.X a_22195_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15472 _1968_.Q a_27095_23163# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15473 a_23726_8181# a_23558_8207# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15474 vssd1 a_13599_13866# _1755_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15475 vssd1 a_22015_11471# _1723_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15476 vccd1 _1329_.S a_5664_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X15477 _1329_.S a_8548_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X15480 _1082_.X a_14379_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X15481 a_12601_17277# _1442_.A a_12529_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15482 a_25455_13469# a_24757_13103# a_25198_13215# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15483 a_10585_29423# a_9595_29423# a_10459_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15485 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15486 _1537_.B a_9871_10391# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X15487 _1325_.A2 a_5731_12567# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X15488 vssd1 a_2623_8181# a_2581_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15489 vssd1 _1325_.A2 a_5903_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X15490 a_23155_24349# a_22291_23983# a_22898_24095# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15491 vssd1 a_6151_22869# _1282_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X15493 vccd1 _0916_.A a_3983_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15495 vssd1 _1849_.CLK a_19439_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15496 a_19057_17999# _1821_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15497 a_14979_17130# _1381_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15499 vssd1 a_26099_16911# a_26267_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15501 a_24661_11849# a_23671_11477# a_24535_11471# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15503 vssd1 a_3578_2741# a_3536_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15505 _1513_.A a_20216_22467# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15507 vccd1 a_19275_3829# a_19191_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15508 vssd1 a_24703_10357# a_24661_10761# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15509 vccd1 _1855_.CLK a_10423_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15510 a_10062_25071# _1274_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X15511 _1153_.X a_21279_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15512 a_7599_1501# a_6817_1135# a_7515_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15513 vssd1 a_14123_31029# a_14081_31433# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15514 _1164_.A2 _0930_.A a_8215_8751# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15515 a_5081_19087# _0925_.A2 _1327_.A1_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15516 _0981_.B a_9894_17429# a_9674_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15517 a_24025_4399# a_23848_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15518 vccd1 a_18371_31055# a_18539_31029# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15519 a_5687_4564# _1756_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15520 a_22369_25615# _1833_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15521 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15522 vccd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE a_9595_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X15523 a_19878_29789# a_19605_29423# a_19793_29423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15524 a_6309_3339# _1291_.A1 a_6223_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X15525 a_10693_6575# _1189_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X15526 vccd1 a_2962_14735# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15527 _1099_.B1 a_18243_13760# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15528 vccd1 a_2915_27613# a_3083_27515# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15530 vssd1 a_22063_18218# _1527_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15531 _1050_.Y _1038_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X15532 a_12886_25615# a_12447_25621# a_12801_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15533 vccd1 a_22983_21482# _1885_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15534 a_3312_32143# a_3063_32143# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X15535 a_8387_13647# _0930_.A _1175_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15536 a_24972_3145# a_24573_2773# a_24846_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15537 vssd1 _1459_.A a_16035_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X15539 vccd1 _1786_.A1 a_5727_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X15540 _1143_.X a_14655_18115# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X15541 vccd1 a_1823_19796# _1777_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15542 a_2765_28335# a_1775_28335# a_2639_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15543 a_25769_23439# a_25235_23445# a_25674_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15544 vccd1 _0998_.A2 a_17595_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15545 vccd1 io_in[1] a_2327_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X15547 a_18180_9295# _0993_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X15548 a_18329_25981# a_18059_25615# a_18239_25615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15550 a_25581_28335# a_24591_28335# a_25455_28701# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15551 a_2040_14191# _1218_.B a_1737_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X15554 _1463_.A a_7383_29967# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X15555 a_15013_28111# _1486_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X15556 a_8356_20407# _0913_.A1 a_8498_20214# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X15557 vssd1 a_2623_2491# _1286_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
R35 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X15560 _1896_.CLK a_18830_29967# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15561 a_13061_18543# _1845_.Q a_12989_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15562 _0921_.B a_3983_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15563 vccd1 a_12743_1403# a_12659_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15564 vccd1 a_8307_14191# _1544_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X15565 vccd1 _1816_.CLK a_3983_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15566 a_10386_8181# a_10218_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15567 vssd1 _1042_.B a_12488_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15568 a_20447_9295# a_20267_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15569 _1451_.B a_10811_29941# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15570 _1317_.X a_5087_10496# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15571 vccd1 _1132_.A a_11159_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15572 vssd1 clkbuf_0_net57.X a_2686_26703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15573 vssd1 _1880_.CLK a_22567_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15574 vssd1 _1147_.C1 a_17139_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X15576 vssd1 a_22438_29535# a_22396_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15578 vssd1 a_21150_23007# a_21108_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15579 a_2965_19453# _1762_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X15581 _1304_.B a_2807_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15583 vssd1 a_15207_20719# _1484_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15584 a_5871_1898# _1368_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15585 _0993_.X a_16159_9867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X15586 vssd1 a_2686_26703# temp1.inv2_2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15587 a_2030_9295# a_1757_9301# a_1945_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15588 a_4765_24759# _1763_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X15589 vssd1 _1234_.A2 a_8112_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15590 a_17956_14191# _1033_.A1 a_17381_14337# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X15591 vccd1 _1218_.B a_6682_7913# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X15592 a_7619_26324# _1373_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15593 vssd1 _1184_.X a_15299_20291# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X15594 a_27038_17567# a_26870_17821# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15596 a_26670_25183# a_26502_25437# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X15597 a_27931_10205# a_27149_9839# a_27847_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15599 a_27245_28335# _1886_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15600 a_8120_27791# a_7847_27791# _1775_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15601 a_17313_21807# _0964_.A a_17231_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15603 a_4209_15279# _1323_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X15604 vssd1 _1189_.B2 a_10464_1385# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15605 a_12575_11471# a_11877_11477# a_12318_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15607 _1077_.D1 a_12447_17024# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15608 a_11842_10089# _1139_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X15609 a_4713_12015# _1301_.A1 a_4495_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X15610 temp1.capload\[15\].cap.Y temp1.capload\[15\].cap.A a_22745_32463# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15612 a_1855_22895# _0923_.Y _0925_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X15613 vssd1 a_15917_5461# _1196_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X15614 vssd1 _1148_.B a_6921_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15615 a_18979_10496# _1182_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X15616 _1492_.A a_18607_26525# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X15617 vssd1 a_26927_25437# a_27095_25339# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15618 _1763_.A2 a_2686_23439# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15619 a_1673_20175# _0930_.B _0930_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X15620 _0989_.B2 a_9247_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15621 vccd1 _2023_.CLK a_1775_6037# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15622 vssd1 _1051_.A1 a_10331_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X15624 vssd1 _0983_.A2 a_10677_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X15625 vssd1 _1760_.A_N a_7847_27791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X15626 clkbuf_1_1__f_net57.X a_1674_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15627 a_10862_3677# a_10589_3311# a_10777_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15628 vccd1 _1210_.B a_5303_9633# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X15629 _1859_.Q a_17527_31867# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15631 a_25589_26703# _1883_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15632 a_21647_10205# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15633 a_11306_31711# a_11138_31965# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15635 a_4796_24893# a_4765_24759# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X15636 vccd1 _1270_.A a_5534_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X15637 a_27548_3311# a_27149_3311# a_27422_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15638 a_25800_20553# a_25401_20181# a_25674_20175# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15639 a_2631_13469# a_1849_13103# a_2547_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15640 _1570_.X a_11752_13353# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15641 vccd1 a_2235_2775# _1850_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X15642 vssd1 _1941_.CLK a_18243_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15643 vccd1 _0951_.B a_19439_8751# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X15644 vssd1 a_1827_32117# _1338_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X15646 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE a_11527_28335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15647 a_16274_24095# a_16106_24349# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15648 vccd1 io_in[7] a_1591_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X15649 a_26927_23261# a_26063_22895# a_26670_23007# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15650 a_21235_1898# _1738_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15651 vssd1 _0965_.X a_14839_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X15652 a_21491_23261# a_20709_22895# a_21407_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15653 a_27153_15279# _1389_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15654 _0932_.A a_3247_12672# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15655 vccd1 a_22622_31029# a_22549_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15657 vssd1 _1876_.CLK a_22291_23983# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15661 vssd1 _1344_.Y a_9135_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15663 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15665 _1382_.X a_15616_18115# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X15667 vssd1 _1785_.X a_5812_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15668 a_6469_20719# a_6186_21041# a_6056_20871# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15670 vssd1 a_10811_29941# a_10769_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15671 a_2686_10383# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15672 vccd1 a_22403_30779# a_22319_30877# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15674 vccd1 a_27479_16733# a_27647_16635# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15675 vccd1 a_2198_2335# a_2125_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15676 vssd1 _1941_.CLK a_17507_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15677 _1291_.A1 a_2623_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15678 vccd1 _1924_.CLK a_23119_8213# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15679 vssd1 _1077_.X a_14379_18793# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X15680 a_13993_24527# a_13459_24533# a_13898_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15681 a_26597_23261# a_26063_22895# a_26502_23261# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15682 vccd1 _1326_.A2 a_4533_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X15683 vccd1 _1041_.A1 a_20907_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15684 a_13057_8897# _1059_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X15685 a_19952_12533# _1183_.B1 a_20081_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X15686 _1387_.A a_23391_16733# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X15687 vssd1 a_17831_11092# _1584_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15688 vssd1 a_23726_8181# a_23684_8585# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15689 _2023_.CLK a_2686_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X15690 vccd1 _1590_.A_N a_17047_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15691 vccd1 _1218_.B _1301_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15692 vccd1 _1782_.A a_6651_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15693 a_23523_9117# a_22825_8751# a_23266_8863# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15694 vccd1 _1301_.A1 _1246_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15695 a_6743_10703# _1298_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15696 a_22081_13621# _1190_.B1 a_22238_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X15697 vccd1 _1965_.Q a_22747_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15698 vccd1 _1324_.A a_6743_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15699 vccd1 a_12035_2986# _1934_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15701 a_2639_4765# a_1941_4399# a_2382_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15702 a_9043_21263# _1544_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15703 vssd1 _1184_.A2 a_19877_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X15704 _1074_.X a_16863_21376# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15705 vccd1 a_10995_19899# a_10911_19997# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15706 a_17257_16395# _0961_.A a_17171_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X15707 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A a_3312_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15708 a_26670_23007# a_26502_23261# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15709 a_11865_15101# _1905_.Q a_11793_15101# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15712 a_13275_32143# _1474_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15713 vssd1 _1882_.CLK a_26799_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15714 vssd1 _1269_.A1 _0981_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15717 a_11877_29423# a_11711_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15718 a_25539_28701# a_24757_28335# a_25455_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15720 a_24661_10761# a_23671_10389# a_24535_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15721 vssd1 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE a_6559_31599# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15722 a_19793_31599# _1540_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15724 a_25306_11293# a_25033_10927# a_25221_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15726 a_14453_9839# a_14287_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15727 vssd1 a_10459_29789# a_10627_29691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15728 vssd1 _1066_.B a_17317_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15729 a_27903_16911# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15730 a_13165_13103# _1219_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15731 vssd1 a_13330_29941# a_13288_30345# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15732 _1132_.C a_10865_18909# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X15733 a_24021_1685# a_23855_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15734 a_18703_27791# _0965_.B1 a_18785_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15735 a_19237_1679# a_18703_1685# a_19142_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15736 vssd1 _1129_.B a_23849_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15738 vssd1 a_2991_25339# _2005_.Q vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15740 vssd1 a_9937_4917# _1011_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X15741 vccd1 a_20782_4511# a_20709_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15742 a_3041_27247# a_2051_27247# a_2915_27613# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15743 _1689_.A a_21091_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15744 a_18313_29257# a_17323_28885# a_18187_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15745 _0923_.Y _1775_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15747 a_7843_8207# a_7663_8207# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15748 vccd1 _1263_.A _1265_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15749 a_15538_25589# a_15370_25615# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15750 vssd1 a_1674_30511# clkbuf_1_1__f_net57.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15751 a_25769_22351# a_25235_22357# a_25674_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15752 a_6867_8545# _1165_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X15756 vccd1 a_20655_28603# a_20571_28701# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15757 vssd1 a_2715_13371# _1218_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15758 vssd1 a_23523_27613# a_23691_27515# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15759 vccd1 a_2639_7119# a_2807_7093# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15761 vccd1 _1307_.X a_4150_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X15762 a_15931_15823# _1034_.D _1034_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15763 a_23903_19796# _1387_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15765 vccd1 _1141_.C a_17415_13760# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X15766 vssd1 a_23303_6031# fanout20.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15767 a_22825_3311# a_22659_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15768 vccd1 a_27463_6843# a_27379_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15769 a_13805_11471# _1143_.X a_13551_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15770 a_10083_7119# a_9301_7125# a_9999_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15771 a_6797_19605# _1325_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X15772 vccd1 _1232_.Y a_4161_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X15773 a_24941_17999# a_24407_18005# a_24846_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15774 _1717_.X a_23667_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X15775 vccd1 _1760_.B a_2309_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X15776 a_2850_15279# _1301_.A1 a_2472_15431# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X15777 _1061_.B a_27739_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15778 _1110_.A a_14103_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X15779 vccd1 a_20379_31029# a_20295_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15780 _1881_.Q a_26175_26427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15781 a_20161_32143# _1896_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15782 _0913_.Y _1242_.B1 a_5455_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15783 vccd1 a_3467_24527# a_3635_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15784 a_5099_24527# _1766_.A0 a_4587_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X15785 _1421_.A a_12396_22057# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15786 _1727_.X a_23483_12381# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15787 a_20387_31965# a_19605_31599# a_20303_31965# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15788 a_2781_21807# _1237_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X15789 vccd1 _1855_.CLK a_9779_29973# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15790 vssd1 a_25455_28701# a_25623_28603# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15792 vssd1 a_3467_24527# a_3635_24501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15793 a_22879_24527# a_22015_24533# a_22622_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15794 _1269_.B1 a_4351_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X15795 a_6717_9001# _1122_.A1 a_6645_9001# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15796 vccd1 _1324_.A _1326_.A3 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15797 vssd1 _1824_.Q a_23573_16189# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15799 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE a_7387_32143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X15800 vssd1 a_23967_3829# a_23925_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15801 vccd1 a_25639_3855# a_25807_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15802 _1084_.C1 a_1626_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X15803 a_25455_2589# a_24757_2223# a_25198_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15804 a_27571_2589# a_26873_2223# a_27314_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15805 vssd1 a_28135_13866# _1975_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15806 vssd1 a_20303_1501# a_20471_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15807 vssd1 a_7867_3829# a_7825_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15808 vssd1 a_12575_8207# a_12743_8181# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15809 temp1.capload\[15\].cap.B a_10506_30511# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15810 a_13544_30511# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X15811 a_14776_24233# _1056_.B1 a_14674_24233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X15812 _0965_.A2 a_16159_20747# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X15813 temp1.inv2_2.Y temp1.inv2_2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15814 a_6641_16189# _1273_.A1 a_6559_15936# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15815 vccd1 a_17647_2388# _1944_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15818 a_1791_13967# _1246_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X15819 a_7737_28335# _1273_.A1 _1274_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X15821 vssd1 _0930_.A a_6747_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X15823 _1122_.A1 _1120_.X a_9779_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15824 a_22549_24527# a_22015_24533# a_22454_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15825 vssd1 _1394_.A a_18100_19203# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X15826 vccd1 _1744_.A_N a_23579_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15827 a_17861_32143# _1841_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X15828 a_5177_14191# _1217_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X15829 a_20947_11471# a_20249_11477# a_20690_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15830 _1205_.A1 a_3063_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15832 vccd1 _0918_.A a_6929_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X15833 vssd1 a_27590_3423# a_27548_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X15834 a_27675_29588# _1463_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15835 vssd1 _1242_.B1 _1306_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15836 a_7442_17429# _1269_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X15837 a_2125_2589# a_1591_2223# a_2030_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15838 vssd1 _1032_.C a_19041_19453# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X15839 vccd1 _0939_.A a_21463_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15840 vccd1 _1015_.A1 a_10603_9117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X15841 a_17170_26819# _1484_.B a_17088_26819# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15842 _1303_.A1 a_4443_20175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X15843 vccd1 a_25455_17821# a_25623_17723# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15844 a_26295_18218# _1693_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15845 a_21003_2767# _1744_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15846 _1684_.A a_22747_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15847 vccd1 a_10459_2589# a_10627_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15848 vccd1 a_25455_9117# a_25623_9019# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15849 vccd1 a_2198_9269# a_2125_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X15850 a_17727_17999# a_17029_18005# a_17470_17973# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15852 vccd1 a_4863_23413# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15853 vccd1 _1249_.A2 a_4719_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15854 a_20911_24349# _1489_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15855 _1761_.X a_27167_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X15856 _1657_.A a_7199_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X15857 a_14545_4949# a_14379_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15858 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE a_7479_28887# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X15859 a_15545_8573# _1109_.B a_15473_8573# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X15860 _1872_.Q a_22403_30779# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15861 vssd1 _1882_.CLK a_25235_22357# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15862 a_14921_25071# _1132_.A a_14839_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15863 _0963_.B a_12226_16341# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X15864 a_12659_8207# a_11877_8213# a_12575_8207# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15865 clkbuf_1_1__f_net57.X a_1674_30511# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15867 vccd1 a_5417_18517# _1254_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15868 a_19487_4564# _1636_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15869 vssd1 a_20303_31965# a_20471_31867# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15871 a_20065_13647# _1191_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X15873 vssd1 a_26175_10107# a_26133_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15875 vccd1 a_3514_25615# clkbuf_1_1__f__0380_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15876 a_25585_18543# a_25419_18543# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15877 a_27399_16042# _1700_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X15878 vssd1 a_11455_3579# a_11413_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15882 vccd1 a_12557_16600# a_12226_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X15883 vccd1 _1267_.A1 a_3707_6144# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15885 a_22383_12381# _1685_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X15886 vssd1 _1768_.A _1074_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15887 a_2225_17455# _1250_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X15888 vccd1 _1127_.A a_16035_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15889 a_25581_20719# a_24591_20719# a_25455_21085# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15891 vccd1 a_27847_12381# a_28015_12283# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15892 vccd1 fanout33.A a_15667_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15893 vssd1 _1242_.B1 _1274_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X15894 a_22825_21807# a_22659_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15895 vssd1 a_24903_19087# a_25071_19061# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15896 vccd1 a_18171_29691# a_18087_29789# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15898 vccd1 _1269_.A1 a_10938_16341# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X15899 vccd1 _1590_.A_N a_16127_6941# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X15901 _1071_.B1 _0987_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15902 vssd1 a_2686_10383# _2023_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15903 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE a_9963_32143# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X15904 _1860_.CLK a_9779_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X15905 _1013_.X a_10648_12675# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15907 a_27421_13103# a_26431_13103# a_27295_13469# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X15908 a_12065_29423# _1902_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X15909 a_23573_16189# a_23303_15823# a_23483_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X15911 vccd1 a_23443_7338# _1676_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15912 vccd1 a_5233_11445# _1796_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X15915 a_17428_30345# a_17029_29973# a_17302_29967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X15916 a_10593_22057# _0921_.B a_10951_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15917 a_27406_15391# a_27238_15645# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15919 vssd1 a_15319_30779# a_15277_30511# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15920 vssd1 a_25623_15547# a_25581_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15921 _1154_.C1 a_19439_8751# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X15922 a_3467_24527# a_2603_24533# a_3210_24501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15923 vccd1 a_8454_15797# _1047_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X15924 a_25030_24349# a_24757_23983# a_24945_23983# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15926 vccd1 _0966_.A2 a_15833_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X15927 vccd1 _1882_.CLK a_26799_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15928 a_12334_4943# a_12061_4949# a_12249_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15929 _1473_.A a_14144_27907# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15930 a_3276_20495# _1257_.B1 a_3185_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X15931 vccd1 a_10506_30511# temp1.capload\[15\].cap.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15932 _0987_.Y _0987_.B a_11067_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15933 vssd1 a_20471_5755# a_20429_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15934 _1191_.A1 a_27923_11195# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15937 _1436_.B a_12743_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15938 _1875_.Q a_21115_27765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15940 vssd1 _1098_.B a_16397_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15941 vccd1 _1816_.CLK a_8215_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15943 vssd1 _1269_.A1 _1766_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15944 a_11793_21263# _1856_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X15945 vssd1 a_15633_19061# _1020_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X15947 a_16616_14441# _1024_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X15948 _1242_.A2 a_7111_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X15949 a_3137_24527# a_2603_24533# a_3042_24527# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15950 a_2331_12879# _1246_.B2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X15951 a_7001_3861# a_6835_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15952 _1436_.B a_12743_11445# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15954 a_27755_11293# a_26891_10927# a_27498_11039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X15955 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z a_17388_27497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X15956 vssd1 _1873_.Q a_18697_26159# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X15957 vssd1 a_27095_23163# a_27053_22895# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15958 a_18969_20175# _1184_.B1 a_19053_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15959 vssd1 a_25255_15797# a_25213_16201# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X15960 vccd1 _1127_.A a_20267_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15961 a_17630_14441# _1032_.X a_17381_14337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X15962 vssd1 a_18107_14954# _1914_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15963 _1074_.C _1764_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15964 a_10596_9839# _1011_.A1 a_10021_9985# vssd1 sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X15965 a_23818_16885# a_23650_16911# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15966 vccd1 _1353_.B a_11711_27791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X15967 a_24075_16911# a_23377_16917# a_23818_16885# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X15968 a_26965_17821# a_26431_17455# a_26870_17821# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X15969 a_20982_8029# a_20709_7663# a_20897_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X15970 a_10140_32463# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X15971 temp1.capload\[9\].cap.Y temp1.capload\[9\].cap.A a_23757_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15972 vssd1 _1330_.X a_21371_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X15973 vssd1 a_10423_23983# _1270_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15974 a_19836_15823# _1127_.X a_19734_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X15975 vssd1 a_5731_7127# _1448_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X15976 a_16904_22467# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15977 a_23759_5853# a_23579_5853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X15978 a_3789_6397# _1267_.A1 a_3707_6144# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15979 vssd1 a_15750_28335# temp1.capload\[6\].cap.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15981 _1529_.A a_20860_19881# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X15982 vccd1 a_10931_2986# _1612_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X15983 vccd1 _1999_.CLK a_9135_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X15985 vccd1 a_2639_6031# a_2807_6005# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X15986 a_14369_17455# _1132_.A a_14287_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X15988 a_21905_5487# a_21739_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15989 vssd1 a_20671_32143# a_20839_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15990 a_10951_22057# _0921_.B a_10593_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15991 vssd1 a_2686_15823# _2009_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X15992 _1506_.B a_18611_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X15993 vccd1 _1021_.A a_13091_19200# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X15995 _1032_.X a_18887_19200# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X15997 a_20522_28879# a_20083_28885# a_20437_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X15998 vccd1 a_24243_23413# a_24159_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X15999 vccd1 _1970_.Q a_22103_16733# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X16000 vssd1 a_20591_1898# _1940_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X16001 _1540_.A a_14927_28701# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X16002 a_23667_17999# a_23487_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X16004 a_15879_25615# a_15097_25621# a_15795_25615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X16005 a_5871_23658# _1375_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16006 vssd1 _1090_.C a_16797_15307# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X16007 vccd1 a_28015_3579# a_27931_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X16008 vccd1 a_1657_10901# _1177_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X16009 a_11803_6575# _1117_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X16010 a_27237_14191# a_26247_14191# a_27111_14557# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X16011 vccd1 a_25623_13371# a_25539_13469# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X16012 vccd1 a_7619_2986# _1955_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X16013 a_7928_27023# _1261_.A1 a_7625_26677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X16014 vccd1 _1544_.A_N a_7755_22351# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X16015 a_12927_13103# _1219_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X16017 a_10283_25071# _1306_.A2 a_9920_25223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X16018 a_18836_23555# _1405_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16019 vssd1 fanout20.X a_25235_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16020 a_2413_29423# a_2143_29789# a_2309_29789# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X16023 a_2125_9295# a_1591_9301# a_2030_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X16025 _1142_.B1 a_10055_21376# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X16026 _1053_.A _2007_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X16027 _1030_.B a_14307_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16028 vccd1 a_5509_17973# _1786_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X16030 vccd1 a_7975_2589# a_8143_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X16031 vccd1 _1047_.C a_12907_7232# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X16032 clkbuf_1_1__f__0380_.A a_3514_25615# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16034 vccd1 a_1674_30511# clkbuf_1_1__f_net57.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X16035 vccd1 _1394_.A a_18182_19203# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X16037 a_17415_3677# _1639_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16038 vssd1 a_18371_32143# a_18539_32117# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16039 vssd1 a_19567_14735# a_19735_14709# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16040 a_27364_21807# a_26965_21807# a_27238_22173# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X16041 vssd1 _1823_.Q a_23481_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X16042 _1044_.X a_11159_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X16043 vssd1 a_24646_19061# a_24604_19465# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X16044 a_4590_1653# a_4422_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X16045 a_26226_4765# a_25787_4399# a_26141_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X16046 vccd1 a_12815_6031# _1639_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16048 _0994_.B2 a_18539_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16051 vssd1 _1882_.CLK a_23211_23445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16052 vccd1 a_11030_27359# a_10957_27613# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X16053 vccd1 a_14370_31599# clkbuf_0_temp1.dcdel_capnode_notouch_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16054 _1877_.Q a_25991_22075# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16057 _1134_.B1 a_15483_23552# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X16058 io_out[1] a_1643_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16059 a_9735_9514# _1759_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X16060 a_17861_31055# _1467_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X16065 a_18697_26159# a_18427_26525# a_18607_26525# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X16066 vccd1 _1205_.Y a_4015_8779# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X16067 _1329_.A0 a_1674_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16069 a_5241_13647# _1217_.B1 a_4709_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X16070 a_16029_29245# a_15759_28879# a_15939_28879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X16071 vssd1 _1855_.CLK a_10423_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16072 _1654_.X a_6739_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X16073 _1880_.CLK a_15886_25071# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X16074 a_20131_21972# _1523_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X16075 a_25823_22173# a_24959_21807# a_25566_21919# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16076 vccd1 a_7295_6031# _1177_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X16077 a_9489_31055# _1860_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X16078 a_18107_21972# _1397_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16079 vssd1 a_22081_14709# _1190_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X16080 a_6808_29673# a_6559_29423# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X16081 vssd1 a_13311_25615# a_13479_25589# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16082 vccd1 a_15115_5487# _1830_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16083 a_23013_8751# _1920_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X16084 a_5629_12015# _1291_.A1 a_5547_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X16085 vssd1 fanout28.A a_16311_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X16086 a_9761_2223# a_9595_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X16087 vccd1 a_23627_6740# _1593_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X16088 a_15089_10499# _1008_.B a_15017_10499# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X16090 vccd1 _1269_.A1 a_7479_17277# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X16091 a_16434_14441# _1099_.D1 a_16185_14337# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X16092 vssd1 _1192_.X a_14287_9001# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X16093 vccd1 _1723_.A_N a_23303_12381# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X16094 a_11983_18909# a_11803_18909# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X16095 a_13173_19453# _1021_.A a_13091_19200# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X16096 a_22879_2767# a_22181_2773# a_22622_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X16097 a_1643_21237# _1260_.B1 a_2706_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16098 a_22707_18218# _1500_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16099 vccd1 _1459_.A a_17047_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X16100 vccd1 _1353_.Y a_8158_29967# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X16101 _1133_.X a_17415_24640# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X16102 vccd1 a_20885_16341# _1179_.C1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X16103 a_14545_3861# a_14379_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X16104 a_19878_29789# a_19439_29423# a_19793_29423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X16105 vccd1 a_10839_10602# _1848_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X16106 a_7019_12265# _1086_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16107 a_19881_31055# a_19347_31061# a_19786_31055# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X16109 vssd1 _1047_.C a_12601_17277# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X16110 _1205_.Y _1170_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X16111 vccd1 _1841_.CLK a_17323_28885# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X16112 a_25493_22173# a_24959_21807# a_25398_22173# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X16113 a_5911_19881# _1780_.B1 a_5693_19605# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X16114 a_10865_18909# a_10699_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X16115 _1012_.Y _1012_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16116 a_17812_7119# _1061_.X a_17710_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X16117 _1590_.A_N a_16035_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X16118 a_11895_19631# _1819_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X16119 _1249_.A2 a_2472_15431# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X16120 a_26225_12937# a_25235_12565# a_26099_12559# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X16122 a_12027_20495# _0956_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X16123 vccd1 _1286_.A1 a_6559_26703# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16124 _1500_.A a_20999_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X16125 _1813_.Q a_10811_8181# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16126 a_22825_21807# a_22659_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X16127 vssd1 a_13551_17999# _0958_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16128 vccd1 _1985_.CLK a_26799_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X16129 a_5625_5792# _1780_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16130 _1393_.A a_18560_18793# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X16131 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16132 _1184_.A2 a_17723_20513# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X16134 a_4931_25437# a_4149_25071# a_4847_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X16135 _1070_.X a_17139_18793# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X16136 a_17276_6351# _1047_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X16137 a_23473_8207# _1916_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X16138 vccd1 _0951_.B a_17541_15307# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X16140 a_10643_8207# a_9779_8213# a_10386_8181# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16141 vssd1 _1047_.C a_15693_12043# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X16142 a_4351_12879# _1217_.A3 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16143 a_17930_28853# a_17762_28879# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X16144 a_20617_28879# a_20083_28885# a_20522_28879# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X16147 vccd1 _1032_.C a_17139_11584# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X16148 vssd1 a_27215_17130# _1389_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X16150 vccd1 _1121_.A1 a_10227_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16151 _1867_.Q a_17895_29941# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16152 temp1.capload\[6\].cap.B a_15750_28335# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16153 vccd1 _1885_.Q a_19928_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X16154 a_22730_18909# a_22291_18543# a_22645_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X16155 a_11023_26922# _1458_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16156 a_22733_20175# a_22199_20181# a_22638_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X16157 _1359_.X a_8395_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X16158 vssd1 _1353_.A _1344_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16159 vssd1 _2009_.CLK a_3983_25071# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16162 vccd1 temp1.capload\[13\].cap_43.LO temp1.capload\[13\].cap.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16163 vccd1 _1073_.A2 a_16301_22057# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X16164 a_23487_17999# _1690_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16165 vssd1 _1797_.Y a_5817_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X16166 vccd1 a_26670_25183# a_26597_25437# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X16167 a_18371_32143# a_17507_32149# a_18114_32117# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16168 vssd1 a_25455_21085# a_25623_20987# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16170 vccd1 _1194_.A2 a_13490_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X16171 a_14741_1135# a_14471_1501# a_14651_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X16172 a_20249_11477# a_20083_11477# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X16173 a_3881_16911# _1291_.B1 a_3965_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16174 a_22546_6031# a_22369_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X16176 a_18085_16395# _0961_.A a_17999_16395# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X16177 a_4263_22895# _1274_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X16178 a_9602_25654# _1329_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X16179 vccd1 a_2686_26703# temp1.inv2_2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16180 _1118_.X a_17139_11584# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X16182 a_25306_11293# a_24867_10927# a_25221_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X16183 vssd1 a_27295_13469# a_27463_13371# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16186 vccd1 a_22879_1679# a_23047_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X16188 a_20211_31055# a_19513_31061# a_19954_31029# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X16190 a_17470_27765# a_17302_27791# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X16191 clkbuf_1_1__f_io_in[0].A a_2962_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16192 a_18243_13760# _1721_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X16193 _1179_.B2 a_21115_11445# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16194 vccd1 a_17470_17973# a_17397_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X16195 a_18170_17705# _1049_.C1 a_18090_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X16196 vssd1 _0963_.B a_13061_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X16197 vccd1 a_7295_17455# a_7442_17429# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X16199 a_26295_2986# _1318_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16200 a_9503_16911# _1768_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 a_24945_1135# vssd1 0.23fF $ **FLOATING
C1 a_27215_1300# vssd1 0.52fF $ **FLOATING
C2 a_26479_1300# vssd1 0.52fF $ **FLOATING
C3 a_25455_1501# vssd1 0.61fF $ **FLOATING
C4 a_25623_1403# vssd1 0.82fF $ **FLOATING
C5 a_25030_1501# vssd1 0.63fF $ **FLOATING
C6 a_25198_1247# vssd1 0.58fF $ **FLOATING
C7 a_24757_1135# vssd1 1.43fF $ **FLOATING
C8 a_24591_1135# vssd1 1.81fF $ **FLOATING
C9 a_22369_1135# vssd1 0.23fF $ **FLOATING
C10 a_23903_1300# vssd1 0.52fF $ **FLOATING
C11 a_22879_1501# vssd1 0.61fF $ **FLOATING
C12 a_23047_1403# vssd1 0.82fF $ **FLOATING
C13 a_22454_1501# vssd1 0.63fF $ **FLOATING
C14 a_22622_1247# vssd1 0.58fF $ **FLOATING
C15 a_22181_1135# vssd1 1.43fF $ **FLOATING
C16 a_22015_1135# vssd1 1.81fF $ **FLOATING
C17 a_19793_1135# vssd1 0.23fF $ **FLOATING
C18 a_21327_1300# vssd1 0.52fF $ **FLOATING
C19 a_20303_1501# vssd1 0.61fF $ **FLOATING
C20 a_20471_1403# vssd1 0.82fF $ **FLOATING
C21 a_19878_1501# vssd1 0.63fF $ **FLOATING
C22 a_20046_1247# vssd1 0.58fF $ **FLOATING
C23 a_19605_1135# vssd1 1.43fF $ **FLOATING
C24 a_19439_1135# vssd1 1.81fF $ **FLOATING
C25 a_17861_1135# vssd1 0.23fF $ **FLOATING
C26 a_18371_1501# vssd1 0.61fF $ **FLOATING
C27 a_18539_1403# vssd1 0.82fF $ **FLOATING
C28 a_17946_1501# vssd1 0.63fF $ **FLOATING
C29 a_18114_1247# vssd1 0.58fF $ **FLOATING
C30 a_17673_1135# vssd1 1.43fF $ **FLOATING
C31 a_17507_1135# vssd1 1.81fF $ **FLOATING
C32 _1945_.D vssd1 1.92fF $ **FLOATING
C33 a_12065_1135# vssd1 0.23fF $ **FLOATING
C34 a_16911_1300# vssd1 0.52fF $ **FLOATING
C35 a_15432_1385# vssd1 0.50fF $ **FLOATING
C36 a_14651_1501# vssd1 0.51fF $ **FLOATING
C37 a_14471_1501# vssd1 0.60fF $ **FLOATING
C38 _1645_.A vssd1 1.14fF $ **FLOATING
C39 a_13599_1300# vssd1 0.52fF $ **FLOATING
C40 a_12575_1501# vssd1 0.61fF $ **FLOATING
C41 a_12743_1403# vssd1 0.82fF $ **FLOATING
C42 a_12150_1501# vssd1 0.63fF $ **FLOATING
C43 a_12318_1247# vssd1 0.58fF $ **FLOATING
C44 a_11877_1135# vssd1 1.43fF $ **FLOATING
C45 a_11711_1135# vssd1 1.81fF $ **FLOATING
C46 _1616_.A vssd1 8.11fF $ **FLOATING
C47 a_7005_1135# vssd1 0.23fF $ **FLOATING
C48 a_10464_1385# vssd1 0.50fF $ **FLOATING
C49 a_9683_1501# vssd1 0.51fF $ **FLOATING
C50 a_9503_1501# vssd1 0.60fF $ **FLOATING
C51 a_7515_1501# vssd1 0.61fF $ **FLOATING
C52 a_7683_1403# vssd1 0.82fF $ **FLOATING
C53 a_7090_1501# vssd1 0.63fF $ **FLOATING
C54 a_7258_1247# vssd1 0.58fF $ **FLOATING
C55 a_6817_1135# vssd1 1.43fF $ **FLOATING
C56 a_6651_1135# vssd1 1.81fF $ **FLOATING
C57 a_4521_1135# vssd1 0.23fF $ **FLOATING
C58 a_5031_1501# vssd1 0.61fF $ **FLOATING
C59 a_5199_1403# vssd1 0.82fF $ **FLOATING
C60 a_4606_1501# vssd1 0.63fF $ **FLOATING
C61 a_4774_1247# vssd1 0.58fF $ **FLOATING
C62 a_4333_1135# vssd1 1.43fF $ **FLOATING
C63 a_4167_1135# vssd1 1.81fF $ **FLOATING
C64 a_1945_1135# vssd1 0.23fF $ **FLOATING
C65 a_2455_1501# vssd1 0.61fF $ **FLOATING
C66 a_2623_1403# vssd1 0.82fF $ **FLOATING
C67 a_2030_1501# vssd1 0.63fF $ **FLOATING
C68 a_2198_1247# vssd1 0.58fF $ **FLOATING
C69 a_1757_1135# vssd1 1.43fF $ **FLOATING
C70 a_1591_1135# vssd1 1.81fF $ **FLOATING
C71 a_24209_1679# vssd1 0.23fF $ **FLOATING
C72 a_22369_1679# vssd1 0.23fF $ **FLOATING
C73 a_19057_1679# vssd1 0.23fF $ **FLOATING
C74 a_17217_1679# vssd1 0.23fF $ **FLOATING
C75 _1957_.D vssd1 3.78fF $ **FLOATING
C76 a_13629_1679# vssd1 0.23fF $ **FLOATING
C77 _1956_.D vssd1 3.61fF $ **FLOATING
C78 a_10133_1679# vssd1 0.23fF $ **FLOATING
C79 a_8293_1679# vssd1 0.23fF $ **FLOATING
C80 a_4337_1679# vssd1 0.23fF $ **FLOATING
C81 a_2497_1679# vssd1 0.23fF $ **FLOATING
C82 a_26387_1898# vssd1 0.52fF $ **FLOATING
C83 a_25743_1898# vssd1 0.52fF $ **FLOATING
C84 a_24719_1679# vssd1 0.61fF $ **FLOATING
C85 a_24887_1653# vssd1 0.82fF $ **FLOATING
C86 a_24294_1679# vssd1 0.63fF $ **FLOATING
C87 a_24462_1653# vssd1 0.58fF $ **FLOATING
C88 a_24021_1685# vssd1 1.43fF $ **FLOATING
C89 a_23855_1685# vssd1 1.81fF $ **FLOATING
C90 a_22879_1679# vssd1 0.61fF $ **FLOATING
C91 a_23047_1653# vssd1 0.82fF $ **FLOATING
C92 a_22454_1679# vssd1 0.63fF $ **FLOATING
C93 a_22622_1653# vssd1 0.58fF $ **FLOATING
C94 a_22181_1685# vssd1 1.43fF $ **FLOATING
C95 _1940_.D vssd1 1.51fF $ **FLOATING
C96 a_22015_1685# vssd1 1.81fF $ **FLOATING
C97 a_21235_1898# vssd1 0.52fF $ **FLOATING
C98 a_20591_1898# vssd1 0.52fF $ **FLOATING
C99 a_19567_1679# vssd1 0.61fF $ **FLOATING
C100 a_19735_1653# vssd1 0.82fF $ **FLOATING
C101 a_19142_1679# vssd1 0.63fF $ **FLOATING
C102 a_19310_1653# vssd1 0.58fF $ **FLOATING
C103 a_18869_1685# vssd1 1.43fF $ **FLOATING
C104 a_18703_1685# vssd1 1.81fF $ **FLOATING
C105 a_17727_1679# vssd1 0.61fF $ **FLOATING
C106 a_17895_1653# vssd1 0.82fF $ **FLOATING
C107 a_17302_1679# vssd1 0.63fF $ **FLOATING
C108 a_17470_1653# vssd1 0.58fF $ **FLOATING
C109 a_17029_1685# vssd1 1.43fF $ **FLOATING
C110 a_16863_1685# vssd1 1.81fF $ **FLOATING
C111 _1665_.A vssd1 0.88fF $ **FLOATING
C112 a_16175_1898# vssd1 0.52fF $ **FLOATING
C113 a_15387_1679# vssd1 0.51fF $ **FLOATING
C114 a_15207_1679# vssd1 0.60fF $ **FLOATING
C115 a_14139_1679# vssd1 0.61fF $ **FLOATING
C116 a_14307_1653# vssd1 0.82fF $ **FLOATING
C117 a_13714_1679# vssd1 0.63fF $ **FLOATING
C118 a_13882_1653# vssd1 0.58fF $ **FLOATING
C119 a_13441_1685# vssd1 1.43fF $ **FLOATING
C120 a_13275_1685# vssd1 1.81fF $ **FLOATING
C121 a_12535_1679# vssd1 0.51fF $ **FLOATING
C122 a_12355_1679# vssd1 0.60fF $ **FLOATING
C123 _1662_.X vssd1 1.00fF $ **FLOATING
C124 a_11759_1898# vssd1 0.52fF $ **FLOATING
C125 a_10643_1679# vssd1 0.61fF $ **FLOATING
C126 a_10811_1653# vssd1 0.82fF $ **FLOATING
C127 a_10218_1679# vssd1 0.63fF $ **FLOATING
C128 a_10386_1653# vssd1 0.58fF $ **FLOATING
C129 a_9945_1685# vssd1 1.43fF $ **FLOATING
C130 _1616_.X vssd1 8.32fF $ **FLOATING
C131 a_9779_1685# vssd1 1.81fF $ **FLOATING
C132 a_8803_1679# vssd1 0.61fF $ **FLOATING
C133 a_8971_1653# vssd1 0.82fF $ **FLOATING
C134 a_8378_1679# vssd1 0.63fF $ **FLOATING
C135 a_8546_1653# vssd1 0.58fF $ **FLOATING
C136 a_8105_1685# vssd1 1.43fF $ **FLOATING
C137 a_7939_1685# vssd1 1.81fF $ **FLOATING
C138 a_7199_1679# vssd1 0.51fF $ **FLOATING
C139 a_7019_1679# vssd1 0.60fF $ **FLOATING
C140 a_5871_1898# vssd1 0.52fF $ **FLOATING
C141 a_4847_1679# vssd1 0.61fF $ **FLOATING
C142 a_5015_1653# vssd1 0.82fF $ **FLOATING
C143 a_4422_1679# vssd1 0.63fF $ **FLOATING
C144 a_4590_1653# vssd1 0.58fF $ **FLOATING
C145 a_4149_1685# vssd1 1.43fF $ **FLOATING
C146 a_3983_1685# vssd1 1.81fF $ **FLOATING
C147 a_3007_1679# vssd1 0.61fF $ **FLOATING
C148 a_3175_1653# vssd1 0.82fF $ **FLOATING
C149 a_2582_1679# vssd1 0.63fF $ **FLOATING
C150 a_2750_1653# vssd1 0.58fF $ **FLOATING
C151 a_2309_1685# vssd1 1.43fF $ **FLOATING
C152 _1651_.X vssd1 11.22fF $ **FLOATING
C153 a_2143_1685# vssd1 1.81fF $ **FLOATING
C154 a_27061_2223# vssd1 0.23fF $ **FLOATING
C155 a_27571_2589# vssd1 0.61fF $ **FLOATING
C156 a_27739_2491# vssd1 0.82fF $ **FLOATING
C157 a_27146_2589# vssd1 0.63fF $ **FLOATING
C158 a_27314_2335# vssd1 0.58fF $ **FLOATING
C159 a_26873_2223# vssd1 1.43fF $ **FLOATING
C160 a_26707_2223# vssd1 1.81fF $ **FLOATING
C161 a_24945_2223# vssd1 0.23fF $ **FLOATING
C162 a_25455_2589# vssd1 0.61fF $ **FLOATING
C163 a_25623_2491# vssd1 0.82fF $ **FLOATING
C164 a_25030_2589# vssd1 0.63fF $ **FLOATING
C165 a_25198_2335# vssd1 0.58fF $ **FLOATING
C166 a_24757_2223# vssd1 1.43fF $ **FLOATING
C167 a_24591_2223# vssd1 1.81fF $ **FLOATING
C168 a_23013_2223# vssd1 0.23fF $ **FLOATING
C169 a_23523_2589# vssd1 0.61fF $ **FLOATING
C170 a_23691_2491# vssd1 0.82fF $ **FLOATING
C171 a_23098_2589# vssd1 0.63fF $ **FLOATING
C172 a_23266_2335# vssd1 0.58fF $ **FLOATING
C173 a_22825_2223# vssd1 1.43fF $ **FLOATING
C174 a_22659_2223# vssd1 1.81fF $ **FLOATING
C175 a_20897_2223# vssd1 0.23fF $ **FLOATING
C176 a_21407_2589# vssd1 0.61fF $ **FLOATING
C177 a_21575_2491# vssd1 0.82fF $ **FLOATING
C178 a_20982_2589# vssd1 0.63fF $ **FLOATING
C179 a_21150_2335# vssd1 0.58fF $ **FLOATING
C180 a_20709_2223# vssd1 1.43fF $ **FLOATING
C181 a_20543_2223# vssd1 1.81fF $ **FLOATING
C182 _1628_.X vssd1 3.69fF $ **FLOATING
C183 _1944_.D vssd1 2.09fF $ **FLOATING
C184 a_16113_2223# vssd1 0.23fF $ **FLOATING
C185 a_19487_2388# vssd1 0.52fF $ **FLOATING
C186 _1628_.A vssd1 2.35fF $ **FLOATING
C187 a_18291_2388# vssd1 0.52fF $ **FLOATING
C188 a_17647_2388# vssd1 0.52fF $ **FLOATING
C189 a_16623_2589# vssd1 0.61fF $ **FLOATING
C190 a_16791_2491# vssd1 0.82fF $ **FLOATING
C191 a_16198_2589# vssd1 0.63fF $ **FLOATING
C192 a_16366_2335# vssd1 0.58fF $ **FLOATING
C193 a_15925_2223# vssd1 1.43fF $ **FLOATING
C194 _1947_.D vssd1 2.37fF $ **FLOATING
C195 a_15759_2223# vssd1 1.81fF $ **FLOATING
C196 _1643_.X vssd1 2.54fF $ **FLOATING
C197 a_11789_2223# vssd1 0.23fF $ **FLOATING
C198 a_15163_2388# vssd1 0.52fF $ **FLOATING
C199 a_14335_2388# vssd1 0.52fF $ **FLOATING
C200 a_13599_2388# vssd1 0.52fF $ **FLOATING
C201 a_12299_2589# vssd1 0.61fF $ **FLOATING
C202 a_12467_2491# vssd1 0.82fF $ **FLOATING
C203 a_11874_2589# vssd1 0.63fF $ **FLOATING
C204 a_12042_2335# vssd1 0.58fF $ **FLOATING
C205 a_11601_2223# vssd1 1.43fF $ **FLOATING
C206 a_11435_2223# vssd1 1.81fF $ **FLOATING
C207 a_9949_2223# vssd1 0.23fF $ **FLOATING
C208 a_10459_2589# vssd1 0.61fF $ **FLOATING
C209 a_10627_2491# vssd1 0.82fF $ **FLOATING
C210 a_10034_2589# vssd1 0.63fF $ **FLOATING
C211 a_10202_2335# vssd1 0.58fF $ **FLOATING
C212 a_9761_2223# vssd1 1.43fF $ **FLOATING
C213 a_9595_2223# vssd1 1.81fF $ **FLOATING
C214 a_7465_2223# vssd1 0.23fF $ **FLOATING
C215 a_7975_2589# vssd1 0.61fF $ **FLOATING
C216 a_8143_2491# vssd1 0.82fF $ **FLOATING
C217 a_7550_2589# vssd1 0.63fF $ **FLOATING
C218 a_7718_2335# vssd1 0.58fF $ **FLOATING
C219 a_7277_2223# vssd1 1.43fF $ **FLOATING
C220 _1952_.D vssd1 9.09fF $ **FLOATING
C221 a_7111_2223# vssd1 1.81fF $ **FLOATING
C222 a_5625_2223# vssd1 0.23fF $ **FLOATING
C223 a_6135_2589# vssd1 0.61fF $ **FLOATING
C224 a_6303_2491# vssd1 0.82fF $ **FLOATING
C225 a_5710_2589# vssd1 0.63fF $ **FLOATING
C226 a_5878_2335# vssd1 0.58fF $ **FLOATING
C227 a_5437_2223# vssd1 1.43fF $ **FLOATING
C228 a_5271_2223# vssd1 1.81fF $ **FLOATING
C229 _1650_.X vssd1 10.31fF $ **FLOATING
C230 a_1945_2223# vssd1 0.23fF $ **FLOATING
C231 a_4531_2589# vssd1 0.51fF $ **FLOATING
C232 a_4351_2589# vssd1 0.60fF $ **FLOATING
C233 a_2455_2589# vssd1 0.61fF $ **FLOATING
C234 a_2623_2491# vssd1 0.97fF $ **FLOATING
C235 a_2030_2589# vssd1 0.63fF $ **FLOATING
C236 a_2198_2335# vssd1 0.58fF $ **FLOATING
C237 a_1757_2223# vssd1 1.43fF $ **FLOATING
C238 a_1591_2223# vssd1 1.81fF $ **FLOATING
C239 a_24761_2767# vssd1 0.23fF $ **FLOATING
C240 a_22369_2767# vssd1 0.23fF $ **FLOATING
C241 _1736_.X vssd1 2.90fF $ **FLOATING
C242 a_18597_2767# vssd1 0.23fF $ **FLOATING
C243 _1629_.X vssd1 2.73fF $ **FLOATING
C244 a_14825_2767# vssd1 0.23fF $ **FLOATING
C245 a_12985_2767# vssd1 0.23fF $ **FLOATING
C246 _1612_.X vssd1 1.87fF $ **FLOATING
C247 _1659_.X vssd1 2.55fF $ **FLOATING
C248 a_8569_2767# vssd1 0.23fF $ **FLOATING
C249 _1654_.X vssd1 9.12fF $ **FLOATING
C250 a_5357_3087# vssd1 0.21fF $ **FLOATING
C251 _1808_.Y vssd1 2.94fF $ **FLOATING
C252 a_26295_2986# vssd1 0.52fF $ **FLOATING
C253 a_25271_2767# vssd1 0.61fF $ **FLOATING
C254 a_25439_2741# vssd1 0.82fF $ **FLOATING
C255 a_24846_2767# vssd1 0.63fF $ **FLOATING
C256 a_25014_2741# vssd1 0.58fF $ **FLOATING
C257 a_24573_2773# vssd1 1.43fF $ **FLOATING
C258 _1992_.D vssd1 2.80fF $ **FLOATING
C259 a_24407_2773# vssd1 1.81fF $ **FLOATING
C260 a_22879_2767# vssd1 0.61fF $ **FLOATING
C261 a_23047_2741# vssd1 0.82fF $ **FLOATING
C262 a_22454_2767# vssd1 0.63fF $ **FLOATING
C263 a_22622_2741# vssd1 0.58fF $ **FLOATING
C264 a_22181_2773# vssd1 1.43fF $ **FLOATING
C265 _1993_.D vssd1 2.32fF $ **FLOATING
C266 a_22015_2773# vssd1 1.81fF $ **FLOATING
C267 a_21183_2767# vssd1 0.51fF $ **FLOATING
C268 a_21003_2767# vssd1 0.60fF $ **FLOATING
C269 a_20407_2986# vssd1 0.52fF $ **FLOATING
C270 a_19107_2767# vssd1 0.61fF $ **FLOATING
C271 a_19275_2741# vssd1 0.82fF $ **FLOATING
C272 a_18682_2767# vssd1 0.63fF $ **FLOATING
C273 a_18850_2741# vssd1 0.58fF $ **FLOATING
C274 a_18409_2773# vssd1 1.43fF $ **FLOATING
C275 _1938_.D vssd1 3.10fF $ **FLOATING
C276 a_18243_2773# vssd1 1.81fF $ **FLOATING
C277 a_17180_2883# vssd1 0.50fF $ **FLOATING
C278 a_15335_2767# vssd1 0.61fF $ **FLOATING
C279 a_15503_2741# vssd1 0.82fF $ **FLOATING
C280 a_14910_2767# vssd1 0.63fF $ **FLOATING
C281 a_15078_2741# vssd1 0.58fF $ **FLOATING
C282 a_14637_2773# vssd1 1.43fF $ **FLOATING
C283 _1934_.D vssd1 1.88fF $ **FLOATING
C284 a_14471_2773# vssd1 1.81fF $ **FLOATING
C285 a_13495_2767# vssd1 0.61fF $ **FLOATING
C286 a_13663_2741# vssd1 0.82fF $ **FLOATING
C287 a_13070_2767# vssd1 0.63fF $ **FLOATING
C288 a_13238_2741# vssd1 0.58fF $ **FLOATING
C289 a_12797_2773# vssd1 1.43fF $ **FLOATING
C290 _1955_.D vssd1 3.01fF $ **FLOATING
C291 a_12631_2773# vssd1 1.81fF $ **FLOATING
C292 a_12035_2986# vssd1 0.52fF $ **FLOATING
C293 a_10931_2986# vssd1 0.52fF $ **FLOATING
C294 a_10287_2986# vssd1 0.52fF $ **FLOATING
C295 a_9079_2767# vssd1 0.61fF $ **FLOATING
C296 a_9247_2741# vssd1 0.82fF $ **FLOATING
C297 a_8654_2767# vssd1 0.63fF $ **FLOATING
C298 a_8822_2741# vssd1 0.58fF $ **FLOATING
C299 a_8381_2773# vssd1 1.43fF $ **FLOATING
C300 a_8215_2773# vssd1 1.81fF $ **FLOATING
C301 a_7619_2986# vssd1 0.52fF $ **FLOATING
C302 a_6739_2767# vssd1 0.51fF $ **FLOATING
C303 a_6559_2767# vssd1 0.60fF $ **FLOATING
C304 a_5165_2828# vssd1 0.45fF $ **FLOATING
C305 a_3325_2767# vssd1 0.23fF $ **FLOATING
C306 a_3835_2767# vssd1 0.61fF $ **FLOATING
C307 a_4003_2741# vssd1 0.82fF $ **FLOATING
C308 a_3410_2767# vssd1 0.63fF $ **FLOATING
C309 a_3578_2741# vssd1 0.58fF $ **FLOATING
C310 a_3137_2773# vssd1 1.43fF $ **FLOATING
C311 _1951_.D vssd1 12.04fF $ **FLOATING
C312 a_2971_2773# vssd1 1.81fF $ **FLOATING
C313 a_2235_2775# vssd1 0.65fF $ **FLOATING
C314 a_27337_3311# vssd1 0.23fF $ **FLOATING
C315 a_27847_3677# vssd1 0.61fF $ **FLOATING
C316 a_28015_3579# vssd1 0.82fF $ **FLOATING
C317 a_27422_3677# vssd1 0.63fF $ **FLOATING
C318 a_27590_3423# vssd1 0.58fF $ **FLOATING
C319 a_27149_3311# vssd1 1.43fF $ **FLOATING
C320 a_26983_3311# vssd1 1.81fF $ **FLOATING
C321 a_25497_3311# vssd1 0.23fF $ **FLOATING
C322 a_26007_3677# vssd1 0.61fF $ **FLOATING
C323 a_26175_3579# vssd1 0.82fF $ **FLOATING
C324 a_25582_3677# vssd1 0.63fF $ **FLOATING
C325 a_25750_3423# vssd1 0.58fF $ **FLOATING
C326 a_25309_3311# vssd1 1.43fF $ **FLOATING
C327 _1990_.D vssd1 3.54fF $ **FLOATING
C328 a_25143_3311# vssd1 1.81fF $ **FLOATING
C329 a_23013_3311# vssd1 0.23fF $ **FLOATING
C330 a_23523_3677# vssd1 0.61fF $ **FLOATING
C331 a_23691_3579# vssd1 0.82fF $ **FLOATING
C332 a_23098_3677# vssd1 0.63fF $ **FLOATING
C333 a_23266_3423# vssd1 0.58fF $ **FLOATING
C334 a_22825_3311# vssd1 1.43fF $ **FLOATING
C335 _1989_.D vssd1 2.14fF $ **FLOATING
C336 a_22659_3311# vssd1 1.81fF $ **FLOATING
C337 _1734_.X vssd1 1.60fF $ **FLOATING
C338 _1738_.X vssd1 1.48fF $ **FLOATING
C339 _1740_.X vssd1 1.17fF $ **FLOATING
C340 _1640_.X vssd1 1.83fF $ **FLOATING
C341 a_15929_3311# vssd1 0.23fF $ **FLOATING
C342 a_21459_3677# vssd1 0.51fF $ **FLOATING
C343 a_21279_3677# vssd1 0.60fF $ **FLOATING
C344 a_20539_3677# vssd1 0.51fF $ **FLOATING
C345 a_20359_3677# vssd1 0.60fF $ **FLOATING
C346 a_19619_3677# vssd1 0.51fF $ **FLOATING
C347 a_19439_3677# vssd1 0.60fF $ **FLOATING
C348 a_18383_3476# vssd1 0.52fF $ **FLOATING
C349 a_17595_3677# vssd1 0.51fF $ **FLOATING
C350 a_17415_3677# vssd1 0.60fF $ **FLOATING
C351 a_16439_3677# vssd1 0.61fF $ **FLOATING
C352 a_16607_3579# vssd1 0.82fF $ **FLOATING
C353 a_16014_3677# vssd1 0.63fF $ **FLOATING
C354 a_16182_3423# vssd1 0.58fF $ **FLOATING
C355 a_15741_3311# vssd1 1.43fF $ **FLOATING
C356 a_15575_3311# vssd1 1.81fF $ **FLOATING
C357 _1642_.X vssd1 1.39fF $ **FLOATING
C358 _1625_.X vssd1 1.11fF $ **FLOATING
C359 _1624_.X vssd1 3.33fF $ **FLOATING
C360 a_10777_3311# vssd1 0.23fF $ **FLOATING
C361 a_14328_3561# vssd1 0.50fF $ **FLOATING
C362 a_13408_3561# vssd1 0.50fF $ **FLOATING
C363 a_12771_3476# vssd1 0.52fF $ **FLOATING
C364 a_11287_3677# vssd1 0.61fF $ **FLOATING
C365 a_11455_3579# vssd1 0.82fF $ **FLOATING
C366 a_10862_3677# vssd1 0.63fF $ **FLOATING
C367 a_11030_3423# vssd1 0.58fF $ **FLOATING
C368 a_10589_3311# vssd1 1.43fF $ **FLOATING
C369 a_10423_3311# vssd1 1.81fF $ **FLOATING
C370 a_5541_3311# vssd1 0.21fF $ **FLOATING
C371 a_9135_3311# vssd1 0.70fF $ **FLOATING
C372 a_7704_3561# vssd1 0.50fF $ **FLOATING
C373 a_6223_3339# vssd1 0.56fF $ **FLOATING
C374 a_5349_3616# vssd1 0.45fF $ **FLOATING
C375 a_2129_3311# vssd1 0.23fF $ **FLOATING
C376 a_3983_3311# vssd1 0.70fF $ **FLOATING
C377 a_2639_3677# vssd1 0.61fF $ **FLOATING
C378 a_2807_3579# vssd1 0.97fF $ **FLOATING
C379 a_2214_3677# vssd1 0.63fF $ **FLOATING
C380 a_2382_3423# vssd1 0.58fF $ **FLOATING
C381 a_1941_3311# vssd1 1.43fF $ **FLOATING
C382 a_1775_3311# vssd1 1.81fF $ **FLOATING
C383 _1367_.X vssd1 12.27fF $ **FLOATING
C384 a_25129_3855# vssd1 0.23fF $ **FLOATING
C385 a_23289_3855# vssd1 0.23fF $ **FLOATING
C386 _1732_.X vssd1 1.85fF $ **FLOATING
C387 _1743_.X vssd1 3.32fF $ **FLOATING
C388 a_18597_3855# vssd1 0.23fF $ **FLOATING
C389 _1637_.X vssd1 1.57fF $ **FLOATING
C390 a_14733_3855# vssd1 0.23fF $ **FLOATING
C391 _1660_.X vssd1 3.22fF $ **FLOATING
C392 _1658_.X vssd1 1.11fF $ **FLOATING
C393 _1611_.X vssd1 1.68fF $ **FLOATING
C394 _1567_.X vssd1 1.82fF $ **FLOATING
C395 a_7189_3855# vssd1 0.23fF $ **FLOATING
C396 a_4805_4175# vssd1 0.21fF $ **FLOATING
C397 a_27215_4074# vssd1 0.52fF $ **FLOATING
C398 a_25639_3855# vssd1 0.61fF $ **FLOATING
C399 a_25807_3829# vssd1 0.82fF $ **FLOATING
C400 a_25214_3855# vssd1 0.63fF $ **FLOATING
C401 a_25382_3829# vssd1 0.58fF $ **FLOATING
C402 a_24941_3861# vssd1 1.43fF $ **FLOATING
C403 a_24775_3861# vssd1 1.81fF $ **FLOATING
C404 a_23799_3855# vssd1 0.61fF $ **FLOATING
C405 a_23967_3829# vssd1 0.82fF $ **FLOATING
C406 a_23374_3855# vssd1 0.63fF $ **FLOATING
C407 a_23542_3829# vssd1 0.58fF $ **FLOATING
C408 a_23101_3861# vssd1 1.43fF $ **FLOATING
C409 _1991_.D vssd1 2.23fF $ **FLOATING
C410 a_22935_3861# vssd1 1.81fF $ **FLOATING
C411 a_22195_3855# vssd1 0.51fF $ **FLOATING
C412 a_22015_3855# vssd1 0.60fF $ **FLOATING
C413 _1743_.A vssd1 0.88fF $ **FLOATING
C414 a_21051_4074# vssd1 0.52fF $ **FLOATING
C415 a_20263_3855# vssd1 0.51fF $ **FLOATING
C416 a_20083_3855# vssd1 0.60fF $ **FLOATING
C417 a_19107_3855# vssd1 0.61fF $ **FLOATING
C418 a_19275_3829# vssd1 0.82fF $ **FLOATING
C419 a_18682_3855# vssd1 0.63fF $ **FLOATING
C420 a_18850_3829# vssd1 0.58fF $ **FLOATING
C421 a_18409_3861# vssd1 1.43fF $ **FLOATING
C422 _1935_.D vssd1 3.18fF $ **FLOATING
C423 a_18243_3861# vssd1 1.81fF $ **FLOATING
C424 a_16904_3971# vssd1 0.50fF $ **FLOATING
C425 a_15243_3855# vssd1 0.61fF $ **FLOATING
C426 a_15411_3829# vssd1 0.82fF $ **FLOATING
C427 a_14818_3855# vssd1 0.63fF $ **FLOATING
C428 a_14986_3829# vssd1 0.58fF $ **FLOATING
C429 a_14545_3861# vssd1 1.43fF $ **FLOATING
C430 a_14379_3861# vssd1 1.81fF $ **FLOATING
C431 a_13643_3855# vssd1 0.70fF $ **FLOATING
C432 a_12351_3855# vssd1 0.51fF $ **FLOATING
C433 a_12171_3855# vssd1 0.60fF $ **FLOATING
C434 a_10327_3855# vssd1 0.51fF $ **FLOATING
C435 a_10147_3855# vssd1 0.60fF $ **FLOATING
C436 a_9360_3971# vssd1 0.50fF $ **FLOATING
C437 a_8723_4074# vssd1 0.52fF $ **FLOATING
C438 a_7699_3855# vssd1 0.61fF $ **FLOATING
C439 a_7867_3829# vssd1 0.82fF $ **FLOATING
C440 a_7274_3855# vssd1 0.63fF $ **FLOATING
C441 a_7442_3829# vssd1 0.58fF $ **FLOATING
C442 a_7001_3861# vssd1 1.43fF $ **FLOATING
C443 a_6835_3861# vssd1 1.81fF $ **FLOATING
C444 io_in[5] vssd1 6.17fF
C445 a_5503_4074# vssd1 0.52fF $ **FLOATING
C446 _1800_.A2 vssd1 1.76fF $ **FLOATING
C447 a_4613_3916# vssd1 0.45fF $ **FLOATING
C448 _1652_.X vssd1 12.88fF $ **FLOATING
C449 a_2129_3855# vssd1 0.23fF $ **FLOATING
C450 a_3748_3971# vssd1 0.50fF $ **FLOATING
C451 a_2639_3855# vssd1 0.61fF $ **FLOATING
C452 a_2807_3829# vssd1 0.97fF $ **FLOATING
C453 a_2214_3855# vssd1 0.63fF $ **FLOATING
C454 a_2382_3829# vssd1 0.58fF $ **FLOATING
C455 a_1941_3861# vssd1 1.43fF $ **FLOATING
C456 a_1775_3861# vssd1 1.81fF $ **FLOATING
C457 a_26141_4399# vssd1 0.23fF $ **FLOATING
C458 a_26651_4765# vssd1 0.61fF $ **FLOATING
C459 a_26819_4667# vssd1 0.82fF $ **FLOATING
C460 a_26226_4765# vssd1 0.63fF $ **FLOATING
C461 a_26394_4511# vssd1 0.58fF $ **FLOATING
C462 a_25953_4399# vssd1 1.43fF $ **FLOATING
C463 a_25787_4399# vssd1 1.81fF $ **FLOATING
C464 _1959_.D vssd1 1.34fF $ **FLOATING
C465 a_24025_4399# vssd1 0.23fF $ **FLOATING
C466 a_20529_4399# vssd1 0.23fF $ **FLOATING
C467 _1670_.A vssd1 1.58fF $ **FLOATING
C468 a_24639_4564# vssd1 0.52fF $ **FLOATING
C469 a_23848_4399# vssd1 0.50fF $ **FLOATING
C470 a_23742_4399# vssd1 0.58fF $ **FLOATING
C471 a_23565_4399# vssd1 0.50fF $ **FLOATING
C472 fanout21.X vssd1 6.78fF $ **FLOATING
C473 a_23246_4399# vssd1 0.54fF $ **FLOATING
C474 a_22195_4765# vssd1 0.51fF $ **FLOATING
C475 a_22015_4765# vssd1 0.60fF $ **FLOATING
C476 a_21039_4765# vssd1 0.61fF $ **FLOATING
C477 a_21207_4667# vssd1 0.82fF $ **FLOATING
C478 a_20614_4765# vssd1 0.63fF $ **FLOATING
C479 a_20782_4511# vssd1 0.58fF $ **FLOATING
C480 a_20341_4399# vssd1 1.43fF $ **FLOATING
C481 _1941_.D vssd1 2.01fF $ **FLOATING
C482 a_20175_4399# vssd1 1.81fF $ **FLOATING
C483 _1941_.CLK vssd1 13.15fF $ **FLOATING
C484 _1636_.X vssd1 3.10fF $ **FLOATING
C485 _1631_.X vssd1 1.49fF $ **FLOATING
C486 a_16573_4399# vssd1 0.23fF $ **FLOATING
C487 _1622_.X vssd1 1.12fF $ **FLOATING
C488 _1619_.X vssd1 1.62fF $ **FLOATING
C489 _1623_.X vssd1 1.16fF $ **FLOATING
C490 _1617_.X vssd1 1.32fF $ **FLOATING
C491 a_9489_4399# vssd1 0.23fF $ **FLOATING
C492 _1636_.A vssd1 1.11fF $ **FLOATING
C493 a_19487_4564# vssd1 0.52fF $ **FLOATING
C494 a_18147_4765# vssd1 0.51fF $ **FLOATING
C495 a_17967_4765# vssd1 0.60fF $ **FLOATING
C496 a_17227_4765# vssd1 0.51fF $ **FLOATING
C497 a_17047_4765# vssd1 0.60fF $ **FLOATING
C498 a_16396_4399# vssd1 0.50fF $ **FLOATING
C499 a_16290_4399# vssd1 0.58fF $ **FLOATING
C500 a_16113_4399# vssd1 0.50fF $ **FLOATING
C501 a_15794_4399# vssd1 0.54fF $ **FLOATING
C502 a_15163_4564# vssd1 0.52fF $ **FLOATING
C503 a_14328_4649# vssd1 0.50fF $ **FLOATING
C504 a_13455_4765# vssd1 0.51fF $ **FLOATING
C505 a_13275_4765# vssd1 0.60fF $ **FLOATING
C506 a_12488_4649# vssd1 0.50fF $ **FLOATING
C507 a_11707_4765# vssd1 0.51fF $ **FLOATING
C508 a_11527_4765# vssd1 0.60fF $ **FLOATING
C509 a_9999_4765# vssd1 0.61fF $ **FLOATING
C510 a_10167_4667# vssd1 0.82fF $ **FLOATING
C511 a_9574_4765# vssd1 0.63fF $ **FLOATING
C512 a_9742_4511# vssd1 0.58fF $ **FLOATING
C513 a_9301_4399# vssd1 1.43fF $ **FLOATING
C514 a_9135_4399# vssd1 1.81fF $ **FLOATING
C515 a_7373_4399# vssd1 0.23fF $ **FLOATING
C516 a_7883_4765# vssd1 0.61fF $ **FLOATING
C517 a_8051_4667# vssd1 0.82fF $ **FLOATING
C518 a_7458_4765# vssd1 0.63fF $ **FLOATING
C519 a_7626_4511# vssd1 0.58fF $ **FLOATING
C520 a_7185_4399# vssd1 1.43fF $ **FLOATING
C521 _1816_.D vssd1 2.38fF $ **FLOATING
C522 a_7019_4399# vssd1 1.81fF $ **FLOATING
C523 _1816_.CLK vssd1 10.56fF $ **FLOATING
C524 _1999_.CLK vssd1 12.08fF $ **FLOATING
C525 a_2129_4399# vssd1 0.23fF $ **FLOATING
C526 a_6283_4399# vssd1 0.70fF $ **FLOATING
C527 a_5687_4564# vssd1 0.52fF $ **FLOATING
C528 a_4116_4649# vssd1 0.50fF $ **FLOATING
C529 a_2639_4765# vssd1 0.61fF $ **FLOATING
C530 a_2807_4667# vssd1 0.97fF $ **FLOATING
C531 a_2214_4765# vssd1 0.63fF $ **FLOATING
C532 a_2382_4511# vssd1 0.58fF $ **FLOATING
C533 a_1941_4399# vssd1 1.43fF $ **FLOATING
C534 a_1775_4399# vssd1 1.81fF $ **FLOATING
C535 a_25589_4943# vssd1 0.23fF $ **FLOATING
C536 _1731_.X vssd1 3.00fF $ **FLOATING
C537 a_23013_4943# vssd1 0.23fF $ **FLOATING
C538 a_17730_4943# vssd1 0.33fF $ **FLOATING
C539 _1668_.X vssd1 4.76fF $ **FLOATING
C540 a_14733_4943# vssd1 0.23fF $ **FLOATING
C541 _1610_.X vssd1 2.28fF $ **FLOATING
C542 a_10094_4943# vssd1 0.33fF $ **FLOATING
C543 a_12249_4943# vssd1 0.23fF $ **FLOATING
C544 _1647_.X vssd1 2.12fF $ **FLOATING
C545 _1566_.X vssd1 1.02fF $ **FLOATING
C546 a_7002_4943# vssd1 0.51fF $ **FLOATING
C547 a_6559_4943# vssd1 0.32fF $ **FLOATING
C548 a_7002_5263# vssd1 0.28fF $ **FLOATING
C549 _1318_.X vssd1 10.49fF $ **FLOATING
C550 a_4163_4943# vssd1 0.25fF $ **FLOATING
C551 _1365_.X vssd1 2.12fF $ **FLOATING
C552 a_2129_4943# vssd1 0.23fF $ **FLOATING
C553 a_26099_4943# vssd1 0.61fF $ **FLOATING
C554 a_26267_4917# vssd1 0.82fF $ **FLOATING
C555 a_25674_4943# vssd1 0.63fF $ **FLOATING
C556 a_25842_4917# vssd1 0.58fF $ **FLOATING
C557 a_25401_4949# vssd1 1.43fF $ **FLOATING
C558 _1960_.D vssd1 2.20fF $ **FLOATING
C559 a_25235_4949# vssd1 1.81fF $ **FLOATING
C560 a_24547_5162# vssd1 0.52fF $ **FLOATING
C561 a_23523_4943# vssd1 0.61fF $ **FLOATING
C562 a_23691_4917# vssd1 0.82fF $ **FLOATING
C563 a_23098_4943# vssd1 0.63fF $ **FLOATING
C564 a_23266_4917# vssd1 0.58fF $ **FLOATING
C565 a_22825_4949# vssd1 1.43fF $ **FLOATING
C566 _1929_.D vssd1 1.96fF $ **FLOATING
C567 a_22659_4949# vssd1 1.81fF $ **FLOATING
C568 _1672_.A vssd1 1.00fF $ **FLOATING
C569 a_22063_5162# vssd1 0.52fF $ **FLOATING
C570 a_20999_4943# vssd1 0.51fF $ **FLOATING
C571 a_20819_4943# vssd1 0.60fF $ **FLOATING
C572 a_20039_5162# vssd1 0.52fF $ **FLOATING
C573 a_19395_5162# vssd1 0.52fF $ **FLOATING
C574 a_18751_5162# vssd1 0.52fF $ **FLOATING
C575 _1150_.B2 vssd1 4.37fF $ **FLOATING
C576 _1150_.A2 vssd1 6.31fF $ **FLOATING
C577 a_17573_4917# vssd1 0.72fF $ **FLOATING
C578 a_16911_5162# vssd1 0.52fF $ **FLOATING
C579 a_15243_4943# vssd1 0.61fF $ **FLOATING
C580 a_15411_4917# vssd1 0.82fF $ **FLOATING
C581 a_14818_4943# vssd1 0.63fF $ **FLOATING
C582 a_14986_4917# vssd1 0.58fF $ **FLOATING
C583 a_14545_4949# vssd1 1.43fF $ **FLOATING
C584 a_14379_4949# vssd1 1.81fF $ **FLOATING
C585 a_13783_5162# vssd1 0.52fF $ **FLOATING
C586 a_12759_4943# vssd1 0.61fF $ **FLOATING
C587 a_12927_4917# vssd1 0.82fF $ **FLOATING
C588 a_12334_4943# vssd1 0.63fF $ **FLOATING
C589 a_12502_4917# vssd1 0.58fF $ **FLOATING
C590 a_12061_4949# vssd1 1.43fF $ **FLOATING
C591 a_11895_4949# vssd1 1.81fF $ **FLOATING
C592 _1646_.X vssd1 1.94fF $ **FLOATING
C593 a_11023_5162# vssd1 0.52fF $ **FLOATING
C594 _0989_.B2 vssd1 3.04fF $ **FLOATING
C595 _0989_.A2 vssd1 5.09fF $ **FLOATING
C596 a_9937_4917# vssd1 0.72fF $ **FLOATING
C597 a_8579_4943# vssd1 0.51fF $ **FLOATING
C598 a_8399_4943# vssd1 0.60fF $ **FLOATING
C599 a_6644_5263# vssd1 1.17fF $ **FLOATING
C600 _1202_.Y vssd1 10.72fF $ **FLOATING
C601 a_5487_5281# vssd1 0.56fF $ **FLOATING
C602 a_4859_5162# vssd1 0.52fF $ **FLOATING
C603 _1802_.X vssd1 0.90fF $ **FLOATING
C604 a_3945_4917# vssd1 0.55fF $ **FLOATING
C605 a_2639_4943# vssd1 0.61fF $ **FLOATING
C606 a_2807_4917# vssd1 0.82fF $ **FLOATING
C607 a_2214_4943# vssd1 0.63fF $ **FLOATING
C608 a_2382_4917# vssd1 0.58fF $ **FLOATING
C609 a_1941_4949# vssd1 1.43fF $ **FLOATING
C610 _2021_.D vssd1 3.03fF $ **FLOATING
C611 a_1775_4949# vssd1 1.81fF $ **FLOATING
C612 a_27337_5487# vssd1 0.23fF $ **FLOATING
C613 a_27847_5853# vssd1 0.61fF $ **FLOATING
C614 a_28015_5755# vssd1 0.82fF $ **FLOATING
C615 a_27422_5853# vssd1 0.63fF $ **FLOATING
C616 a_27590_5599# vssd1 0.58fF $ **FLOATING
C617 a_27149_5487# vssd1 1.43fF $ **FLOATING
C618 a_26983_5487# vssd1 1.81fF $ **FLOATING
C619 a_24945_5487# vssd1 0.23fF $ **FLOATING
C620 a_25455_5853# vssd1 0.61fF $ **FLOATING
C621 a_25623_5755# vssd1 0.82fF $ **FLOATING
C622 a_25030_5853# vssd1 0.63fF $ **FLOATING
C623 a_25198_5599# vssd1 0.58fF $ **FLOATING
C624 a_24757_5487# vssd1 1.43fF $ **FLOATING
C625 a_24591_5487# vssd1 1.81fF $ **FLOATING
C626 _1730_.X vssd1 1.09fF $ **FLOATING
C627 a_22093_5487# vssd1 0.23fF $ **FLOATING
C628 a_23759_5853# vssd1 0.51fF $ **FLOATING
C629 a_23579_5853# vssd1 0.60fF $ **FLOATING
C630 a_22603_5853# vssd1 0.61fF $ **FLOATING
C631 a_22771_5755# vssd1 0.82fF $ **FLOATING
C632 a_22178_5853# vssd1 0.63fF $ **FLOATING
C633 a_22346_5599# vssd1 0.58fF $ **FLOATING
C634 a_21905_5487# vssd1 1.43fF $ **FLOATING
C635 _1923_.D vssd1 2.31fF $ **FLOATING
C636 a_21739_5487# vssd1 1.81fF $ **FLOATING
C637 a_19793_5487# vssd1 0.23fF $ **FLOATING
C638 a_20303_5853# vssd1 0.61fF $ **FLOATING
C639 a_20471_5755# vssd1 0.82fF $ **FLOATING
C640 a_19878_5853# vssd1 0.63fF $ **FLOATING
C641 a_20046_5599# vssd1 0.58fF $ **FLOATING
C642 a_19605_5487# vssd1 1.43fF $ **FLOATING
C643 _1942_.D vssd1 2.17fF $ **FLOATING
C644 a_19439_5487# vssd1 1.81fF $ **FLOATING
C645 _1607_.X vssd1 1.47fF $ **FLOATING
C646 _1607_.B vssd1 12.74fF $ **FLOATING
C647 _1633_.X vssd1 1.05fF $ **FLOATING
C648 a_16074_5737# vssd1 0.33fF $ **FLOATING
C649 _1066_.B vssd1 7.57fF $ **FLOATING
C650 a_13130_5737# vssd1 0.33fF $ **FLOATING
C651 _1067_.B vssd1 4.78fF $ **FLOATING
C652 _1356_.X vssd1 4.64fF $ **FLOATING
C653 a_9489_5487# vssd1 0.23fF $ **FLOATING
C654 a_18468_5737# vssd1 0.50fF $ **FLOATING
C655 a_17319_5853# vssd1 0.51fF $ **FLOATING
C656 a_17139_5853# vssd1 0.60fF $ **FLOATING
C657 _1195_.B2 vssd1 5.51fF $ **FLOATING
C658 _1195_.A2 vssd1 5.67fF $ **FLOATING
C659 a_15917_5461# vssd1 0.72fF $ **FLOATING
C660 a_15115_5487# vssd1 0.70fF $ **FLOATING
C661 a_14287_5487# vssd1 0.62fF $ **FLOATING
C662 _1194_.B2 vssd1 3.32fF $ **FLOATING
C663 _1194_.A2 vssd1 4.88fF $ **FLOATING
C664 a_12973_5461# vssd1 0.72fF $ **FLOATING
C665 a_11711_5487# vssd1 0.62fF $ **FLOATING
C666 a_11023_5652# vssd1 0.52fF $ **FLOATING
C667 a_9999_5853# vssd1 0.61fF $ **FLOATING
C668 a_10167_5755# vssd1 0.82fF $ **FLOATING
C669 a_9574_5853# vssd1 0.63fF $ **FLOATING
C670 a_9742_5599# vssd1 0.58fF $ **FLOATING
C671 a_9301_5487# vssd1 1.43fF $ **FLOATING
C672 _2001_.D vssd1 2.72fF $ **FLOATING
C673 a_9135_5487# vssd1 1.81fF $ **FLOATING
C674 _1565_.X vssd1 2.41fF $ **FLOATING
C675 a_5817_5487# vssd1 0.21fF $ **FLOATING
C676 _1798_.Y vssd1 3.20fF $ **FLOATING
C677 a_8307_5487# vssd1 0.70fF $ **FLOATING
C678 a_7711_5652# vssd1 0.52fF $ **FLOATING
C679 a_6831_5853# vssd1 0.51fF $ **FLOATING
C680 a_6651_5853# vssd1 0.60fF $ **FLOATING
C681 a_5625_5792# vssd1 0.45fF $ **FLOATING
C682 _1366_.X vssd1 11.04fF $ **FLOATING
C683 a_4069_5737# vssd1 0.24fF $ **FLOATING
C684 _1804_.Y vssd1 2.23fF $ **FLOATING
C685 a_4760_5737# vssd1 0.50fF $ **FLOATING
C686 io_in[6] vssd1 5.10fF
C687 a_3111_5652# vssd1 0.52fF $ **FLOATING
C688 a_2327_5487# vssd1 0.70fF $ **FLOATING
C689 io_in[1] vssd1 2.36fF
C690 a_1591_5487# vssd1 0.70fF $ **FLOATING
C691 io_in[2] vssd1 1.25fF
C692 a_25589_6031# vssd1 0.23fF $ **FLOATING
C693 _1674_.X vssd1 3.18fF $ **FLOATING
C694 fanout20.X vssd1 11.25fF $ **FLOATING
C695 a_22829_6031# vssd1 0.23fF $ **FLOATING
C696 a_17270_6031# vssd1 0.33fF $ **FLOATING
C697 a_15614_6031# vssd1 0.33fF $ **FLOATING
C698 _1745_.X vssd1 3.84fF $ **FLOATING
C699 _1807_.Y vssd1 8.31fF $ **FLOATING
C700 _1621_.X vssd1 1.99fF $ **FLOATING
C701 a_11877_6031# vssd1 0.21fF $ **FLOATING
C702 a_11793_6031# vssd1 0.17fF $ **FLOATING
C703 _1639_.X vssd1 15.10fF $ **FLOATING
C704 a_10133_6031# vssd1 0.23fF $ **FLOATING
C705 a_7742_6031# vssd1 0.32fF $ **FLOATING
C706 a_7828_6351# vssd1 0.34fF $ **FLOATING
C707 a_7295_6351# vssd1 0.28fF $ **FLOATING
C708 _1783_.X vssd1 3.32fF $ **FLOATING
C709 a_2129_6031# vssd1 0.23fF $ **FLOATING
C710 a_26099_6031# vssd1 0.61fF $ **FLOATING
C711 a_26267_6005# vssd1 0.82fF $ **FLOATING
C712 a_25674_6031# vssd1 0.63fF $ **FLOATING
C713 a_25842_6005# vssd1 0.58fF $ **FLOATING
C714 a_25401_6037# vssd1 1.43fF $ **FLOATING
C715 a_25235_6037# vssd1 1.81fF $ **FLOATING
C716 _1674_.A vssd1 2.02fF $ **FLOATING
C717 a_24087_6250# vssd1 0.52fF $ **FLOATING
C718 a_23303_6031# vssd1 0.70fF $ **FLOATING
C719 a_22652_6031# vssd1 0.50fF $ **FLOATING
C720 a_22546_6031# vssd1 0.58fF $ **FLOATING
C721 a_22369_6031# vssd1 0.50fF $ **FLOATING
C722 a_22050_6031# vssd1 0.54fF $ **FLOATING
C723 a_20907_6031# vssd1 0.51fF $ **FLOATING
C724 a_20727_6031# vssd1 0.60fF $ **FLOATING
C725 a_20131_6250# vssd1 0.52fF $ **FLOATING
C726 a_18151_6031# vssd1 0.70fF $ **FLOATING
C727 _0998_.B2 vssd1 6.01fF $ **FLOATING
C728 _0998_.A2 vssd1 4.86fF $ **FLOATING
C729 a_17113_6005# vssd1 0.72fF $ **FLOATING
C730 _0994_.B2 vssd1 5.72fF $ **FLOATING
C731 _0994_.A2 vssd1 5.28fF $ **FLOATING
C732 a_15457_6005# vssd1 0.72fF $ **FLOATING
C733 a_14283_6031# vssd1 0.51fF $ **FLOATING
C734 a_14103_6031# vssd1 0.60fF $ **FLOATING
C735 a_12815_6031# vssd1 0.70fF $ **FLOATING
C736 a_11711_6031# vssd1 0.97fF $ **FLOATING
C737 _1145_.A1 vssd1 4.45fF $ **FLOATING
C738 _1145_.B2 vssd1 3.10fF $ **FLOATING
C739 a_10643_6031# vssd1 0.61fF $ **FLOATING
C740 a_10811_6005# vssd1 0.82fF $ **FLOATING
C741 a_10218_6031# vssd1 0.63fF $ **FLOATING
C742 a_10386_6005# vssd1 0.58fF $ **FLOATING
C743 a_9945_6037# vssd1 1.43fF $ **FLOATING
C744 a_9779_6037# vssd1 1.81fF $ **FLOATING
C745 a_8859_6144# vssd1 0.62fF $ **FLOATING
C746 _1188_.B vssd1 5.14fF $ **FLOATING
C747 a_7295_6031# vssd1 1.14fF $ **FLOATING
C748 a_6607_6250# vssd1 0.52fF $ **FLOATING
C749 a_4627_6031# vssd1 0.70fF $ **FLOATING
C750 a_3707_6144# vssd1 0.62fF $ **FLOATING
C751 a_2639_6031# vssd1 0.61fF $ **FLOATING
C752 a_2807_6005# vssd1 0.97fF $ **FLOATING
C753 a_2214_6031# vssd1 0.63fF $ **FLOATING
C754 a_2382_6005# vssd1 0.58fF $ **FLOATING
C755 a_1941_6037# vssd1 1.43fF $ **FLOATING
C756 _2019_.D vssd1 2.92fF $ **FLOATING
C757 a_1775_6037# vssd1 1.81fF $ **FLOATING
C758 a_26785_6575# vssd1 0.23fF $ **FLOATING
C759 a_27295_6941# vssd1 0.61fF $ **FLOATING
C760 a_27463_6843# vssd1 0.82fF $ **FLOATING
C761 a_26870_6941# vssd1 0.63fF $ **FLOATING
C762 a_27038_6687# vssd1 0.58fF $ **FLOATING
C763 a_26597_6575# vssd1 1.43fF $ **FLOATING
C764 a_26431_6575# vssd1 1.81fF $ **FLOATING
C765 a_24945_6575# vssd1 0.23fF $ **FLOATING
C766 a_25455_6941# vssd1 0.61fF $ **FLOATING
C767 a_25623_6843# vssd1 0.82fF $ **FLOATING
C768 a_25030_6941# vssd1 0.63fF $ **FLOATING
C769 a_25198_6687# vssd1 0.58fF $ **FLOATING
C770 a_24757_6575# vssd1 1.43fF $ **FLOATING
C771 a_24591_6575# vssd1 1.81fF $ **FLOATING
C772 _1593_.X vssd1 1.76fF $ **FLOATING
C773 a_22093_6575# vssd1 0.23fF $ **FLOATING
C774 a_23627_6740# vssd1 0.52fF $ **FLOATING
C775 a_22603_6941# vssd1 0.61fF $ **FLOATING
C776 a_22771_6843# vssd1 0.82fF $ **FLOATING
C777 a_22178_6941# vssd1 0.63fF $ **FLOATING
C778 a_22346_6687# vssd1 0.58fF $ **FLOATING
C779 a_21905_6575# vssd1 1.43fF $ **FLOATING
C780 a_21739_6575# vssd1 1.81fF $ **FLOATING
C781 _1667_.X vssd1 1.67fF $ **FLOATING
C782 _1609_.X vssd1 2.38fF $ **FLOATING
C783 _1065_.B vssd1 8.58fF $ **FLOATING
C784 _1063_.B vssd1 6.17fF $ **FLOATING
C785 a_13120_6825# vssd1 0.26fF $ **FLOATING
C786 _1117_.B vssd1 3.82fF $ **FLOATING
C787 a_10681_6825# vssd1 0.21fF $ **FLOATING
C788 a_10597_6825# vssd1 0.17fF $ **FLOATING
C789 _1144_.X vssd1 1.47fF $ **FLOATING
C790 _1144_.B vssd1 5.38fF $ **FLOATING
C791 _1753_.X vssd1 2.32fF $ **FLOATING
C792 _1756_.X vssd1 1.91fF $ **FLOATING
C793 _1368_.X vssd1 2.62fF $ **FLOATING
C794 a_4341_6621# vssd1 0.43fF $ **FLOATING
C795 a_1945_6575# vssd1 0.23fF $ **FLOATING
C796 a_20539_6941# vssd1 0.51fF $ **FLOATING
C797 a_20359_6941# vssd1 0.60fF $ **FLOATING
C798 a_19619_6941# vssd1 0.51fF $ **FLOATING
C799 a_19439_6941# vssd1 0.60fF $ **FLOATING
C800 a_18239_6941# vssd1 0.51fF $ **FLOATING
C801 a_18059_6941# vssd1 0.60fF $ **FLOATING
C802 a_17319_6941# vssd1 0.51fF $ **FLOATING
C803 a_17139_6941# vssd1 0.60fF $ **FLOATING
C804 a_16307_6941# vssd1 0.51fF $ **FLOATING
C805 a_16127_6941# vssd1 0.60fF $ **FLOATING
C806 a_15299_6575# vssd1 0.62fF $ **FLOATING
C807 a_14471_6575# vssd1 0.62fF $ **FLOATING
C808 _1068_.A1 vssd1 3.58fF $ **FLOATING
C809 _1065_.X vssd1 1.75fF $ **FLOATING
C810 _1068_.C1 vssd1 1.80fF $ **FLOATING
C811 _1068_.D1 vssd1 1.43fF $ **FLOATING
C812 a_12689_6721# vssd1 0.67fF $ **FLOATING
C813 a_11803_6575# vssd1 0.62fF $ **FLOATING
C814 a_10515_6575# vssd1 0.97fF $ **FLOATING
C815 _1189_.B2 vssd1 4.17fF $ **FLOATING
C816 _1189_.C1 vssd1 1.31fF $ **FLOATING
C817 a_9687_6575# vssd1 0.62fF $ **FLOATING
C818 a_8447_6740# vssd1 0.52fF $ **FLOATING
C819 a_7803_6740# vssd1 0.52fF $ **FLOATING
C820 a_6555_6941# vssd1 0.51fF $ **FLOATING
C821 a_6375_6941# vssd1 0.60fF $ **FLOATING
C822 a_5588_6825# vssd1 0.50fF $ **FLOATING
C823 a_4447_6581# vssd1 0.67fF $ **FLOATING
C824 a_2455_6941# vssd1 0.61fF $ **FLOATING
C825 a_2623_6843# vssd1 0.82fF $ **FLOATING
C826 a_2030_6941# vssd1 0.63fF $ **FLOATING
C827 a_2198_6687# vssd1 0.58fF $ **FLOATING
C828 a_1757_6575# vssd1 1.43fF $ **FLOATING
C829 a_1591_6575# vssd1 1.81fF $ **FLOATING
C830 a_24945_7119# vssd1 0.23fF $ **FLOATING
C831 _1676_.X vssd1 2.42fF $ **FLOATING
C832 _1744_.X vssd1 1.11fF $ **FLOATING
C833 a_17812_7119# vssd1 0.26fF $ **FLOATING
C834 a_14549_7119# vssd1 0.23fF $ **FLOATING
C835 _1657_.X vssd1 3.53fF $ **FLOATING
C836 _1649_.X vssd1 5.91fF $ **FLOATING
C837 a_9489_7119# vssd1 0.23fF $ **FLOATING
C838 _1359_.X vssd1 0.88fF $ **FLOATING
C839 _1171_.Y vssd1 1.65fF $ **FLOATING
C840 a_6835_7439# vssd1 0.18fF $ **FLOATING
C841 a_4061_7119# vssd1 0.23fF $ **FLOATING
C842 a_2129_7119# vssd1 0.23fF $ **FLOATING
C843 a_25455_7119# vssd1 0.61fF $ **FLOATING
C844 a_25623_7093# vssd1 0.82fF $ **FLOATING
C845 a_25030_7119# vssd1 0.63fF $ **FLOATING
C846 a_25198_7093# vssd1 0.58fF $ **FLOATING
C847 a_24757_7125# vssd1 1.43fF $ **FLOATING
C848 a_24591_7125# vssd1 1.81fF $ **FLOATING
C849 a_23443_7338# vssd1 0.52fF $ **FLOATING
C850 a_22799_7338# vssd1 0.52fF $ **FLOATING
C851 a_22015_7119# vssd1 0.70fF $ **FLOATING
C852 _1597_.A vssd1 1.58fF $ **FLOATING
C853 a_21235_7338# vssd1 0.52fF $ **FLOATING
C854 _1747_.A vssd1 0.88fF $ **FLOATING
C855 a_20591_7338# vssd1 0.52fF $ **FLOATING
C856 a_19803_7119# vssd1 0.51fF $ **FLOATING
C857 a_19623_7119# vssd1 0.60fF $ **FLOATING
C858 _1744_.A_N vssd1 11.28fF $ **FLOATING
C859 a_18795_7232# vssd1 0.62fF $ **FLOATING
C860 _1061_.B vssd1 7.10fF $ **FLOATING
C861 _1744_.B vssd1 6.72fF $ **FLOATING
C862 _1061_.X vssd1 1.21fF $ **FLOATING
C863 _1064_.D1 vssd1 2.12fF $ **FLOATING
C864 a_17381_7093# vssd1 0.67fF $ **FLOATING
C865 a_16035_7119# vssd1 0.70fF $ **FLOATING
C866 a_15059_7119# vssd1 0.61fF $ **FLOATING
C867 a_15227_7093# vssd1 0.82fF $ **FLOATING
C868 a_14634_7119# vssd1 0.63fF $ **FLOATING
C869 a_14802_7093# vssd1 0.58fF $ **FLOATING
C870 a_14361_7125# vssd1 1.43fF $ **FLOATING
C871 a_14195_7125# vssd1 1.81fF $ **FLOATING
C872 a_12907_7232# vssd1 0.62fF $ **FLOATING
C873 _1039_.B vssd1 5.25fF $ **FLOATING
C874 _1657_.A vssd1 5.08fF $ **FLOATING
C875 a_11759_7338# vssd1 0.52fF $ **FLOATING
C876 _1649_.A vssd1 4.22fF $ **FLOATING
C877 a_11023_7338# vssd1 0.52fF $ **FLOATING
C878 a_9999_7119# vssd1 0.61fF $ **FLOATING
C879 a_10167_7093# vssd1 0.82fF $ **FLOATING
C880 a_9574_7119# vssd1 0.63fF $ **FLOATING
C881 a_9742_7093# vssd1 0.58fF $ **FLOATING
C882 a_9301_7125# vssd1 1.43fF $ **FLOATING
C883 _1812_.D vssd1 1.39fF $ **FLOATING
C884 a_9135_7125# vssd1 1.81fF $ **FLOATING
C885 a_8395_7119# vssd1 0.51fF $ **FLOATING
C886 a_8215_7119# vssd1 0.60fF $ **FLOATING
C887 a_5731_7127# vssd1 0.65fF $ **FLOATING
C888 a_4571_7119# vssd1 0.61fF $ **FLOATING
C889 a_4739_7093# vssd1 0.82fF $ **FLOATING
C890 a_4146_7119# vssd1 0.63fF $ **FLOATING
C891 a_4314_7093# vssd1 0.58fF $ **FLOATING
C892 a_3873_7125# vssd1 1.43fF $ **FLOATING
C893 _2020_.D vssd1 1.64fF $ **FLOATING
C894 a_3707_7125# vssd1 1.81fF $ **FLOATING
C895 a_2639_7119# vssd1 0.61fF $ **FLOATING
C896 a_2807_7093# vssd1 0.97fF $ **FLOATING
C897 a_2214_7119# vssd1 0.63fF $ **FLOATING
C898 a_2382_7093# vssd1 0.58fF $ **FLOATING
C899 a_1941_7125# vssd1 1.43fF $ **FLOATING
C900 a_1775_7125# vssd1 1.81fF $ **FLOATING
C901 a_26141_7663# vssd1 0.23fF $ **FLOATING
C902 a_26651_8029# vssd1 0.61fF $ **FLOATING
C903 a_26819_7931# vssd1 0.82fF $ **FLOATING
C904 a_26226_8029# vssd1 0.63fF $ **FLOATING
C905 a_26394_7775# vssd1 0.58fF $ **FLOATING
C906 a_25953_7663# vssd1 1.43fF $ **FLOATING
C907 a_25787_7663# vssd1 1.81fF $ **FLOATING
C908 _1982_.CLK vssd1 7.70fF $ **FLOATING
C909 _1982_.D vssd1 1.34fF $ **FLOATING
C910 _1675_.X vssd1 1.14fF $ **FLOATING
C911 a_20897_7663# vssd1 0.23fF $ **FLOATING
C912 a_24639_7828# vssd1 0.52fF $ **FLOATING
C913 a_23351_7828# vssd1 0.52fF $ **FLOATING
C914 a_22563_8029# vssd1 0.51fF $ **FLOATING
C915 a_22383_8029# vssd1 0.60fF $ **FLOATING
C916 a_21407_8029# vssd1 0.61fF $ **FLOATING
C917 a_21575_7931# vssd1 0.82fF $ **FLOATING
C918 a_20982_8029# vssd1 0.63fF $ **FLOATING
C919 a_21150_7775# vssd1 0.58fF $ **FLOATING
C920 a_20709_7663# vssd1 1.43fF $ **FLOATING
C921 _1996_.D vssd1 1.02fF $ **FLOATING
C922 a_20543_7663# vssd1 1.81fF $ **FLOATING
C923 _1111_.B vssd1 4.79fF $ **FLOATING
C924 _1592_.X vssd1 3.38fF $ **FLOATING
C925 _1594_.X vssd1 2.20fF $ **FLOATING
C926 a_16156_7913# vssd1 0.26fF $ **FLOATING
C927 _0988_.X vssd1 4.93fF $ **FLOATING
C928 _1749_.X vssd1 2.21fF $ **FLOATING
C929 _1148_.B vssd1 4.86fF $ **FLOATING
C930 _1614_.X vssd1 4.02fF $ **FLOATING
C931 _1751_.X vssd1 3.41fF $ **FLOATING
C932 _1752_.X vssd1 1.22fF $ **FLOATING
C933 _1809_.B vssd1 3.35fF $ **FLOATING
C934 _1173_.X vssd1 2.52fF $ **FLOATING
C935 a_5629_7913# vssd1 0.21fF $ **FLOATING
C936 a_4715_7913# vssd1 0.25fF $ **FLOATING
C937 a_2037_7663# vssd1 0.23fF $ **FLOATING
C938 a_19439_7663# vssd1 0.62fF $ **FLOATING
C939 a_18560_7913# vssd1 0.50fF $ **FLOATING
C940 a_17456_7913# vssd1 0.50fF $ **FLOATING
C941 _1041_.A1 vssd1 7.09fF $ **FLOATING
C942 _1041_.C1 vssd1 2.03fF $ **FLOATING
C943 a_15725_7809# vssd1 0.67fF $ **FLOATING
C944 a_14319_7691# vssd1 0.56fF $ **FLOATING
C945 _1749_.A vssd1 2.74fF $ **FLOATING
C946 a_13599_7828# vssd1 0.52fF $ **FLOATING
C947 a_12539_7663# vssd1 0.70fF $ **FLOATING
C948 a_11711_7663# vssd1 0.62fF $ **FLOATING
C949 _1614_.A vssd1 3.49fF $ **FLOATING
C950 a_11115_7828# vssd1 0.52fF $ **FLOATING
C951 a_10471_7828# vssd1 0.52fF $ **FLOATING
C952 a_9683_8029# vssd1 0.51fF $ **FLOATING
C953 a_9503_8029# vssd1 0.60fF $ **FLOATING
C954 _1750_.X vssd1 1.19fF $ **FLOATING
C955 a_8447_7828# vssd1 0.52fF $ **FLOATING
C956 a_7659_8029# vssd1 0.51fF $ **FLOATING
C957 a_7479_8029# vssd1 0.60fF $ **FLOATING
C958 a_6600_7913# vssd1 0.50fF $ **FLOATING
C959 a_5547_7913# vssd1 0.80fF $ **FLOATING
C960 a_4497_7637# vssd1 0.55fF $ **FLOATING
C961 a_2547_8029# vssd1 0.61fF $ **FLOATING
C962 a_2715_7931# vssd1 0.97fF $ **FLOATING
C963 a_2122_8029# vssd1 0.63fF $ **FLOATING
C964 a_2290_7775# vssd1 0.58fF $ **FLOATING
C965 a_1849_7663# vssd1 1.43fF $ **FLOATING
C966 a_1683_7663# vssd1 1.81fF $ **FLOATING
C967 a_25313_8207# vssd1 0.23fF $ **FLOATING
C968 a_23473_8207# vssd1 0.23fF $ **FLOATING
C969 _1599_.X vssd1 2.86fF $ **FLOATING
C970 _1582_.X vssd1 2.19fF $ **FLOATING
C971 _1040_.X vssd1 1.71fF $ **FLOATING
C972 a_14453_8207# vssd1 0.21fF $ **FLOATING
C973 a_14369_8207# vssd1 0.17fF $ **FLOATING
C974 a_12065_8207# vssd1 0.23fF $ **FLOATING
C975 a_10133_8207# vssd1 0.23fF $ **FLOATING
C976 _1364_.X vssd1 3.77fF $ **FLOATING
C977 _1564_.X vssd1 2.10fF $ **FLOATING
C978 _1168_.X vssd1 2.47fF $ **FLOATING
C979 _1355_.X vssd1 4.35fF $ **FLOATING
C980 a_4167_8527# vssd1 0.21fF $ **FLOATING
C981 a_1945_8207# vssd1 0.23fF $ **FLOATING
C982 a_25823_8207# vssd1 0.61fF $ **FLOATING
C983 a_25991_8181# vssd1 0.82fF $ **FLOATING
C984 a_25398_8207# vssd1 0.63fF $ **FLOATING
C985 a_25566_8181# vssd1 0.58fF $ **FLOATING
C986 a_25125_8213# vssd1 1.43fF $ **FLOATING
C987 a_24959_8213# vssd1 1.81fF $ **FLOATING
C988 a_23983_8207# vssd1 0.61fF $ **FLOATING
C989 a_24151_8181# vssd1 0.82fF $ **FLOATING
C990 a_23558_8207# vssd1 0.63fF $ **FLOATING
C991 a_23726_8181# vssd1 0.58fF $ **FLOATING
C992 a_23285_8213# vssd1 1.43fF $ **FLOATING
C993 _1916_.D vssd1 1.30fF $ **FLOATING
C994 a_23119_8213# vssd1 1.81fF $ **FLOATING
C995 _1580_.A vssd1 1.72fF $ **FLOATING
C996 a_22063_8426# vssd1 0.52fF $ **FLOATING
C997 a_20867_8426# vssd1 0.52fF $ **FLOATING
C998 _1582_.A vssd1 1.30fF $ **FLOATING
C999 a_20223_8426# vssd1 0.52fF $ **FLOATING
C1000 a_19388_8323# vssd1 0.50fF $ **FLOATING
C1001 a_18560_8323# vssd1 0.50fF $ **FLOATING
C1002 a_17691_8320# vssd1 0.62fF $ **FLOATING
C1003 _1040_.B vssd1 7.85fF $ **FLOATING
C1004 a_16863_8320# vssd1 0.62fF $ **FLOATING
C1005 _1146_.B vssd1 7.16fF $ **FLOATING
C1006 a_15391_8320# vssd1 0.62fF $ **FLOATING
C1007 _1109_.B vssd1 4.96fF $ **FLOATING
C1008 a_14287_8207# vssd1 0.97fF $ **FLOATING
C1009 _1149_.A1 vssd1 8.70fF $ **FLOATING
C1010 _1149_.C1 vssd1 1.73fF $ **FLOATING
C1011 a_13551_8215# vssd1 0.65fF $ **FLOATING
C1012 a_12575_8207# vssd1 0.61fF $ **FLOATING
C1013 a_12743_8181# vssd1 0.82fF $ **FLOATING
C1014 a_12150_8207# vssd1 0.63fF $ **FLOATING
C1015 a_12318_8181# vssd1 0.58fF $ **FLOATING
C1016 a_11877_8213# vssd1 1.43fF $ **FLOATING
C1017 a_11711_8213# vssd1 1.81fF $ **FLOATING
C1018 a_10643_8207# vssd1 0.61fF $ **FLOATING
C1019 a_10811_8181# vssd1 0.82fF $ **FLOATING
C1020 a_10218_8207# vssd1 0.63fF $ **FLOATING
C1021 a_10386_8181# vssd1 0.58fF $ **FLOATING
C1022 a_9945_8213# vssd1 1.43fF $ **FLOATING
C1023 _1813_.D vssd1 1.13fF $ **FLOATING
C1024 a_9779_8213# vssd1 1.81fF $ **FLOATING
C1025 _1907_.CLK vssd1 12.25fF $ **FLOATING
C1026 a_8855_8207# vssd1 0.51fF $ **FLOATING
C1027 a_8675_8207# vssd1 0.60fF $ **FLOATING
C1028 a_7843_8207# vssd1 0.51fF $ **FLOATING
C1029 a_7663_8207# vssd1 0.60fF $ **FLOATING
C1030 a_6867_8545# vssd1 0.56fF $ **FLOATING
C1031 a_5404_8323# vssd1 0.50fF $ **FLOATING
C1032 a_2455_8207# vssd1 0.61fF $ **FLOATING
C1033 a_2623_8181# vssd1 0.97fF $ **FLOATING
C1034 a_2030_8207# vssd1 0.63fF $ **FLOATING
C1035 a_2198_8181# vssd1 0.58fF $ **FLOATING
C1036 a_1757_8213# vssd1 1.43fF $ **FLOATING
C1037 a_1591_8213# vssd1 1.81fF $ **FLOATING
C1038 a_27061_8751# vssd1 0.23fF $ **FLOATING
C1039 a_27571_9117# vssd1 0.61fF $ **FLOATING
C1040 a_27739_9019# vssd1 0.82fF $ **FLOATING
C1041 a_27146_9117# vssd1 0.63fF $ **FLOATING
C1042 a_27314_8863# vssd1 0.58fF $ **FLOATING
C1043 a_26873_8751# vssd1 1.43fF $ **FLOATING
C1044 a_26707_8751# vssd1 1.81fF $ **FLOATING
C1045 a_24945_8751# vssd1 0.23fF $ **FLOATING
C1046 a_25455_9117# vssd1 0.61fF $ **FLOATING
C1047 a_25623_9019# vssd1 0.82fF $ **FLOATING
C1048 a_25030_9117# vssd1 0.63fF $ **FLOATING
C1049 a_25198_8863# vssd1 0.58fF $ **FLOATING
C1050 a_24757_8751# vssd1 1.43fF $ **FLOATING
C1051 _1924_.D vssd1 3.02fF $ **FLOATING
C1052 a_24591_8751# vssd1 1.81fF $ **FLOATING
C1053 a_23013_8751# vssd1 0.23fF $ **FLOATING
C1054 a_23523_9117# vssd1 0.61fF $ **FLOATING
C1055 a_23691_9019# vssd1 0.82fF $ **FLOATING
C1056 a_23098_9117# vssd1 0.63fF $ **FLOATING
C1057 a_23266_8863# vssd1 0.58fF $ **FLOATING
C1058 a_22825_8751# vssd1 1.43fF $ **FLOATING
C1059 _1920_.D vssd1 1.40fF $ **FLOATING
C1060 a_22659_8751# vssd1 1.81fF $ **FLOATING
C1061 _1924_.CLK vssd1 10.88fF $ **FLOATING
C1062 _1591_.X vssd1 3.50fF $ **FLOATING
C1063 _1605_.X vssd1 3.43fF $ **FLOATING
C1064 _1152_.B vssd1 5.69fF $ **FLOATING
C1065 _1062_.X vssd1 1.58fF $ **FLOATING
C1066 a_16481_8751# vssd1 0.23fF $ **FLOATING
C1067 a_21787_8916# vssd1 0.52fF $ **FLOATING
C1068 a_21143_8916# vssd1 0.52fF $ **FLOATING
C1069 a_20308_9001# vssd1 0.50fF $ **FLOATING
C1070 a_19439_8751# vssd1 0.62fF $ **FLOATING
C1071 a_17967_8751# vssd1 0.62fF $ **FLOATING
C1072 a_16991_9117# vssd1 0.61fF $ **FLOATING
C1073 a_17159_9019# vssd1 0.82fF $ **FLOATING
C1074 a_16566_9117# vssd1 0.63fF $ **FLOATING
C1075 a_16734_8863# vssd1 0.58fF $ **FLOATING
C1076 a_16293_8751# vssd1 1.43fF $ **FLOATING
C1077 a_16127_8751# vssd1 1.81fF $ **FLOATING
C1078 _1849_.CLK vssd1 10.82fF $ **FLOATING
C1079 _1059_.B vssd1 7.12fF $ **FLOATING
C1080 _1196_.C vssd1 2.74fF $ **FLOATING
C1081 _1196_.D vssd1 2.94fF $ **FLOATING
C1082 a_13488_9001# vssd1 0.26fF $ **FLOATING
C1083 _1043_.B vssd1 6.62fF $ **FLOATING
C1084 _1042_.B vssd1 4.90fF $ **FLOATING
C1085 _1362_.X vssd1 1.17fF $ **FLOATING
C1086 a_8215_8751# vssd1 0.18fF $ **FLOATING
C1087 _1058_.B vssd1 6.05fF $ **FLOATING
C1088 _1205_.Y vssd1 1.21fF $ **FLOATING
C1089 _1205_.A1 vssd1 1.08fF $ **FLOATING
C1090 a_15299_8751# vssd1 0.62fF $ **FLOATING
C1091 a_14287_9001# vssd1 0.70fF $ **FLOATING
C1092 _1060_.C1 vssd1 2.15fF $ **FLOATING
C1093 _1059_.X vssd1 1.67fF $ **FLOATING
C1094 a_13057_8897# vssd1 0.67fF $ **FLOATING
C1095 a_12171_8751# vssd1 0.62fF $ **FLOATING
C1096 a_11343_8751# vssd1 0.62fF $ **FLOATING
C1097 a_10603_9117# vssd1 0.51fF $ **FLOATING
C1098 a_10423_9117# vssd1 0.60fF $ **FLOATING
C1099 a_9595_8751# vssd1 0.62fF $ **FLOATING
C1100 _1813_.Q vssd1 2.76fF $ **FLOATING
C1101 _1165_.A vssd1 2.60fF $ **FLOATING
C1102 _1165_.C vssd1 1.81fF $ **FLOATING
C1103 a_6467_9001# vssd1 0.70fF $ **FLOATING
C1104 a_5496_9001# vssd1 0.50fF $ **FLOATING
C1105 a_4015_8779# vssd1 0.56fF $ **FLOATING
C1106 a_3063_8751# vssd1 0.62fF $ **FLOATING
C1107 a_24853_9295# vssd1 0.23fF $ **FLOATING
C1108 _1578_.X vssd1 2.66fF $ **FLOATING
C1109 _1604_.X vssd1 1.08fF $ **FLOATING
C1110 a_18180_9295# vssd1 0.26fF $ **FLOATING
C1111 _1598_.X vssd1 1.76fF $ **FLOATING
C1112 input3.X vssd1 5.65fF $ **FLOATING
C1113 a_26387_9514# vssd1 0.52fF $ **FLOATING
C1114 a_25363_9295# vssd1 0.61fF $ **FLOATING
C1115 a_25531_9269# vssd1 0.82fF $ **FLOATING
C1116 a_24938_9295# vssd1 0.63fF $ **FLOATING
C1117 a_25106_9269# vssd1 0.58fF $ **FLOATING
C1118 a_24665_9301# vssd1 1.43fF $ **FLOATING
C1119 _1678_.X vssd1 1.42fF $ **FLOATING
C1120 a_24499_9301# vssd1 1.81fF $ **FLOATING
C1121 a_23443_9514# vssd1 0.52fF $ **FLOATING
C1122 _1601_.A vssd1 1.84fF $ **FLOATING
C1123 a_22707_9514# vssd1 0.52fF $ **FLOATING
C1124 a_22063_9514# vssd1 0.52fF $ **FLOATING
C1125 a_21187_9295# vssd1 0.70fF $ **FLOATING
C1126 a_20447_9295# vssd1 0.51fF $ **FLOATING
C1127 a_20267_9295# vssd1 0.60fF $ **FLOATING
C1128 a_19112_9411# vssd1 0.50fF $ **FLOATING
C1129 _1112_.A1 vssd1 7.22fF $ **FLOATING
C1130 _1112_.B1 vssd1 2.07fF $ **FLOATING
C1131 _1112_.D1 vssd1 2.05fF $ **FLOATING
C1132 a_17749_9269# vssd1 0.67fF $ **FLOATING
C1133 a_16863_9295# vssd1 0.70fF $ **FLOATING
C1134 a_16175_9514# vssd1 0.52fF $ **FLOATING
C1135 io_in[3] vssd1 8.61fF
C1136 _1057_.X vssd1 1.75fF $ **FLOATING
C1137 a_11934_9295# vssd1 0.33fF $ **FLOATING
C1138 _1801_.Y vssd1 6.75fF $ **FLOATING
C1139 _1192_.X vssd1 2.10fF $ **FLOATING
C1140 _1759_.X vssd1 3.60fF $ **FLOATING
C1141 a_3979_9295# vssd1 0.25fF $ **FLOATING
C1142 _1210_.B vssd1 4.12fF $ **FLOATING
C1143 a_1945_9295# vssd1 0.23fF $ **FLOATING
C1144 a_15115_9408# vssd1 0.62fF $ **FLOATING
C1145 _1057_.B vssd1 5.65fF $ **FLOATING
C1146 a_14379_9408# vssd1 0.62fF $ **FLOATING
C1147 _1030_.B vssd1 5.40fF $ **FLOATING
C1148 _1801_.B vssd1 16.54fF $ **FLOATING
C1149 a_12815_9295# vssd1 1.20fF $ **FLOATING
C1150 _1192_.A2 vssd1 5.42fF $ **FLOATING
C1151 a_11777_9269# vssd1 0.72fF $ **FLOATING
C1152 a_10511_9295# vssd1 0.51fF $ **FLOATING
C1153 _1568_.B vssd1 5.03fF $ **FLOATING
C1154 a_10331_9295# vssd1 0.60fF $ **FLOATING
C1155 _1759_.A vssd1 0.90fF $ **FLOATING
C1156 a_9735_9514# vssd1 0.52fF $ **FLOATING
C1157 a_8947_9295# vssd1 0.51fF $ **FLOATING
C1158 a_8767_9295# vssd1 0.60fF $ **FLOATING
C1159 a_7980_9411# vssd1 0.50fF $ **FLOATING
C1160 _1562_.A vssd1 4.38fF $ **FLOATING
C1161 a_6559_9295# vssd1 1.20fF $ **FLOATING
C1162 a_5303_9633# vssd1 0.56fF $ **FLOATING
C1163 a_3761_9269# vssd1 0.55fF $ **FLOATING
C1164 a_2455_9295# vssd1 0.61fF $ **FLOATING
C1165 a_2623_9269# vssd1 0.97fF $ **FLOATING
C1166 a_2030_9295# vssd1 0.63fF $ **FLOATING
C1167 a_2198_9269# vssd1 0.58fF $ **FLOATING
C1168 a_1757_9301# vssd1 1.43fF $ **FLOATING
C1169 a_1591_9301# vssd1 1.81fF $ **FLOATING
C1170 a_27337_9839# vssd1 0.23fF $ **FLOATING
C1171 a_27847_10205# vssd1 0.61fF $ **FLOATING
C1172 a_28015_10107# vssd1 0.82fF $ **FLOATING
C1173 a_27422_10205# vssd1 0.63fF $ **FLOATING
C1174 a_27590_9951# vssd1 0.58fF $ **FLOATING
C1175 a_27149_9839# vssd1 1.43fF $ **FLOATING
C1176 _1926_.D vssd1 3.10fF $ **FLOATING
C1177 a_26983_9839# vssd1 1.81fF $ **FLOATING
C1178 a_25497_9839# vssd1 0.23fF $ **FLOATING
C1179 a_26007_10205# vssd1 0.61fF $ **FLOATING
C1180 a_26175_10107# vssd1 0.82fF $ **FLOATING
C1181 a_25582_10205# vssd1 0.63fF $ **FLOATING
C1182 a_25750_9951# vssd1 0.58fF $ **FLOATING
C1183 a_25309_9839# vssd1 1.43fF $ **FLOATING
C1184 _1927_.D vssd1 2.44fF $ **FLOATING
C1185 a_25143_9839# vssd1 1.81fF $ **FLOATING
C1186 _1717_.X vssd1 1.83fF $ **FLOATING
C1187 _1677_.X vssd1 2.94fF $ **FLOATING
C1188 _1590_.X vssd1 1.41fF $ **FLOATING
C1189 a_23667_10205# vssd1 0.51fF $ **FLOATING
C1190 a_23487_10205# vssd1 0.60fF $ **FLOATING
C1191 a_22747_10205# vssd1 0.51fF $ **FLOATING
C1192 a_22567_10205# vssd1 0.60fF $ **FLOATING
C1193 a_21827_10205# vssd1 0.51fF $ **FLOATING
C1194 a_21647_10205# vssd1 0.60fF $ **FLOATING
C1195 a_20815_10205# vssd1 0.51fF $ **FLOATING
C1196 a_20635_10205# vssd1 0.60fF $ **FLOATING
C1197 _1590_.A_N vssd1 15.42fF $ **FLOATING
C1198 a_19439_9839# vssd1 0.65fF $ **FLOATING
C1199 _0993_.X vssd1 7.99fF $ **FLOATING
C1200 a_7749_9839# vssd1 0.17fF $ **FLOATING
C1201 a_14641_9839# vssd1 0.23fF $ **FLOATING
C1202 a_18059_9839# vssd1 0.70fF $ **FLOATING
C1203 a_17139_9839# vssd1 1.20fF $ **FLOATING
C1204 a_16159_9867# vssd1 0.56fF $ **FLOATING
C1205 a_15151_10205# vssd1 0.61fF $ **FLOATING
C1206 a_15319_10107# vssd1 0.82fF $ **FLOATING
C1207 a_14726_10205# vssd1 0.63fF $ **FLOATING
C1208 a_14894_9951# vssd1 0.58fF $ **FLOATING
C1209 a_14453_9839# vssd1 1.43fF $ **FLOATING
C1210 a_14287_9839# vssd1 1.81fF $ **FLOATING
C1211 _1069_.C vssd1 3.61fF $ **FLOATING
C1212 _1069_.D vssd1 1.90fF $ **FLOATING
C1213 _1069_.B vssd1 1.25fF $ **FLOATING
C1214 a_11842_10089# vssd1 0.33fF $ **FLOATING
C1215 a_10452_10089# vssd1 0.26fF $ **FLOATING
C1216 a_4669_9839# vssd1 0.19fF $ **FLOATING
C1217 _1083_.A vssd1 5.61fF $ **FLOATING
C1218 _1563_.X vssd1 2.90fF $ **FLOATING
C1219 _1159_.X vssd1 14.15fF $ **FLOATING
C1220 a_6645_10089# vssd1 0.24fF $ **FLOATING
C1221 _1172_.X vssd1 2.35fF $ **FLOATING
C1222 a_2405_9839# vssd1 0.23fF $ **FLOATING
C1223 a_12723_10089# vssd1 0.70fF $ **FLOATING
C1224 _0992_.A2 vssd1 5.84fF $ **FLOATING
C1225 a_11685_9813# vssd1 0.72fF $ **FLOATING
C1226 _1011_.A1 vssd1 4.47fF $ **FLOATING
C1227 _1011_.B1 vssd1 2.80fF $ **FLOATING
C1228 a_10021_9985# vssd1 0.67fF $ **FLOATING
C1229 a_9176_10089# vssd1 0.50fF $ **FLOATING
C1230 _1563_.A vssd1 1.00fF $ **FLOATING
C1231 a_8447_10004# vssd1 0.52fF $ **FLOATING
C1232 a_7531_9813# vssd1 0.55fF $ **FLOATING
C1233 a_5639_10089# vssd1 0.70fF $ **FLOATING
C1234 a_4519_9991# vssd1 0.74fF $ **FLOATING
C1235 a_3095_9867# vssd1 0.56fF $ **FLOATING
C1236 a_2228_9839# vssd1 0.50fF $ **FLOATING
C1237 a_2122_9839# vssd1 0.58fF $ **FLOATING
C1238 a_1945_9839# vssd1 0.50fF $ **FLOATING
C1239 a_1626_9839# vssd1 0.54fF $ **FLOATING
C1240 io_in[4] vssd1 1.35fF
C1241 _1728_.X vssd1 3.14fF $ **FLOATING
C1242 _1720_.X vssd1 2.04fF $ **FLOATING
C1243 a_24025_10383# vssd1 0.23fF $ **FLOATING
C1244 _1602_.X vssd1 3.19fF $ **FLOATING
C1245 _1008_.X vssd1 2.93fF $ **FLOATING
C1246 a_26203_10602# vssd1 0.52fF $ **FLOATING
C1247 _1720_.A vssd1 2.00fF $ **FLOATING
C1248 a_25559_10602# vssd1 0.52fF $ **FLOATING
C1249 a_24535_10383# vssd1 0.61fF $ **FLOATING
C1250 a_24703_10357# vssd1 0.82fF $ **FLOATING
C1251 a_24110_10383# vssd1 0.63fF $ **FLOATING
C1252 a_24278_10357# vssd1 0.58fF $ **FLOATING
C1253 a_23837_10389# vssd1 1.43fF $ **FLOATING
C1254 a_23671_10389# vssd1 1.81fF $ **FLOATING
C1255 a_22935_10383# vssd1 0.70fF $ **FLOATING
C1256 a_22195_10383# vssd1 0.51fF $ **FLOATING
C1257 _1719_.B vssd1 6.41fF $ **FLOATING
C1258 a_22015_10383# vssd1 0.60fF $ **FLOATING
C1259 a_20676_10499# vssd1 0.50fF $ **FLOATING
C1260 a_19807_10496# vssd1 0.62fF $ **FLOATING
C1261 _1129_.B vssd1 6.73fF $ **FLOATING
C1262 a_18979_10496# vssd1 0.62fF $ **FLOATING
C1263 _1182_.B vssd1 5.34fF $ **FLOATING
C1264 a_18151_10496# vssd1 0.62fF $ **FLOATING
C1265 _1080_.B vssd1 6.59fF $ **FLOATING
C1266 a_16863_10496# vssd1 0.62fF $ **FLOATING
C1267 _1089_.B vssd1 5.64fF $ **FLOATING
C1268 a_15943_10496# vssd1 0.62fF $ **FLOATING
C1269 _1102_.B vssd1 6.49fF $ **FLOATING
C1270 a_14839_10499# vssd1 0.70fF $ **FLOATING
C1271 _1008_.A vssd1 2.42fF $ **FLOATING
C1272 _1008_.B vssd1 2.52fF $ **FLOATING
C1273 a_12525_10383# vssd1 0.23fF $ **FLOATING
C1274 a_6997_10383# vssd1 0.23fF $ **FLOATING
C1275 a_6743_10383# vssd1 0.39fF $ **FLOATING
C1276 _1561_.X vssd1 2.74fF $ **FLOATING
C1277 _1126_.Y vssd1 15.16fF $ **FLOATING
C1278 a_6743_10703# vssd1 0.59fF $ **FLOATING
C1279 _1317_.X vssd1 4.99fF $ **FLOATING
C1280 a_14103_10383# vssd1 0.70fF $ **FLOATING
C1281 a_13035_10383# vssd1 0.61fF $ **FLOATING
C1282 a_13203_10357# vssd1 0.82fF $ **FLOATING
C1283 a_12610_10383# vssd1 0.63fF $ **FLOATING
C1284 a_12778_10357# vssd1 0.58fF $ **FLOATING
C1285 a_12337_10389# vssd1 1.43fF $ **FLOATING
C1286 _1848_.D vssd1 1.58fF $ **FLOATING
C1287 a_12171_10389# vssd1 1.81fF $ **FLOATING
C1288 a_10839_10602# vssd1 0.52fF $ **FLOATING
C1289 a_9871_10391# vssd1 0.65fF $ **FLOATING
C1290 _1532_.A vssd1 12.43fF $ **FLOATING
C1291 a_9275_10602# vssd1 0.52fF $ **FLOATING
C1292 a_8440_10499# vssd1 0.50fF $ **FLOATING
C1293 a_5087_10496# vssd1 0.62fF $ **FLOATING
C1294 a_2686_10383# vssd1 4.03fF $ **FLOATING
C1295 a_1775_10496# vssd1 0.62fF $ **FLOATING
C1296 a_27245_10927# vssd1 0.23fF $ **FLOATING
C1297 a_27755_11293# vssd1 0.61fF $ **FLOATING
C1298 a_27923_11195# vssd1 0.82fF $ **FLOATING
C1299 a_27330_11293# vssd1 0.63fF $ **FLOATING
C1300 a_27498_11039# vssd1 0.58fF $ **FLOATING
C1301 a_27057_10927# vssd1 1.43fF $ **FLOATING
C1302 a_26891_10927# vssd1 1.81fF $ **FLOATING
C1303 a_25221_10927# vssd1 0.23fF $ **FLOATING
C1304 a_25731_11293# vssd1 0.61fF $ **FLOATING
C1305 a_25899_11195# vssd1 0.82fF $ **FLOATING
C1306 a_25306_11293# vssd1 0.63fF $ **FLOATING
C1307 a_25474_11039# vssd1 0.58fF $ **FLOATING
C1308 a_25033_10927# vssd1 1.43fF $ **FLOATING
C1309 a_24867_10927# vssd1 1.81fF $ **FLOATING
C1310 a_23013_10927# vssd1 0.23fF $ **FLOATING
C1311 a_23523_11293# vssd1 0.61fF $ **FLOATING
C1312 a_23691_11195# vssd1 0.82fF $ **FLOATING
C1313 a_23098_11293# vssd1 0.63fF $ **FLOATING
C1314 a_23266_11039# vssd1 0.58fF $ **FLOATING
C1315 a_22825_10927# vssd1 1.43fF $ **FLOATING
C1316 a_22659_10927# vssd1 1.81fF $ **FLOATING
C1317 _1587_.X vssd1 2.92fF $ **FLOATING
C1318 _0973_.B vssd1 6.37fF $ **FLOATING
C1319 _1584_.X vssd1 3.65fF $ **FLOATING
C1320 _1155_.C vssd1 3.24fF $ **FLOATING
C1321 _1155_.B vssd1 3.14fF $ **FLOATING
C1322 _1037_.B vssd1 6.19fF $ **FLOATING
C1323 _1088_.B vssd1 6.94fF $ **FLOATING
C1324 a_10331_10927# vssd1 0.18fF $ **FLOATING
C1325 _1197_.D vssd1 2.22fF $ **FLOATING
C1326 _1197_.B vssd1 3.56fF $ **FLOATING
C1327 a_12384_11177# vssd1 0.26fF $ **FLOATING
C1328 _1439_.X vssd1 3.93fF $ **FLOATING
C1329 _1560_.X vssd1 1.02fF $ **FLOATING
C1330 a_4253_10927# vssd1 0.17fF $ **FLOATING
C1331 a_2897_10927# vssd1 0.44fF $ **FLOATING
C1332 a_8325_10901# vssd1 0.61fF $ **FLOATING
C1333 _1162_.X vssd1 2.73fF $ **FLOATING
C1334 a_6277_11177# vssd1 0.24fF $ **FLOATING
C1335 _1797_.Y vssd1 2.99fF $ **FLOATING
C1336 _1684_.A vssd1 1.57fF $ **FLOATING
C1337 a_22063_11092# vssd1 0.52fF $ **FLOATING
C1338 a_21136_11177# vssd1 0.50fF $ **FLOATING
C1339 a_20267_10927# vssd1 0.62fF $ **FLOATING
C1340 a_19480_11177# vssd1 0.50fF $ **FLOATING
C1341 a_18607_11293# vssd1 0.51fF $ **FLOATING
C1342 a_18427_11293# vssd1 0.60fF $ **FLOATING
C1343 _1583_.X vssd1 1.00fF $ **FLOATING
C1344 a_17831_11092# vssd1 0.52fF $ **FLOATING
C1345 a_16863_11177# vssd1 0.70fF $ **FLOATING
C1346 a_16035_10927# vssd1 0.62fF $ **FLOATING
C1347 a_15207_10927# vssd1 0.62fF $ **FLOATING
C1348 a_14467_11293# vssd1 0.51fF $ **FLOATING
C1349 a_14287_11293# vssd1 0.60fF $ **FLOATING
C1350 a_13183_11177# vssd1 0.70fF $ **FLOATING
C1351 _1572_.B vssd1 2.99fF $ **FLOATING
C1352 _1045_.B1 vssd1 1.78fF $ **FLOATING
C1353 _1045_.C1 vssd1 1.67fF $ **FLOATING
C1354 a_11953_11073# vssd1 0.67fF $ **FLOATING
C1355 a_11299_11092# vssd1 0.52fF $ **FLOATING
C1356 _1051_.A1 vssd1 4.40fF $ **FLOATING
C1357 a_9591_11293# vssd1 0.51fF $ **FLOATING
C1358 a_9411_11293# vssd1 0.60fF $ **FLOATING
C1359 a_7896_11079# vssd1 0.59fF $ **FLOATING
C1360 a_5361_11191# vssd1 0.60fF $ **FLOATING
C1361 a_5261_10973# vssd1 0.49fF $ **FLOATING
C1362 a_3065_11177# vssd1 0.39fF $ **FLOATING
C1363 _1207_.B1_N vssd1 5.35fF $ **FLOATING
C1364 a_1814_11177# vssd1 0.33fF $ **FLOATING
C1365 _1226_.A2 vssd1 3.61fF $ **FLOATING
C1366 a_4035_10901# vssd1 0.55fF $ **FLOATING
C1367 _1226_.A1 vssd1 5.54fF $ **FLOATING
C1368 _1226_.B1 vssd1 6.21fF $ **FLOATING
C1369 a_2696_11177# vssd1 0.63fF $ **FLOATING
C1370 _1170_.B2 vssd1 3.19fF $ **FLOATING
C1371 _1170_.B1 vssd1 3.90fF $ **FLOATING
C1372 _1170_.A2 vssd1 15.36fF $ **FLOATING
C1373 _1170_.A3 vssd1 15.38fF $ **FLOATING
C1374 a_1657_10901# vssd1 0.72fF $ **FLOATING
C1375 _1716_.X vssd1 2.54fF $ **FLOATING
C1376 a_24025_11471# vssd1 0.23fF $ **FLOATING
C1377 _1680_.X vssd1 1.91fF $ **FLOATING
C1378 a_20437_11471# vssd1 0.23fF $ **FLOATING
C1379 _1586_.X vssd1 4.52fF $ **FLOATING
C1380 a_16064_11471# vssd1 0.26fF $ **FLOATING
C1381 a_13999_11471# vssd1 0.35fF $ **FLOATING
C1382 a_13805_11471# vssd1 0.25fF $ **FLOATING
C1383 a_13551_11471# vssd1 0.38fF $ **FLOATING
C1384 a_10227_11471# vssd1 0.38fF $ **FLOATING
C1385 a_9779_11471# vssd1 0.38fF $ **FLOATING
C1386 a_7656_11471# vssd1 0.17fF $ **FLOATING
C1387 a_12065_11471# vssd1 0.23fF $ **FLOATING
C1388 a_9779_11791# vssd1 0.55fF $ **FLOATING
C1389 a_8955_11791# vssd1 0.27fF $ **FLOATING
C1390 a_7573_11791# vssd1 0.42fF $ **FLOATING
C1391 _1125_.X vssd1 3.95fF $ **FLOATING
C1392 a_5451_11471# vssd1 0.25fF $ **FLOATING
C1393 a_27623_11471# vssd1 0.51fF $ **FLOATING
C1394 a_27443_11471# vssd1 0.60fF $ **FLOATING
C1395 a_26479_11690# vssd1 0.52fF $ **FLOATING
C1396 a_24535_11471# vssd1 0.61fF $ **FLOATING
C1397 a_24703_11445# vssd1 0.82fF $ **FLOATING
C1398 a_24110_11471# vssd1 0.63fF $ **FLOATING
C1399 a_24278_11445# vssd1 0.58fF $ **FLOATING
C1400 a_23837_11477# vssd1 1.43fF $ **FLOATING
C1401 _1966_.D vssd1 1.80fF $ **FLOATING
C1402 a_23671_11477# vssd1 1.81fF $ **FLOATING
C1403 a_23075_11690# vssd1 0.52fF $ **FLOATING
C1404 a_22015_11471# vssd1 0.70fF $ **FLOATING
C1405 a_20947_11471# vssd1 0.61fF $ **FLOATING
C1406 a_21115_11445# vssd1 0.82fF $ **FLOATING
C1407 a_20522_11471# vssd1 0.63fF $ **FLOATING
C1408 a_20690_11445# vssd1 0.58fF $ **FLOATING
C1409 a_20249_11477# vssd1 1.43fF $ **FLOATING
C1410 a_20083_11477# vssd1 1.81fF $ **FLOATING
C1411 _1586_.A vssd1 1.20fF $ **FLOATING
C1412 a_19487_11690# vssd1 0.52fF $ **FLOATING
C1413 a_18551_11809# vssd1 0.56fF $ **FLOATING
C1414 a_17139_11584# vssd1 0.62fF $ **FLOATING
C1415 _1119_.A1 vssd1 7.00fF $ **FLOATING
C1416 _1119_.C1 vssd1 4.48fF $ **FLOATING
C1417 _1118_.X vssd1 1.33fF $ **FLOATING
C1418 a_15633_11445# vssd1 0.67fF $ **FLOATING
C1419 a_14839_11471# vssd1 0.70fF $ **FLOATING
C1420 _1156_.D vssd1 2.34fF $ **FLOATING
C1421 _1156_.C vssd1 3.78fF $ **FLOATING
C1422 a_12575_11471# vssd1 0.61fF $ **FLOATING
C1423 a_12743_11445# vssd1 0.82fF $ **FLOATING
C1424 a_12150_11471# vssd1 0.63fF $ **FLOATING
C1425 a_12318_11445# vssd1 0.58fF $ **FLOATING
C1426 a_11877_11477# vssd1 1.43fF $ **FLOATING
C1427 a_11711_11477# vssd1 1.81fF $ **FLOATING
C1428 _1121_.A1 vssd1 8.33fF $ **FLOATING
C1429 a_8818_11703# vssd1 0.60fF $ **FLOATING
C1430 _1164_.A2 vssd1 2.54fF $ **FLOATING
C1431 _1156_.Y vssd1 5.20fF $ **FLOATING
C1432 a_6651_11587# vssd1 0.70fF $ **FLOATING
C1433 _1124_.X vssd1 2.37fF $ **FLOATING
C1434 _1796_.X vssd1 5.87fF $ **FLOATING
C1435 _1782_.X vssd1 6.01fF $ **FLOATING
C1436 a_5233_11445# vssd1 0.55fF $ **FLOATING
C1437 _1177_.B vssd1 4.50fF $ **FLOATING
C1438 _1177_.C vssd1 6.53fF $ **FLOATING
C1439 a_2644_11587# vssd1 0.50fF $ **FLOATING
C1440 _1221_.A vssd1 6.50fF $ **FLOATING
C1441 _1221_.B vssd1 5.54fF $ **FLOATING
C1442 a_1816_11587# vssd1 0.50fF $ **FLOATING
C1443 _1782_.A vssd1 13.75fF $ **FLOATING
C1444 a_27337_12015# vssd1 0.23fF $ **FLOATING
C1445 a_27847_12381# vssd1 0.61fF $ **FLOATING
C1446 a_28015_12283# vssd1 0.82fF $ **FLOATING
C1447 a_27422_12381# vssd1 0.63fF $ **FLOATING
C1448 a_27590_12127# vssd1 0.58fF $ **FLOATING
C1449 a_27149_12015# vssd1 1.43fF $ **FLOATING
C1450 a_26983_12015# vssd1 1.81fF $ **FLOATING
C1451 _1978_.D vssd1 1.85fF $ **FLOATING
C1452 _1727_.X vssd1 2.50fF $ **FLOATING
C1453 _1680_.A vssd1 0.97fF $ **FLOATING
C1454 _1681_.X vssd1 2.45fF $ **FLOATING
C1455 _1577_.X vssd1 2.37fF $ **FLOATING
C1456 _1577_.B vssd1 11.17fF $ **FLOATING
C1457 _1135_.B vssd1 5.79fF $ **FLOATING
C1458 _1128_.B vssd1 6.22fF $ **FLOATING
C1459 _1098_.B vssd1 7.48fF $ **FLOATING
C1460 _0991_.X vssd1 5.03fF $ **FLOATING
C1461 _1025_.B vssd1 3.53fF $ **FLOATING
C1462 _1438_.X vssd1 1.53fF $ **FLOATING
C1463 a_10515_12015# vssd1 0.18fF $ **FLOATING
C1464 a_8178_12015# vssd1 0.20fF $ **FLOATING
C1465 _1847_.D vssd1 1.22fF $ **FLOATING
C1466 _1571_.X vssd1 4.03fF $ **FLOATING
C1467 _1086_.Y vssd1 6.05fF $ **FLOATING
C1468 a_7019_12265# vssd1 0.39fF $ **FLOATING
C1469 a_4713_12015# vssd1 0.17fF $ **FLOATING
C1470 _1321_.C vssd1 12.35fF $ **FLOATING
C1471 a_1857_12265# vssd1 0.21fF $ **FLOATING
C1472 a_24639_12180# vssd1 0.52fF $ **FLOATING
C1473 a_23483_12381# vssd1 0.51fF $ **FLOATING
C1474 a_23303_12381# vssd1 0.60fF $ **FLOATING
C1475 a_22563_12381# vssd1 0.51fF $ **FLOATING
C1476 a_22383_12381# vssd1 0.60fF $ **FLOATING
C1477 a_21643_12381# vssd1 0.51fF $ **FLOATING
C1478 a_21463_12381# vssd1 0.60fF $ **FLOATING
C1479 a_20676_12265# vssd1 0.50fF $ **FLOATING
C1480 a_19439_12015# vssd1 0.62fF $ **FLOATING
C1481 a_18243_12015# vssd1 0.62fF $ **FLOATING
C1482 a_17323_12015# vssd1 0.62fF $ **FLOATING
C1483 a_16495_12015# vssd1 0.62fF $ **FLOATING
C1484 a_15607_12043# vssd1 0.56fF $ **FLOATING
C1485 a_14747_12015# vssd1 0.62fF $ **FLOATING
C1486 _1569_.A vssd1 2.76fF $ **FLOATING
C1487 a_13047_12180# vssd1 0.52fF $ **FLOATING
C1488 a_12259_12381# vssd1 0.51fF $ **FLOATING
C1489 _1438_.B vssd1 2.59fF $ **FLOATING
C1490 a_12079_12381# vssd1 0.60fF $ **FLOATING
C1491 a_11299_12180# vssd1 0.52fF $ **FLOATING
C1492 _1015_.A1 vssd1 3.27fF $ **FLOATING
C1493 a_9779_12015# vssd1 0.70fF $ **FLOATING
C1494 a_9183_12180# vssd1 0.52fF $ **FLOATING
C1495 _1084_.C1 vssd1 7.26fF $ **FLOATING
C1496 _1084_.B1 vssd1 1.93fF $ **FLOATING
C1497 _1084_.A1 vssd1 3.72fF $ **FLOATING
C1498 a_7993_11989# vssd1 0.89fF $ **FLOATING
C1499 _1086_.B vssd1 4.78fF $ **FLOATING
C1500 _1086_.A vssd1 4.49fF $ **FLOATING
C1501 a_5547_12015# vssd1 0.62fF $ **FLOATING
C1502 _1216_.A2 vssd1 1.96fF $ **FLOATING
C1503 a_4495_11989# vssd1 0.55fF $ **FLOATING
C1504 a_1775_12265# vssd1 0.80fF $ **FLOATING
C1505 _1177_.Y vssd1 2.81fF $ **FLOATING
C1506 _1208_.A1 vssd1 7.31fF $ **FLOATING
C1507 _1715_.X vssd1 1.46fF $ **FLOATING
C1508 a_25589_12559# vssd1 0.23fF $ **FLOATING
C1509 a_22504_12559# vssd1 0.26fF $ **FLOATING
C1510 _1154_.X vssd1 3.60fF $ **FLOATING
C1511 a_20081_12559# vssd1 0.20fF $ **FLOATING
C1512 a_19069_12559# vssd1 0.20fF $ **FLOATING
C1513 a_17029_12559# vssd1 0.21fF $ **FLOATING
C1514 a_16945_12559# vssd1 0.17fF $ **FLOATING
C1515 a_15512_12559# vssd1 0.26fF $ **FLOATING
C1516 _0999_.X vssd1 2.57fF $ **FLOATING
C1517 _1573_.X vssd1 3.93fF $ **FLOATING
C1518 a_12893_12559# vssd1 0.23fF $ **FLOATING
C1519 a_8395_12559# vssd1 0.25fF $ **FLOATING
C1520 a_6981_12559# vssd1 0.39fF $ **FLOATING
C1521 a_6559_12559# vssd1 0.86fF $ **FLOATING
C1522 _1013_.X vssd1 1.38fF $ **FLOATING
C1523 _1158_.X vssd1 3.53fF $ **FLOATING
C1524 a_28135_12778# vssd1 0.52fF $ **FLOATING
C1525 a_27347_12559# vssd1 0.51fF $ **FLOATING
C1526 a_27167_12559# vssd1 0.60fF $ **FLOATING
C1527 a_26099_12559# vssd1 0.61fF $ **FLOATING
C1528 a_26267_12533# vssd1 0.82fF $ **FLOATING
C1529 a_25674_12559# vssd1 0.63fF $ **FLOATING
C1530 a_25842_12533# vssd1 0.58fF $ **FLOATING
C1531 a_25401_12565# vssd1 1.43fF $ **FLOATING
C1532 _1965_.D vssd1 3.15fF $ **FLOATING
C1533 a_25235_12565# vssd1 1.81fF $ **FLOATING
C1534 a_24039_12559# vssd1 0.70fF $ **FLOATING
C1535 fanout24.A vssd1 10.40fF $ **FLOATING
C1536 a_23443_12778# vssd1 0.52fF $ **FLOATING
C1537 _1154_.A1 vssd1 2.98fF $ **FLOATING
C1538 _1154_.C1 vssd1 3.26fF $ **FLOATING
C1539 a_22073_12533# vssd1 0.67fF $ **FLOATING
C1540 a_21127_12897# vssd1 0.56fF $ **FLOATING
C1541 _1183_.B1 vssd1 2.52fF $ **FLOATING
C1542 _1183_.A2 vssd1 8.28fF $ **FLOATING
C1543 a_19952_12533# vssd1 0.65fF $ **FLOATING
C1544 _0974_.B1 vssd1 1.77fF $ **FLOATING
C1545 _0974_.A2 vssd1 6.16fF $ **FLOATING
C1546 a_18940_12533# vssd1 0.65fF $ **FLOATING
C1547 a_17967_12672# vssd1 0.62fF $ **FLOATING
C1548 _1965_.Q vssd1 6.19fF $ **FLOATING
C1549 a_16863_12559# vssd1 0.97fF $ **FLOATING
C1550 _0999_.C1 vssd1 3.83fF $ **FLOATING
C1551 _1103_.A1 vssd1 9.63fF $ **FLOATING
C1552 _1103_.D1 vssd1 1.88fF $ **FLOATING
C1553 a_15081_12533# vssd1 0.67fF $ **FLOATING
C1554 _1573_.A vssd1 1.40fF $ **FLOATING
C1555 a_14427_12778# vssd1 0.52fF $ **FLOATING
C1556 a_13403_12559# vssd1 0.61fF $ **FLOATING
C1557 a_13571_12533# vssd1 0.82fF $ **FLOATING
C1558 a_12978_12559# vssd1 0.63fF $ **FLOATING
C1559 a_13146_12533# vssd1 0.58fF $ **FLOATING
C1560 a_12705_12565# vssd1 1.43fF $ **FLOATING
C1561 _1911_.D vssd1 1.05fF $ **FLOATING
C1562 a_12539_12565# vssd1 1.81fF $ **FLOATING
C1563 a_11711_12672# vssd1 0.62fF $ **FLOATING
C1564 _1092_.B vssd1 5.28fF $ **FLOATING
C1565 a_10648_12675# vssd1 0.50fF $ **FLOATING
C1566 a_9879_12675# vssd1 0.48fF $ **FLOATING
C1567 a_9687_12919# vssd1 0.48fF $ **FLOATING
C1568 _1794_.Y vssd1 2.68fF $ **FLOATING
C1569 a_4351_12559# vssd1 0.61fF $ **FLOATING
C1570 _1123_.X vssd1 4.80fF $ **FLOATING
C1571 a_4601_12879# vssd1 0.16fF $ **FLOATING
C1572 a_4351_12879# vssd1 0.19fF $ **FLOATING
C1573 a_2331_12879# vssd1 0.21fF $ **FLOATING
C1574 a_8177_12533# vssd1 0.55fF $ **FLOATING
C1575 _0903_.C vssd1 2.67fF $ **FLOATING
C1576 a_5731_12567# vssd1 0.65fF $ **FLOATING
C1577 _1252_.A vssd1 1.29fF $ **FLOATING
C1578 a_3247_12672# vssd1 0.62fF $ **FLOATING
C1579 _1222_.B1 vssd1 1.20fF $ **FLOATING
C1580 _1222_.A1 vssd1 5.74fF $ **FLOATING
C1581 a_2195_12533# vssd1 0.79fF $ **FLOATING
C1582 a_26785_13103# vssd1 0.23fF $ **FLOATING
C1583 a_27295_13469# vssd1 0.61fF $ **FLOATING
C1584 a_27463_13371# vssd1 0.82fF $ **FLOATING
C1585 a_26870_13469# vssd1 0.63fF $ **FLOATING
C1586 a_27038_13215# vssd1 0.58fF $ **FLOATING
C1587 a_26597_13103# vssd1 1.43fF $ **FLOATING
C1588 a_26431_13103# vssd1 1.81fF $ **FLOATING
C1589 a_24945_13103# vssd1 0.23fF $ **FLOATING
C1590 a_25455_13469# vssd1 0.61fF $ **FLOATING
C1591 a_25623_13371# vssd1 0.82fF $ **FLOATING
C1592 a_25030_13469# vssd1 0.63fF $ **FLOATING
C1593 a_25198_13215# vssd1 0.58fF $ **FLOATING
C1594 a_24757_13103# vssd1 1.43fF $ **FLOATING
C1595 _1980_.D vssd1 2.28fF $ **FLOATING
C1596 a_24591_13103# vssd1 1.81fF $ **FLOATING
C1597 _1709_.X vssd1 1.88fF $ **FLOATING
C1598 _1079_.B vssd1 4.37fF $ **FLOATING
C1599 _1007_.X vssd1 4.25fF $ **FLOATING
C1600 a_20157_13353# vssd1 0.21fF $ **FLOATING
C1601 a_20073_13353# vssd1 0.17fF $ **FLOATING
C1602 _1147_.X vssd1 1.83fF $ **FLOATING
C1603 a_17305_13353# vssd1 0.21fF $ **FLOATING
C1604 a_17221_13353# vssd1 0.17fF $ **FLOATING
C1605 _0997_.X vssd1 7.02fF $ **FLOATING
C1606 a_13165_13103# vssd1 0.21fF $ **FLOATING
C1607 _1120_.X vssd1 4.18fF $ **FLOATING
C1608 _1120_.D vssd1 1.78fF $ **FLOATING
C1609 _1120_.B vssd1 3.67fF $ **FLOATING
C1610 _1570_.X vssd1 2.42fF $ **FLOATING
C1611 _1436_.X vssd1 1.90fF $ **FLOATING
C1612 a_9323_13103# vssd1 0.27fF $ **FLOATING
C1613 a_7381_13103# vssd1 0.21fF $ **FLOATING
C1614 a_8031_13353# vssd1 0.44fF $ **FLOATING
C1615 _1791_.Y vssd1 6.60fF $ **FLOATING
C1616 a_23759_13469# vssd1 0.51fF $ **FLOATING
C1617 _1685_.B vssd1 6.01fF $ **FLOATING
C1618 a_23579_13469# vssd1 0.60fF $ **FLOATING
C1619 _1685_.A_N vssd1 12.90fF $ **FLOATING
C1620 a_22563_13469# vssd1 0.51fF $ **FLOATING
C1621 _1977_.Q vssd1 6.60fF $ **FLOATING
C1622 a_22383_13469# vssd1 0.60fF $ **FLOATING
C1623 a_21095_13103# vssd1 0.62fF $ **FLOATING
C1624 a_19991_13103# vssd1 0.97fF $ **FLOATING
C1625 _1007_.A1 vssd1 4.41fF $ **FLOATING
C1626 a_18459_13131# vssd1 0.56fF $ **FLOATING
C1627 a_17139_13103# vssd1 0.97fF $ **FLOATING
C1628 _1147_.C1 vssd1 2.49fF $ **FLOATING
C1629 a_15883_13131# vssd1 0.56fF $ **FLOATING
C1630 a_14287_13353# vssd1 0.70fF $ **FLOATING
C1631 a_12927_13103# vssd1 0.71fF $ **FLOATING
C1632 a_11752_13353# vssd1 0.50fF $ **FLOATING
C1633 a_10971_13469# vssd1 0.51fF $ **FLOATING
C1634 _1436_.B vssd1 4.20fF $ **FLOATING
C1635 a_10791_13469# vssd1 0.60fF $ **FLOATING
C1636 a_10195_13268# vssd1 0.52fF $ **FLOATING
C1637 _1198_.A1 vssd1 6.82fF $ **FLOATING
C1638 _1198_.A2 vssd1 6.80fF $ **FLOATING
C1639 _1198_.B2 vssd1 3.36fF $ **FLOATING
C1640 a_9186_13255# vssd1 0.60fF $ **FLOATING
C1641 _1052_.B1 vssd1 3.47fF $ **FLOATING
C1642 a_7189_13408# vssd1 0.45fF $ **FLOATING
C1643 _1795_.X vssd1 1.81fF $ **FLOATING
C1644 a_6324_13353# vssd1 0.50fF $ **FLOATING
C1645 a_5269_13367# vssd1 0.60fF $ **FLOATING
C1646 a_5169_13149# vssd1 0.49fF $ **FLOATING
C1647 a_4259_13103# vssd1 0.65fF $ **FLOATING
C1648 a_2037_13103# vssd1 0.23fF $ **FLOATING
C1649 a_2547_13469# vssd1 0.61fF $ **FLOATING
C1650 a_2715_13371# vssd1 0.97fF $ **FLOATING
C1651 a_2122_13469# vssd1 0.63fF $ **FLOATING
C1652 a_2290_13215# vssd1 0.58fF $ **FLOATING
C1653 a_1849_13103# vssd1 1.43fF $ **FLOATING
C1654 a_1683_13103# vssd1 1.81fF $ **FLOATING
C1655 _2023_.CLK vssd1 15.15fF $ **FLOATING
C1656 _1713_.X vssd1 1.30fF $ **FLOATING
C1657 a_25589_13647# vssd1 0.23fF $ **FLOATING
C1658 _1711_.X vssd1 1.02fF $ **FLOATING
C1659 a_22238_13647# vssd1 0.33fF $ **FLOATING
C1660 a_20065_13647# vssd1 0.21fF $ **FLOATING
C1661 a_19981_13647# vssd1 0.17fF $ **FLOATING
C1662 _1006_.X vssd1 1.71fF $ **FLOATING
C1663 _1191_.X vssd1 5.02fF $ **FLOATING
C1664 a_14643_13647# vssd1 0.35fF $ **FLOATING
C1665 a_14449_13647# vssd1 0.25fF $ **FLOATING
C1666 a_14195_13647# vssd1 0.38fF $ **FLOATING
C1667 _1050_.Y vssd1 5.30fF $ **FLOATING
C1668 _1755_.X vssd1 8.73fF $ **FLOATING
C1669 a_10791_13647# vssd1 0.39fF $ **FLOATING
C1670 a_8387_13647# vssd1 0.38fF $ **FLOATING
C1671 a_7939_13647# vssd1 0.38fF $ **FLOATING
C1672 a_5241_13647# vssd1 0.29fF $ **FLOATING
C1673 a_4709_13647# vssd1 0.53fF $ **FLOATING
C1674 a_12065_13647# vssd1 0.23fF $ **FLOATING
C1675 _1434_.X vssd1 1.90fF $ **FLOATING
C1676 _1175_.Y vssd1 5.07fF $ **FLOATING
C1677 a_7939_13967# vssd1 0.55fF $ **FLOATING
C1678 a_6747_13967# vssd1 0.27fF $ **FLOATING
C1679 a_4877_13967# vssd1 0.16fF $ **FLOATING
C1680 a_4627_13967# vssd1 0.25fF $ **FLOATING
C1681 a_3247_13967# vssd1 0.29fF $ **FLOATING
C1682 a_1791_13967# vssd1 0.33fF $ **FLOATING
C1683 _1703_.A vssd1 1.64fF $ **FLOATING
C1684 a_28135_13866# vssd1 0.52fF $ **FLOATING
C1685 a_27347_13647# vssd1 0.51fF $ **FLOATING
C1686 a_27167_13647# vssd1 0.60fF $ **FLOATING
C1687 a_26099_13647# vssd1 0.61fF $ **FLOATING
C1688 a_26267_13621# vssd1 0.82fF $ **FLOATING
C1689 a_25674_13647# vssd1 0.63fF $ **FLOATING
C1690 a_25842_13621# vssd1 0.58fF $ **FLOATING
C1691 a_25401_13653# vssd1 1.43fF $ **FLOATING
C1692 _1986_.D vssd1 2.80fF $ **FLOATING
C1693 a_25235_13653# vssd1 1.81fF $ **FLOATING
C1694 _1686_.A vssd1 0.92fF $ **FLOATING
C1695 a_24087_13866# vssd1 0.52fF $ **FLOATING
C1696 a_23299_13647# vssd1 0.51fF $ **FLOATING
C1697 a_23119_13647# vssd1 0.60fF $ **FLOATING
C1698 _1006_.B2 vssd1 3.71fF $ **FLOATING
C1699 a_22081_13621# vssd1 0.72fF $ **FLOATING
C1700 a_21327_13866# vssd1 0.52fF $ **FLOATING
C1701 a_19899_13647# vssd1 0.97fF $ **FLOATING
C1702 _1191_.A1 vssd1 5.52fF $ **FLOATING
C1703 _1191_.B1 vssd1 1.59fF $ **FLOATING
C1704 a_19103_13985# vssd1 0.56fF $ **FLOATING
C1705 a_18243_13760# vssd1 0.62fF $ **FLOATING
C1706 a_17415_13760# vssd1 0.62fF $ **FLOATING
C1707 _1023_.B vssd1 6.34fF $ **FLOATING
C1708 a_15483_13760# vssd1 0.62fF $ **FLOATING
C1709 _1019_.B vssd1 7.32fF $ **FLOATING
C1710 _1050_.C vssd1 3.10fF $ **FLOATING
C1711 _1050_.B vssd1 4.02fF $ **FLOATING
C1712 _1755_.A vssd1 7.31fF $ **FLOATING
C1713 a_13599_13866# vssd1 0.52fF $ **FLOATING
C1714 a_12575_13647# vssd1 0.61fF $ **FLOATING
C1715 a_12743_13621# vssd1 0.82fF $ **FLOATING
C1716 a_12150_13647# vssd1 0.63fF $ **FLOATING
C1717 a_12318_13621# vssd1 0.58fF $ **FLOATING
C1718 a_11877_13653# vssd1 1.43fF $ **FLOATING
C1719 _1906_.D vssd1 1.74fF $ **FLOATING
C1720 a_11711_13653# vssd1 1.81fF $ **FLOATING
C1721 _1010_.A vssd1 16.38fF $ **FLOATING
C1722 a_9912_13763# vssd1 0.50fF $ **FLOATING
C1723 _1012_.B vssd1 2.96fF $ **FLOATING
C1724 _1175_.B2 vssd1 3.84fF $ **FLOATING
C1725 _1012_.Y vssd1 2.44fF $ **FLOATING
C1726 a_6610_13879# vssd1 0.60fF $ **FLOATING
C1727 _1246_.B1 vssd1 3.27fF $ **FLOATING
C1728 _1246_.B2 vssd1 8.48fF $ **FLOATING
C1729 _1246_.A3 vssd1 2.86fF $ **FLOATING
C1730 _1246_.A2 vssd1 4.17fF $ **FLOATING
C1731 a_1641_13879# vssd1 0.72fF $ **FLOATING
C1732 a_26601_14191# vssd1 0.23fF $ **FLOATING
C1733 a_27111_14557# vssd1 0.61fF $ **FLOATING
C1734 a_27279_14459# vssd1 0.82fF $ **FLOATING
C1735 a_26686_14557# vssd1 0.63fF $ **FLOATING
C1736 a_26854_14303# vssd1 0.58fF $ **FLOATING
C1737 a_26413_14191# vssd1 1.43fF $ **FLOATING
C1738 a_26247_14191# vssd1 1.81fF $ **FLOATING
C1739 _1707_.X vssd1 1.82fF $ **FLOATING
C1740 _1984_.D vssd1 1.54fF $ **FLOATING
C1741 _1725_.X vssd1 1.72fF $ **FLOATING
C1742 _1153_.X vssd1 1.57fF $ **FLOATING
C1743 _1153_.A vssd1 13.04fF $ **FLOATING
C1744 _1136_.B vssd1 5.71fF $ **FLOATING
C1745 _1110_.X vssd1 3.01fF $ **FLOATING
C1746 _1110_.A vssd1 11.98fF $ **FLOATING
C1747 a_17812_14441# vssd1 0.26fF $ **FLOATING
C1748 a_16616_14441# vssd1 0.26fF $ **FLOATING
C1749 a_13304_14441# vssd1 0.26fF $ **FLOATING
C1750 _1038_.X vssd1 1.52fF $ **FLOATING
C1751 _1044_.X vssd1 2.21fF $ **FLOATING
C1752 _1558_.X vssd1 1.20fF $ **FLOATING
C1753 a_25283_14356# vssd1 0.52fF $ **FLOATING
C1754 _1722_.A vssd1 1.50fF $ **FLOATING
C1755 a_24639_14356# vssd1 0.52fF $ **FLOATING
C1756 a_23299_14557# vssd1 0.51fF $ **FLOATING
C1757 a_23119_14557# vssd1 0.60fF $ **FLOATING
C1758 a_22379_14557# vssd1 0.51fF $ **FLOATING
C1759 _1721_.B vssd1 7.95fF $ **FLOATING
C1760 a_22199_14557# vssd1 0.60fF $ **FLOATING
C1761 a_21279_14191# vssd1 0.62fF $ **FLOATING
C1762 a_20267_14191# vssd1 0.62fF $ **FLOATING
C1763 a_18519_14191# vssd1 0.62fF $ **FLOATING
C1764 _1033_.A2 vssd1 3.95fF $ **FLOATING
C1765 _1033_.A1 vssd1 6.99fF $ **FLOATING
C1766 _1033_.B1 vssd1 4.20fF $ **FLOATING
C1767 a_17381_14337# vssd1 0.67fF $ **FLOATING
C1768 _1099_.B1 vssd1 1.72fF $ **FLOATING
C1769 _1099_.D1 vssd1 2.08fF $ **FLOATING
C1770 a_16185_14337# vssd1 0.67fF $ **FLOATING
C1771 a_15387_14557# vssd1 0.51fF $ **FLOATING
C1772 a_15207_14557# vssd1 0.60fF $ **FLOATING
C1773 a_14467_14557# vssd1 0.51fF $ **FLOATING
C1774 _1440_.B vssd1 5.64fF $ **FLOATING
C1775 a_14287_14557# vssd1 0.60fF $ **FLOATING
C1776 _1038_.A1 vssd1 4.03fF $ **FLOATING
C1777 _1038_.C1 vssd1 3.25fF $ **FLOATING
C1778 _1038_.D1 vssd1 3.48fF $ **FLOATING
C1779 a_12873_14337# vssd1 0.67fF $ **FLOATING
C1780 _1263_.A vssd1 8.92fF $ **FLOATING
C1781 a_11159_14191# vssd1 0.62fF $ **FLOATING
C1782 a_10188_14441# vssd1 0.50fF $ **FLOATING
C1783 a_9167_14219# vssd1 0.56fF $ **FLOATING
C1784 a_8307_14191# vssd1 0.65fF $ **FLOATING
C1785 a_7571_14191# vssd1 0.65fF $ **FLOATING
C1786 a_6463_14441# vssd1 0.25fF $ **FLOATING
C1787 _1810_.X vssd1 2.98fF $ **FLOATING
C1788 a_5177_14441# vssd1 0.20fF $ **FLOATING
C1789 a_4173_14441# vssd1 0.19fF $ **FLOATING
C1790 a_1955_14441# vssd1 0.25fF $ **FLOATING
C1791 _1810_.A2 vssd1 3.44fF $ **FLOATING
C1792 a_6245_14165# vssd1 0.55fF $ **FLOATING
C1793 _1217_.B1 vssd1 2.98fF $ **FLOATING
C1794 _1217_.A2 vssd1 3.86fF $ **FLOATING
C1795 _1217_.A3 vssd1 5.56fF $ **FLOATING
C1796 a_5048_14165# vssd1 0.65fF $ **FLOATING
C1797 _1279_.A1 vssd1 6.52fF $ **FLOATING
C1798 a_4036_14165# vssd1 0.85fF $ **FLOATING
C1799 a_3063_14191# vssd1 0.62fF $ **FLOATING
C1800 _1223_.A2 vssd1 6.02fF $ **FLOATING
C1801 _1223_.B1 vssd1 1.35fF $ **FLOATING
C1802 a_1737_14165# vssd1 0.55fF $ **FLOATING
C1803 a_22238_14735# vssd1 0.33fF $ **FLOATING
C1804 a_20858_14735# vssd1 0.33fF $ **FLOATING
C1805 a_24301_14735# vssd1 0.23fF $ **FLOATING
C1806 _1190_.X vssd1 2.01fF $ **FLOATING
C1807 _1830_.Q vssd1 4.30fF $ **FLOATING
C1808 a_17352_14735# vssd1 0.26fF $ **FLOATING
C1809 a_19057_14735# vssd1 0.23fF $ **FLOATING
C1810 a_13948_14735# vssd1 0.26fF $ **FLOATING
C1811 _1104_.X vssd1 5.72fF $ **FLOATING
C1812 a_27807_14735# vssd1 0.51fF $ **FLOATING
C1813 a_27627_14735# vssd1 0.60fF $ **FLOATING
C1814 a_24811_14735# vssd1 0.61fF $ **FLOATING
C1815 a_24979_14709# vssd1 0.82fF $ **FLOATING
C1816 a_24386_14735# vssd1 0.63fF $ **FLOATING
C1817 a_24554_14709# vssd1 0.58fF $ **FLOATING
C1818 a_24113_14741# vssd1 1.43fF $ **FLOATING
C1819 _1979_.D vssd1 2.06fF $ **FLOATING
C1820 a_23947_14741# vssd1 1.81fF $ **FLOATING
C1821 a_23167_14954# vssd1 0.52fF $ **FLOATING
C1822 _1979_.Q vssd1 3.57fF $ **FLOATING
C1823 _1190_.B1 vssd1 2.74fF $ **FLOATING
C1824 a_22081_14709# vssd1 0.72fF $ **FLOATING
C1825 _0952_.A1 vssd1 17.20fF $ **FLOATING
C1826 _0952_.A2 vssd1 4.85fF $ **FLOATING
C1827 a_20701_14709# vssd1 0.72fF $ **FLOATING
C1828 a_19567_14735# vssd1 0.61fF $ **FLOATING
C1829 a_19735_14709# vssd1 0.82fF $ **FLOATING
C1830 a_19142_14735# vssd1 0.63fF $ **FLOATING
C1831 a_19310_14709# vssd1 0.58fF $ **FLOATING
C1832 a_18869_14741# vssd1 1.43fF $ **FLOATING
C1833 a_18703_14741# vssd1 1.81fF $ **FLOATING
C1834 _1830_.CLK vssd1 14.57fF $ **FLOATING
C1835 a_18107_14954# vssd1 0.52fF $ **FLOATING
C1836 _1091_.B1 vssd1 2.86fF $ **FLOATING
C1837 _1091_.C1 vssd1 2.37fF $ **FLOATING
C1838 a_16921_14709# vssd1 0.67fF $ **FLOATING
C1839 _1401_.A vssd1 1.08fF $ **FLOATING
C1840 a_16083_14954# vssd1 0.52fF $ **FLOATING
C1841 a_15115_14851# vssd1 0.70fF $ **FLOATING
C1842 _1091_.X vssd1 1.20fF $ **FLOATING
C1843 _1104_.C vssd1 1.21fF $ **FLOATING
C1844 _1104_.D vssd1 1.77fF $ **FLOATING
C1845 _1108_.X vssd1 1.87fF $ **FLOATING
C1846 a_10594_14735# vssd1 0.36fF $ **FLOATING
C1847 a_10397_14735# vssd1 0.25fF $ **FLOATING
C1848 a_10147_14735# vssd1 0.39fF $ **FLOATING
C1849 a_1965_14735# vssd1 0.19fF $ **FLOATING
C1850 a_8301_15055# vssd1 0.21fF $ **FLOATING
C1851 _1793_.Y vssd1 9.37fF $ **FLOATING
C1852 _1108_.A1 vssd1 2.82fF $ **FLOATING
C1853 _1108_.C1 vssd1 1.36fF $ **FLOATING
C1854 a_13517_14709# vssd1 0.67fF $ **FLOATING
C1855 _1441_.A vssd1 1.77fF $ **FLOATING
C1856 a_12587_14954# vssd1 0.52fF $ **FLOATING
C1857 a_11711_14848# vssd1 0.62fF $ **FLOATING
C1858 a_10814_14709# vssd1 0.65fF $ **FLOATING
C1859 a_9429_15033# vssd1 0.61fF $ **FLOATING
C1860 _1122_.A1 vssd1 6.61fF $ **FLOATING
C1861 a_9000_14967# vssd1 0.59fF $ **FLOATING
C1862 _1793_.A2 vssd1 2.56fF $ **FLOATING
C1863 a_8109_14796# vssd1 0.45fF $ **FLOATING
C1864 a_7201_14851# vssd1 0.60fF $ **FLOATING
C1865 _1218_.B vssd1 11.98fF $ **FLOATING
C1866 a_7101_14735# vssd1 0.49fF $ **FLOATING
C1867 a_5455_14735# vssd1 0.70fF $ **FLOATING
C1868 _0932_.A vssd1 2.31fF $ **FLOATING
C1869 a_2962_14735# vssd1 4.03fF $ **FLOATING
C1870 io_in[0] vssd1 7.82fF
C1871 _1247_.B1 vssd1 1.63fF $ **FLOATING
C1872 a_1828_14709# vssd1 0.85fF $ **FLOATING
C1873 a_27153_15279# vssd1 0.23fF $ **FLOATING
C1874 a_27663_15645# vssd1 0.61fF $ **FLOATING
C1875 a_27831_15547# vssd1 0.82fF $ **FLOATING
C1876 a_27238_15645# vssd1 0.63fF $ **FLOATING
C1877 a_27406_15391# vssd1 0.58fF $ **FLOATING
C1878 a_26965_15279# vssd1 1.43fF $ **FLOATING
C1879 a_26799_15279# vssd1 1.81fF $ **FLOATING
C1880 _1975_.Q vssd1 4.35fF $ **FLOATING
C1881 a_24945_15279# vssd1 0.23fF $ **FLOATING
C1882 a_25455_15645# vssd1 0.61fF $ **FLOATING
C1883 a_25623_15547# vssd1 0.82fF $ **FLOATING
C1884 a_25030_15645# vssd1 0.63fF $ **FLOATING
C1885 a_25198_15391# vssd1 0.58fF $ **FLOATING
C1886 a_24757_15279# vssd1 1.43fF $ **FLOATING
C1887 _1975_.D vssd1 2.70fF $ **FLOATING
C1888 a_24591_15279# vssd1 1.81fF $ **FLOATING
C1889 _1706_.X vssd1 2.13fF $ **FLOATING
C1890 _1046_.B vssd1 5.98fF $ **FLOATING
C1891 _1574_.X vssd1 1.55fF $ **FLOATING
C1892 _0951_.B vssd1 11.65fF $ **FLOATING
C1893 _1399_.X vssd1 2.48fF $ **FLOATING
C1894 a_14776_15529# vssd1 0.26fF $ **FLOATING
C1895 _1095_.X vssd1 1.59fF $ **FLOATING
C1896 _1846_.Q vssd1 3.57fF $ **FLOATING
C1897 a_12249_15279# vssd1 0.23fF $ **FLOATING
C1898 a_23671_15279# vssd1 0.70fF $ **FLOATING
C1899 a_22931_15645# vssd1 0.51fF $ **FLOATING
C1900 a_22751_15645# vssd1 0.60fF $ **FLOATING
C1901 a_21463_15279# vssd1 0.62fF $ **FLOATING
C1902 a_20267_15279# vssd1 0.62fF $ **FLOATING
C1903 a_19480_15529# vssd1 0.50fF $ **FLOATING
C1904 a_18427_15279# vssd1 0.62fF $ **FLOATING
C1905 a_17541_15307# vssd1 0.71fF $ **FLOATING
C1906 a_16711_15307# vssd1 0.56fF $ **FLOATING
C1907 a_15531_15444# vssd1 0.52fF $ **FLOATING
C1908 _1095_.B1 vssd1 3.09fF $ **FLOATING
C1909 _1095_.C1 vssd1 3.33fF $ **FLOATING
C1910 a_14345_15425# vssd1 0.67fF $ **FLOATING
C1911 a_12759_15645# vssd1 0.61fF $ **FLOATING
C1912 a_12927_15547# vssd1 0.82fF $ **FLOATING
C1913 a_12334_15645# vssd1 0.63fF $ **FLOATING
C1914 a_12502_15391# vssd1 0.58fF $ **FLOATING
C1915 a_12061_15279# vssd1 1.43fF $ **FLOATING
C1916 a_11895_15279# vssd1 1.81fF $ **FLOATING
C1917 _0987_.Y vssd1 10.35fF $ **FLOATING
C1918 a_11067_15529# vssd1 0.39fF $ **FLOATING
C1919 a_9889_15253# vssd1 0.61fF $ **FLOATING
C1920 _1199_.A1 vssd1 1.98fF $ **FLOATING
C1921 _1199_.X vssd1 7.60fF $ **FLOATING
C1922 a_8209_15529# vssd1 0.24fF $ **FLOATING
C1923 _1790_.Y vssd1 1.87fF $ **FLOATING
C1924 a_7649_15279# vssd1 0.23fF $ **FLOATING
C1925 a_4209_15279# vssd1 0.19fF $ **FLOATING
C1926 a_5829_15529# vssd1 0.19fF $ **FLOATING
C1927 _1278_.X vssd1 1.23fF $ **FLOATING
C1928 a_2778_15529# vssd1 0.22fF $ **FLOATING
C1929 a_9460_15431# vssd1 0.59fF $ **FLOATING
C1930 a_7472_15279# vssd1 0.50fF $ **FLOATING
C1931 a_7366_15279# vssd1 0.58fF $ **FLOATING
C1932 a_7189_15279# vssd1 0.50fF $ **FLOATING
C1933 _1316_.X vssd1 6.80fF $ **FLOATING
C1934 a_6870_15279# vssd1 0.54fF $ **FLOATING
C1935 _1316_.A vssd1 2.73fF $ **FLOATING
C1936 _1289_.B1 vssd1 7.68fF $ **FLOATING
C1937 a_5692_15253# vssd1 0.85fF $ **FLOATING
C1938 _1278_.A1 vssd1 1.28fF $ **FLOATING
C1939 a_4059_15431# vssd1 0.74fF $ **FLOATING
C1940 _1219_.A2 vssd1 9.20fF $ **FLOATING
C1941 _1219_.B1 vssd1 3.07fF $ **FLOATING
C1942 a_2472_15431# vssd1 0.70fF $ **FLOATING
C1943 a_1591_15279# vssd1 0.70fF $ **FLOATING
C1944 io_in[7] vssd1 1.41fF
C1945 _1974_.Q vssd1 6.35fF $ **FLOATING
C1946 a_24577_15823# vssd1 0.23fF $ **FLOATING
C1947 _1723_.X vssd1 1.38fF $ **FLOATING
C1948 a_21032_15823# vssd1 0.26fF $ **FLOATING
C1949 a_19836_15823# vssd1 0.26fF $ **FLOATING
C1950 a_17904_15823# vssd1 0.26fF $ **FLOATING
C1951 a_15931_15823# vssd1 0.35fF $ **FLOATING
C1952 a_15737_15823# vssd1 0.25fF $ **FLOATING
C1953 a_15483_15823# vssd1 0.38fF $ **FLOATING
C1954 _1034_.Y vssd1 6.15fF $ **FLOATING
C1955 _1097_.X vssd1 2.38fF $ **FLOATING
C1956 a_12637_15823# vssd1 0.19fF $ **FLOATING
C1957 _1071_.X vssd1 4.09fF $ **FLOATING
C1958 _0987_.B vssd1 3.54fF $ **FLOATING
C1959 _1705_.A vssd1 1.09fF $ **FLOATING
C1960 a_28043_16042# vssd1 0.52fF $ **FLOATING
C1961 a_27399_16042# vssd1 0.52fF $ **FLOATING
C1962 a_25087_15823# vssd1 0.61fF $ **FLOATING
C1963 a_25255_15797# vssd1 0.82fF $ **FLOATING
C1964 a_24662_15823# vssd1 0.63fF $ **FLOATING
C1965 a_24830_15797# vssd1 0.58fF $ **FLOATING
C1966 a_24389_15829# vssd1 1.43fF $ **FLOATING
C1967 _1701_.X vssd1 1.94fF $ **FLOATING
C1968 a_24223_15829# vssd1 1.81fF $ **FLOATING
C1969 a_23483_15823# vssd1 0.51fF $ **FLOATING
C1970 a_23303_15823# vssd1 0.60fF $ **FLOATING
C1971 a_22195_15823# vssd1 0.51fF $ **FLOATING
C1972 _1723_.B vssd1 5.80fF $ **FLOATING
C1973 a_22015_15823# vssd1 0.60fF $ **FLOATING
C1974 _1723_.A_N vssd1 12.18fF $ **FLOATING
C1975 _1081_.B1 vssd1 1.19fF $ **FLOATING
C1976 _1081_.C1 vssd1 1.92fF $ **FLOATING
C1977 _1081_.D1 vssd1 5.49fF $ **FLOATING
C1978 a_20601_15797# vssd1 0.67fF $ **FLOATING
C1979 _1130_.C1 vssd1 2.58fF $ **FLOATING
C1980 _1130_.D1 vssd1 3.27fF $ **FLOATING
C1981 a_19405_15797# vssd1 0.67fF $ **FLOATING
C1982 a_18611_15823# vssd1 0.70fF $ **FLOATING
C1983 _1029_.B1 vssd1 3.50fF $ **FLOATING
C1984 _1028_.X vssd1 1.31fF $ **FLOATING
C1985 a_17473_15797# vssd1 0.67fF $ **FLOATING
C1986 _1034_.D vssd1 1.84fF $ **FLOATING
C1987 _1029_.X vssd1 1.32fF $ **FLOATING
C1988 a_13551_15936# vssd1 0.62fF $ **FLOATING
C1989 _1071_.B1 vssd1 11.11fF $ **FLOATING
C1990 a_12500_15797# vssd1 0.85fF $ **FLOATING
C1991 a_11711_15831# vssd1 0.65fF $ **FLOATING
C1992 _1371_.A vssd1 4.34fF $ **FLOATING
C1993 a_11023_16042# vssd1 0.52fF $ **FLOATING
C1994 a_9963_15939# vssd1 0.86fF $ **FLOATING
C1995 _1314_.X vssd1 4.84fF $ **FLOATING
C1996 a_4897_15823# vssd1 0.24fF $ **FLOATING
C1997 a_1769_15823# vssd1 0.24fF $ **FLOATING
C1998 _1289_.A2 vssd1 2.15fF $ **FLOATING
C1999 a_8785_15974# vssd1 0.70fF $ **FLOATING
C2000 a_8307_15823# vssd1 0.79fF $ **FLOATING
C2001 a_8454_15797# vssd1 0.80fF $ **FLOATING
C2002 a_7387_15823# vssd1 0.99fF $ **FLOATING
C2003 a_6559_15936# vssd1 0.62fF $ **FLOATING
C2004 a_2686_15823# vssd1 4.03fF $ **FLOATING
C2005 clkbuf_1_1__f_io_in[0].A vssd1 6.74fF $ **FLOATING
C2006 _1298_.A1 vssd1 8.53fF $ **FLOATING
C2007 _1824_.Q vssd1 4.69fF $ **FLOATING
C2008 a_26969_16367# vssd1 0.23fF $ **FLOATING
C2009 a_27479_16733# vssd1 0.61fF $ **FLOATING
C2010 a_27647_16635# vssd1 0.82fF $ **FLOATING
C2011 a_27054_16733# vssd1 0.63fF $ **FLOATING
C2012 a_27222_16479# vssd1 0.58fF $ **FLOATING
C2013 a_26781_16367# vssd1 1.43fF $ **FLOATING
C2014 a_26615_16367# vssd1 1.81fF $ **FLOATING
C2015 a_25129_16367# vssd1 0.23fF $ **FLOATING
C2016 a_25639_16733# vssd1 0.61fF $ **FLOATING
C2017 a_25807_16635# vssd1 0.82fF $ **FLOATING
C2018 a_25214_16733# vssd1 0.63fF $ **FLOATING
C2019 a_25382_16479# vssd1 0.58fF $ **FLOATING
C2020 a_24941_16367# vssd1 1.43fF $ **FLOATING
C2021 _1985_.D vssd1 2.15fF $ **FLOATING
C2022 a_24775_16367# vssd1 1.81fF $ **FLOATING
C2023 _1985_.CLK vssd1 9.90fF $ **FLOATING
C2024 a_21042_16617# vssd1 0.33fF $ **FLOATING
C2025 _0939_.A vssd1 16.42fF $ **FLOATING
C2026 _1193_.X vssd1 4.69fF $ **FLOATING
C2027 a_16209_16617# vssd1 0.21fF $ **FLOATING
C2028 a_14641_16367# vssd1 0.23fF $ **FLOATING
C2029 a_23391_16733# vssd1 0.51fF $ **FLOATING
C2030 a_23211_16733# vssd1 0.60fF $ **FLOATING
C2031 a_22103_16733# vssd1 0.51fF $ **FLOATING
C2032 a_21923_16733# vssd1 0.60fF $ **FLOATING
C2033 _1985_.Q vssd1 4.09fF $ **FLOATING
C2034 a_20885_16341# vssd1 0.72fF $ **FLOATING
C2035 a_19471_16395# vssd1 0.56fF $ **FLOATING
C2036 a_17999_16395# vssd1 0.56fF $ **FLOATING
C2037 a_17171_16395# vssd1 0.56fF $ **FLOATING
C2038 a_16127_16617# vssd1 0.80fF $ **FLOATING
C2039 a_15151_16733# vssd1 0.61fF $ **FLOATING
C2040 a_15319_16635# vssd1 0.82fF $ **FLOATING
C2041 a_14726_16733# vssd1 0.63fF $ **FLOATING
C2042 a_14894_16479# vssd1 0.58fF $ **FLOATING
C2043 a_14453_16367# vssd1 1.43fF $ **FLOATING
C2044 _1850_.D vssd1 2.19fF $ **FLOATING
C2045 a_14287_16367# vssd1 1.81fF $ **FLOATING
C2046 _1850_.CLK vssd1 19.45fF $ **FLOATING
C2047 _1035_.X vssd1 1.64fF $ **FLOATING
C2048 _0935_.X vssd1 17.95fF $ **FLOATING
C2049 a_13367_16367# vssd1 0.62fF $ **FLOATING
C2050 a_12557_16600# vssd1 0.70fF $ **FLOATING
C2051 a_12079_16367# vssd1 0.79fF $ **FLOATING
C2052 a_12226_16341# vssd1 0.80fF $ **FLOATING
C2053 a_11269_16600# vssd1 0.70fF $ **FLOATING
C2054 a_10791_16367# vssd1 0.79fF $ **FLOATING
C2055 a_10938_16341# vssd1 0.80fF $ **FLOATING
C2056 a_9613_16600# vssd1 0.70fF $ **FLOATING
C2057 a_9135_16367# vssd1 0.79fF $ **FLOATING
C2058 a_9282_16341# vssd1 0.80fF $ **FLOATING
C2059 a_8307_16367# vssd1 0.65fF $ **FLOATING
C2060 a_7657_16617# vssd1 0.24fF $ **FLOATING
C2061 a_6923_16617# vssd1 0.25fF $ **FLOATING
C2062 _1789_.X vssd1 6.39fF $ **FLOATING
C2063 a_5911_16617# vssd1 0.25fF $ **FLOATING
C2064 a_2047_16617# vssd1 0.25fF $ **FLOATING
C2065 _1789_.A1 vssd1 1.26fF $ **FLOATING
C2066 a_6705_16341# vssd1 0.55fF $ **FLOATING
C2067 _1265_.A2 vssd1 1.47fF $ **FLOATING
C2068 _1265_.A1 vssd1 4.33fF $ **FLOATING
C2069 a_5693_16341# vssd1 0.55fF $ **FLOATING
C2070 a_4899_16733# vssd1 0.51fF $ **FLOATING
C2071 a_4719_16733# vssd1 0.60fF $ **FLOATING
C2072 _1324_.A vssd1 7.02fF $ **FLOATING
C2073 a_2971_16367# vssd1 1.20fF $ **FLOATING
C2074 _0917_.A vssd1 8.59fF $ **FLOATING
C2075 a_1829_16341# vssd1 0.55fF $ **FLOATING
C2076 _1700_.X vssd1 1.38fF $ **FLOATING
C2077 _1389_.X vssd1 1.45fF $ **FLOATING
C2078 a_25589_16911# vssd1 0.23fF $ **FLOATING
C2079 a_23565_16911# vssd1 0.23fF $ **FLOATING
C2080 a_19973_16911# vssd1 0.21fF $ **FLOATING
C2081 a_19889_16911# vssd1 0.17fF $ **FLOATING
C2082 a_18685_16911# vssd1 0.21fF $ **FLOATING
C2083 a_18601_16911# vssd1 0.17fF $ **FLOATING
C2084 _1027_.X vssd1 1.19fF $ **FLOATING
C2085 _1101_.X vssd1 3.11fF $ **FLOATING
C2086 a_10279_16911# vssd1 0.59fF $ **FLOATING
C2087 a_9921_16911# vssd1 0.48fF $ **FLOATING
C2088 a_9503_16911# vssd1 0.66fF $ **FLOATING
C2089 a_6588_16911# vssd1 0.24fF $ **FLOATING
C2090 a_4932_16911# vssd1 0.24fF $ **FLOATING
C2091 a_3965_16911# vssd1 0.21fF $ **FLOATING
C2092 a_3881_16911# vssd1 0.17fF $ **FLOATING
C2093 a_2505_16911# vssd1 0.32fF $ **FLOATING
C2094 _1788_.X vssd1 1.67fF $ **FLOATING
C2095 a_28083_16911# vssd1 0.51fF $ **FLOATING
C2096 a_27903_16911# vssd1 0.60fF $ **FLOATING
C2097 _1389_.A vssd1 2.58fF $ **FLOATING
C2098 a_27215_17130# vssd1 0.52fF $ **FLOATING
C2099 a_26099_16911# vssd1 0.61fF $ **FLOATING
C2100 a_26267_16885# vssd1 0.82fF $ **FLOATING
C2101 a_25674_16911# vssd1 0.63fF $ **FLOATING
C2102 a_25842_16885# vssd1 0.58fF $ **FLOATING
C2103 a_25401_16917# vssd1 1.43fF $ **FLOATING
C2104 a_25235_16917# vssd1 1.81fF $ **FLOATING
C2105 a_24075_16911# vssd1 0.61fF $ **FLOATING
C2106 a_24243_16885# vssd1 0.82fF $ **FLOATING
C2107 a_23650_16911# vssd1 0.63fF $ **FLOATING
C2108 a_23818_16885# vssd1 0.58fF $ **FLOATING
C2109 a_23377_16917# vssd1 1.43fF $ **FLOATING
C2110 _1831_.D vssd1 4.98fF $ **FLOATING
C2111 a_23211_16917# vssd1 1.81fF $ **FLOATING
C2112 a_22195_16911# vssd1 0.51fF $ **FLOATING
C2113 _1390_.B vssd1 5.31fF $ **FLOATING
C2114 a_22015_16911# vssd1 0.60fF $ **FLOATING
C2115 a_21091_16911# vssd1 0.51fF $ **FLOATING
C2116 a_20911_16911# vssd1 0.60fF $ **FLOATING
C2117 a_19807_16911# vssd1 0.97fF $ **FLOATING
C2118 _0953_.C1 vssd1 1.84fF $ **FLOATING
C2119 a_18519_16911# vssd1 0.97fF $ **FLOATING
C2120 _1179_.B1 vssd1 5.41fF $ **FLOATING
C2121 _1179_.B2 vssd1 4.39fF $ **FLOATING
C2122 _1179_.C1 vssd1 1.78fF $ **FLOATING
C2123 a_17139_17024# vssd1 0.62fF $ **FLOATING
C2124 a_16083_17130# vssd1 0.52fF $ **FLOATING
C2125 _1381_.A vssd1 0.91fF $ **FLOATING
C2126 a_14979_17130# vssd1 0.52fF $ **FLOATING
C2127 a_14144_17027# vssd1 0.50fF $ **FLOATING
C2128 a_13275_17024# vssd1 0.62fF $ **FLOATING
C2129 a_12447_17024# vssd1 0.62fF $ **FLOATING
C2130 a_11711_16919# vssd1 0.65fF $ **FLOATING
C2131 a_10667_16885# vssd1 1.08fF $ **FLOATING
C2132 a_8624_17027# vssd1 0.50fF $ **FLOATING
C2133 a_7479_17277# vssd1 0.89fF $ **FLOATING
C2134 a_3799_16911# vssd1 0.97fF $ **FLOATING
C2135 _1291_.A1 vssd1 17.47fF $ **FLOATING
C2136 _1291_.B1 vssd1 2.01fF $ **FLOATING
C2137 _1291_.B2 vssd1 2.40fF $ **FLOATING
C2138 _1230_.A4 vssd1 2.94fF $ **FLOATING
C2139 _1249_.A2 vssd1 7.50fF $ **FLOATING
C2140 _1249_.A1 vssd1 4.56fF $ **FLOATING
C2141 _1230_.B1 vssd1 3.97fF $ **FLOATING
C2142 a_2287_16885# vssd1 0.53fF $ **FLOATING
C2143 _1277_.A vssd1 6.33fF $ **FLOATING
C2144 _1277_.B vssd1 6.41fF $ **FLOATING
C2145 a_26785_17455# vssd1 0.23fF $ **FLOATING
C2146 a_27295_17821# vssd1 0.61fF $ **FLOATING
C2147 a_27463_17723# vssd1 0.82fF $ **FLOATING
C2148 a_26870_17821# vssd1 0.63fF $ **FLOATING
C2149 a_27038_17567# vssd1 0.58fF $ **FLOATING
C2150 a_26597_17455# vssd1 1.43fF $ **FLOATING
C2151 a_26431_17455# vssd1 1.81fF $ **FLOATING
C2152 _1914_.Q vssd1 6.29fF $ **FLOATING
C2153 a_24945_17455# vssd1 0.23fF $ **FLOATING
C2154 a_25455_17821# vssd1 0.61fF $ **FLOATING
C2155 a_25623_17723# vssd1 0.82fF $ **FLOATING
C2156 a_25030_17821# vssd1 0.63fF $ **FLOATING
C2157 a_25198_17567# vssd1 0.58fF $ **FLOATING
C2158 a_24757_17455# vssd1 1.43fF $ **FLOATING
C2159 _1914_.D vssd1 4.96fF $ **FLOATING
C2160 a_24591_17455# vssd1 1.81fF $ **FLOATING
C2161 _1127_.X vssd1 1.67fF $ **FLOATING
C2162 _1127_.A vssd1 15.85fF $ **FLOATING
C2163 _1890_.Q vssd1 7.91fF $ **FLOATING
C2164 a_18272_17705# vssd1 0.26fF $ **FLOATING
C2165 _1049_.X vssd1 3.52fF $ **FLOATING
C2166 _1090_.X vssd1 1.95fF $ **FLOATING
C2167 _1090_.C vssd1 15.18fF $ **FLOATING
C2168 _1398_.X vssd1 1.52fF $ **FLOATING
C2169 _1047_.C vssd1 16.03fF $ **FLOATING
C2170 a_9674_17705# vssd1 0.36fF $ **FLOATING
C2171 a_9477_17705# vssd1 0.25fF $ **FLOATING
C2172 a_9227_17705# vssd1 0.39fF $ **FLOATING
C2173 a_3155_17455# vssd1 0.18fF $ **FLOATING
C2174 a_6553_17705# vssd1 0.24fF $ **FLOATING
C2175 a_23395_17455# vssd1 0.70fF $ **FLOATING
C2176 a_22659_17455# vssd1 0.70fF $ **FLOATING
C2177 _1391_.A vssd1 1.20fF $ **FLOATING
C2178 a_21695_17620# vssd1 0.52fF $ **FLOATING
C2179 a_20267_17455# vssd1 0.62fF $ **FLOATING
C2180 a_19480_17705# vssd1 0.50fF $ **FLOATING
C2181 _1049_.B1 vssd1 2.57fF $ **FLOATING
C2182 _1049_.C1 vssd1 2.13fF $ **FLOATING
C2183 a_17841_17601# vssd1 0.67fF $ **FLOATING
C2184 a_17047_17455# vssd1 0.70fF $ **FLOATING
C2185 a_16219_17455# vssd1 0.62fF $ **FLOATING
C2186 a_15479_17821# vssd1 0.51fF $ **FLOATING
C2187 a_15299_17821# vssd1 0.60fF $ **FLOATING
C2188 a_14287_17455# vssd1 0.62fF $ **FLOATING
C2189 a_13399_17483# vssd1 0.56fF $ **FLOATING
C2190 a_11693_17821# vssd1 0.85fF $ **FLOATING
C2191 a_11527_17821# vssd1 0.60fF $ **FLOATING
C2192 a_10731_17483# vssd1 0.56fF $ **FLOATING
C2193 a_9894_17429# vssd1 0.65fF $ **FLOATING
C2194 a_7295_17455# vssd1 0.91fF $ **FLOATING
C2195 a_7442_17429# vssd1 1.31fF $ **FLOATING
C2196 a_5455_17455# vssd1 0.65fF $ **FLOATING
C2197 a_2225_17705# vssd1 0.21fF $ **FLOATING
C2198 a_3983_17455# vssd1 0.99fF $ **FLOATING
C2199 _0916_.A vssd1 8.70fF $ **FLOATING
C2200 _1323_.A2 vssd1 3.06fF $ **FLOATING
C2201 a_2143_17705# vssd1 0.80fF $ **FLOATING
C2202 _1250_.A1 vssd1 4.67fF $ **FLOATING
C2203 _1250_.B2 vssd1 3.60fF $ **FLOATING
C2204 _1976_.Q vssd1 4.02fF $ **FLOATING
C2205 a_24761_17999# vssd1 0.23fF $ **FLOATING
C2206 _1527_.X vssd1 2.78fF $ **FLOATING
C2207 a_19057_17999# vssd1 0.23fF $ **FLOATING
C2208 _1820_.Q vssd1 4.68fF $ **FLOATING
C2209 a_17217_17999# vssd1 0.23fF $ **FLOATING
C2210 _1382_.X vssd1 1.21fF $ **FLOATING
C2211 _1143_.X vssd1 3.89fF $ **FLOATING
C2212 _1693_.A vssd1 1.69fF $ **FLOATING
C2213 a_26295_18218# vssd1 0.52fF $ **FLOATING
C2214 a_25271_17999# vssd1 0.61fF $ **FLOATING
C2215 a_25439_17973# vssd1 0.82fF $ **FLOATING
C2216 a_24846_17999# vssd1 0.63fF $ **FLOATING
C2217 a_25014_17973# vssd1 0.58fF $ **FLOATING
C2218 a_24573_18005# vssd1 1.43fF $ **FLOATING
C2219 _1976_.D vssd1 3.02fF $ **FLOATING
C2220 a_24407_18005# vssd1 1.81fF $ **FLOATING
C2221 a_23667_17999# vssd1 0.51fF $ **FLOATING
C2222 a_23487_17999# vssd1 0.60fF $ **FLOATING
C2223 _1500_.A vssd1 1.27fF $ **FLOATING
C2224 a_22707_18218# vssd1 0.52fF $ **FLOATING
C2225 _1527_.A vssd1 1.92fF $ **FLOATING
C2226 a_22063_18218# vssd1 0.52fF $ **FLOATING
C2227 a_20999_17999# vssd1 0.51fF $ **FLOATING
C2228 a_20819_17999# vssd1 0.60fF $ **FLOATING
C2229 a_19567_17999# vssd1 0.61fF $ **FLOATING
C2230 a_19735_17973# vssd1 0.82fF $ **FLOATING
C2231 a_19142_17999# vssd1 0.63fF $ **FLOATING
C2232 a_19310_17973# vssd1 0.58fF $ **FLOATING
C2233 a_18869_18005# vssd1 1.43fF $ **FLOATING
C2234 _1821_.D vssd1 3.01fF $ **FLOATING
C2235 a_18703_18005# vssd1 1.81fF $ **FLOATING
C2236 a_17727_17999# vssd1 0.61fF $ **FLOATING
C2237 a_17895_17973# vssd1 0.82fF $ **FLOATING
C2238 a_17302_17999# vssd1 0.63fF $ **FLOATING
C2239 a_17470_17973# vssd1 0.58fF $ **FLOATING
C2240 a_17029_18005# vssd1 1.43fF $ **FLOATING
C2241 a_16863_18005# vssd1 1.81fF $ **FLOATING
C2242 a_15616_18115# vssd1 0.50fF $ **FLOATING
C2243 _1821_.Q vssd1 4.78fF $ **FLOATING
C2244 a_14655_18115# vssd1 0.70fF $ **FLOATING
C2245 _1143_.A vssd1 3.39fF $ **FLOATING
C2246 a_8807_17999# vssd1 0.59fF $ **FLOATING
C2247 a_8449_17999# vssd1 0.48fF $ **FLOATING
C2248 a_8031_17999# vssd1 0.66fF $ **FLOATING
C2249 _1820_.D vssd1 3.59fF $ **FLOATING
C2250 a_5727_17999# vssd1 0.25fF $ **FLOATING
C2251 a_4517_17999# vssd1 0.21fF $ **FLOATING
C2252 a_4433_17999# vssd1 0.17fF $ **FLOATING
C2253 a_2861_17999# vssd1 0.21fF $ **FLOATING
C2254 a_2777_17999# vssd1 0.17fF $ **FLOATING
C2255 _1786_.X vssd1 6.52fF $ **FLOATING
C2256 a_13551_17999# vssd1 1.20fF $ **FLOATING
C2257 a_12189_18150# vssd1 0.70fF $ **FLOATING
C2258 a_11711_17999# vssd1 0.79fF $ **FLOATING
C2259 a_11858_17973# vssd1 0.80fF $ **FLOATING
C2260 a_11023_18218# vssd1 0.52fF $ **FLOATING
C2261 a_10188_18115# vssd1 0.50fF $ **FLOATING
C2262 a_9195_17973# vssd1 1.08fF $ **FLOATING
C2263 a_6927_17999# vssd1 0.99fF $ **FLOATING
C2264 _1786_.A1 vssd1 3.97fF $ **FLOATING
C2265 a_5509_17973# vssd1 0.55fF $ **FLOATING
C2266 a_4351_17999# vssd1 0.97fF $ **FLOATING
C2267 _1267_.A1 vssd1 13.60fF $ **FLOATING
C2268 _1267_.B1 vssd1 2.05fF $ **FLOATING
C2269 _1267_.B2 vssd1 1.77fF $ **FLOATING
C2270 a_2695_17999# vssd1 0.97fF $ **FLOATING
C2271 _1281_.A1 vssd1 8.68fF $ **FLOATING
C2272 _1281_.B1 vssd1 2.66fF $ **FLOATING
C2273 a_25773_18543# vssd1 0.23fF $ **FLOATING
C2274 a_26283_18909# vssd1 0.61fF $ **FLOATING
C2275 a_26451_18811# vssd1 0.82fF $ **FLOATING
C2276 a_25858_18909# vssd1 0.63fF $ **FLOATING
C2277 a_26026_18655# vssd1 0.58fF $ **FLOATING
C2278 a_25585_18543# vssd1 1.43fF $ **FLOATING
C2279 a_25419_18543# vssd1 1.81fF $ **FLOATING
C2280 _1971_.D vssd1 1.18fF $ **FLOATING
C2281 a_22645_18543# vssd1 0.23fF $ **FLOATING
C2282 _1695_.A vssd1 2.61fF $ **FLOATING
C2283 a_24639_18708# vssd1 0.52fF $ **FLOATING
C2284 a_23155_18909# vssd1 0.61fF $ **FLOATING
C2285 a_23323_18811# vssd1 0.82fF $ **FLOATING
C2286 a_22730_18909# vssd1 0.63fF $ **FLOATING
C2287 a_22898_18655# vssd1 0.58fF $ **FLOATING
C2288 a_22457_18543# vssd1 1.43fF $ **FLOATING
C2289 a_22291_18543# vssd1 1.81fF $ **FLOATING
C2290 _1151_.X vssd1 3.40fF $ **FLOATING
C2291 a_19928_18793# vssd1 0.26fF $ **FLOATING
C2292 _1138_.X vssd1 2.80fF $ **FLOATING
C2293 _1070_.X vssd1 3.66fF $ **FLOATING
C2294 a_17221_18793# vssd1 0.21fF $ **FLOATING
C2295 a_21463_18543# vssd1 0.62fF $ **FLOATING
C2296 _1138_.B1 vssd1 3.59fF $ **FLOATING
C2297 _1138_.C1 vssd1 2.82fF $ **FLOATING
C2298 a_19497_18689# vssd1 0.67fF $ **FLOATING
C2299 a_18560_18793# vssd1 0.50fF $ **FLOATING
C2300 a_17139_18793# vssd1 0.80fF $ **FLOATING
C2301 _1070_.A2 vssd1 6.55fF $ **FLOATING
C2302 a_16311_18543# vssd1 0.70fF $ **FLOATING
C2303 a_15299_18543# vssd1 0.65fF $ **FLOATING
C2304 _1082_.X vssd1 6.24fF $ **FLOATING
C2305 _1082_.D vssd1 4.38fF $ **FLOATING
C2306 _1094_.X vssd1 2.51fF $ **FLOATING
C2307 _1376_.X vssd1 1.29fF $ **FLOATING
C2308 _1442_.A vssd1 4.70fF $ **FLOATING
C2309 a_8027_18793# vssd1 0.25fF $ **FLOATING
C2310 a_5635_18793# vssd1 0.25fF $ **FLOATING
C2311 a_4533_18793# vssd1 0.20fF $ **FLOATING
C2312 a_3069_18793# vssd1 0.19fF $ **FLOATING
C2313 a_1781_18793# vssd1 0.19fF $ **FLOATING
C2314 a_14379_18793# vssd1 0.70fF $ **FLOATING
C2315 a_12907_18543# vssd1 0.62fF $ **FLOATING
C2316 a_11983_18909# vssd1 0.51fF $ **FLOATING
C2317 a_11803_18909# vssd1 0.60fF $ **FLOATING
C2318 a_10865_18909# vssd1 0.67fF $ **FLOATING
C2319 a_10699_18543# vssd1 0.64fF $ **FLOATING
C2320 a_9360_18793# vssd1 0.50fF $ **FLOATING
C2321 _1255_.A1 vssd1 12.34fF $ **FLOATING
C2322 a_7809_18517# vssd1 0.55fF $ **FLOATING
C2323 a_6835_18543# vssd1 0.99fF $ **FLOATING
C2324 a_5417_18517# vssd1 0.55fF $ **FLOATING
C2325 _1326_.A2 vssd1 1.59fF $ **FLOATING
C2326 _1326_.A3 vssd1 1.72fF $ **FLOATING
C2327 a_4404_18517# vssd1 0.65fF $ **FLOATING
C2328 _1300_.B1 vssd1 5.25fF $ **FLOATING
C2329 _1300_.A1 vssd1 1.26fF $ **FLOATING
C2330 _1300_.A2 vssd1 2.37fF $ **FLOATING
C2331 a_2932_18517# vssd1 0.85fF $ **FLOATING
C2332 a_1644_18517# vssd1 0.85fF $ **FLOATING
C2333 _1826_.Q vssd1 4.65fF $ **FLOATING
C2334 a_24393_19087# vssd1 0.23fF $ **FLOATING
C2335 _1032_.X vssd1 3.36fF $ **FLOATING
C2336 _1105_.X vssd1 4.31fF $ **FLOATING
C2337 a_16064_19087# vssd1 0.26fF $ **FLOATING
C2338 _1020_.X vssd1 1.98fF $ **FLOATING
C2339 _1031_.X vssd1 4.46fF $ **FLOATING
C2340 _1107_.X vssd1 2.47fF $ **FLOATING
C2341 a_9037_19087# vssd1 0.24fF $ **FLOATING
C2342 a_5817_19087# vssd1 0.24fF $ **FLOATING
C2343 a_5081_19087# vssd1 0.24fF $ **FLOATING
C2344 a_4161_19087# vssd1 0.24fF $ **FLOATING
C2345 a_10765_19407# vssd1 0.18fF $ **FLOATING
C2346 a_10515_19407# vssd1 0.22fF $ **FLOATING
C2347 _1280_.Y vssd1 2.35fF $ **FLOATING
C2348 a_1965_19087# vssd1 0.19fF $ **FLOATING
C2349 a_3249_19453# vssd1 0.19fF $ **FLOATING
C2350 a_24903_19087# vssd1 0.61fF $ **FLOATING
C2351 a_25071_19061# vssd1 0.82fF $ **FLOATING
C2352 a_24478_19087# vssd1 0.63fF $ **FLOATING
C2353 a_24646_19061# vssd1 0.58fF $ **FLOATING
C2354 a_24205_19093# vssd1 1.43fF $ **FLOATING
C2355 _1826_.D vssd1 2.58fF $ **FLOATING
C2356 a_24039_19093# vssd1 1.81fF $ **FLOATING
C2357 a_23115_19087# vssd1 0.51fF $ **FLOATING
C2358 _1696_.B vssd1 6.96fF $ **FLOATING
C2359 a_22935_19087# vssd1 0.60fF $ **FLOATING
C2360 a_22195_19087# vssd1 0.51fF $ **FLOATING
C2361 a_22015_19087# vssd1 0.60fF $ **FLOATING
C2362 a_20860_19203# vssd1 0.50fF $ **FLOATING
C2363 a_20079_19087# vssd1 0.51fF $ **FLOATING
C2364 a_19899_19087# vssd1 0.60fF $ **FLOATING
C2365 a_18887_19200# vssd1 0.62fF $ **FLOATING
C2366 a_18100_19203# vssd1 0.50fF $ **FLOATING
C2367 _1394_.A vssd1 6.77fF $ **FLOATING
C2368 a_17231_19200# vssd1 0.62fF $ **FLOATING
C2369 _1020_.A2 vssd1 5.52fF $ **FLOATING
C2370 _1020_.B1 vssd1 1.36fF $ **FLOATING
C2371 _1020_.D1 vssd1 2.72fF $ **FLOATING
C2372 a_15633_19061# vssd1 0.67fF $ **FLOATING
C2373 a_14747_19200# vssd1 0.62fF $ **FLOATING
C2374 a_13919_19200# vssd1 0.62fF $ **FLOATING
C2375 a_13091_19200# vssd1 0.62fF $ **FLOATING
C2376 a_12061_19087# vssd1 0.67fF $ **FLOATING
C2377 a_11895_19087# vssd1 0.64fF $ **FLOATING
C2378 a_9779_19087# vssd1 0.70fF $ **FLOATING
C2379 fanout28.A vssd1 22.84fF $ **FLOATING
C2380 _1234_.A1 vssd1 12.15fF $ **FLOATING
C2381 a_6927_19087# vssd1 1.20fF $ **FLOATING
C2382 _1301_.A1 vssd1 12.77fF $ **FLOATING
C2383 _1254_.A2 vssd1 2.01fF $ **FLOATING
C2384 _1254_.B1 vssd1 1.37fF $ **FLOATING
C2385 _1231_.B1 vssd1 11.47fF $ **FLOATING
C2386 _1231_.B2 vssd1 2.23fF $ **FLOATING
C2387 a_2966_19131# vssd1 0.54fF $ **FLOATING
C2388 a_2836_19319# vssd1 0.64fF $ **FLOATING
C2389 a_1828_19061# vssd1 0.85fF $ **FLOATING
C2390 _1967_.Q vssd1 6.33fF $ **FLOATING
C2391 a_27337_19631# vssd1 0.23fF $ **FLOATING
C2392 a_27847_19997# vssd1 0.61fF $ **FLOATING
C2393 a_28015_19899# vssd1 0.82fF $ **FLOATING
C2394 a_27422_19997# vssd1 0.63fF $ **FLOATING
C2395 a_27590_19743# vssd1 0.58fF $ **FLOATING
C2396 a_27149_19631# vssd1 1.43fF $ **FLOATING
C2397 _1967_.D vssd1 4.39fF $ **FLOATING
C2398 a_26983_19631# vssd1 1.81fF $ **FLOATING
C2399 _1387_.X vssd1 3.33fF $ **FLOATING
C2400 _1393_.X vssd1 1.61fF $ **FLOATING
C2401 _1528_.A vssd1 8.07fF $ **FLOATING
C2402 _1032_.C vssd1 13.79fF $ **FLOATING
C2403 _1387_.A vssd1 2.17fF $ **FLOATING
C2404 a_23903_19796# vssd1 0.52fF $ **FLOATING
C2405 _1385_.A vssd1 1.78fF $ **FLOATING
C2406 a_22983_19796# vssd1 0.52fF $ **FLOATING
C2407 _1689_.A vssd1 2.14fF $ **FLOATING
C2408 a_22339_19796# vssd1 0.52fF $ **FLOATING
C2409 _1393_.A vssd1 2.40fF $ **FLOATING
C2410 a_21695_19796# vssd1 0.52fF $ **FLOATING
C2411 a_20860_19881# vssd1 0.50fF $ **FLOATING
C2412 a_19619_19997# vssd1 0.51fF $ **FLOATING
C2413 _1403_.B vssd1 7.36fF $ **FLOATING
C2414 a_19439_19997# vssd1 0.60fF $ **FLOATING
C2415 a_18151_19631# vssd1 0.65fF $ **FLOATING
C2416 a_17444_19881# vssd1 0.26fF $ **FLOATING
C2417 _1024_.X vssd1 2.74fF $ **FLOATING
C2418 _0985_.X vssd1 6.22fF $ **FLOATING
C2419 _0985_.A vssd1 3.72fF $ **FLOATING
C2420 _1100_.X vssd1 4.23fF $ **FLOATING
C2421 _1024_.A2 vssd1 7.82fF $ **FLOATING
C2422 _1024_.D1 vssd1 3.50fF $ **FLOATING
C2423 a_17013_19777# vssd1 0.67fF $ **FLOATING
C2424 a_15575_19881# vssd1 0.70fF $ **FLOATING
C2425 a_14747_19631# vssd1 0.62fF $ **FLOATING
C2426 a_12815_19631# vssd1 0.65fF $ **FLOATING
C2427 _1141_.C vssd1 14.64fF $ **FLOATING
C2428 _1905_.Q vssd1 4.03fF $ **FLOATING
C2429 a_10317_19631# vssd1 0.23fF $ **FLOATING
C2430 a_11895_19631# vssd1 0.62fF $ **FLOATING
C2431 a_10827_19997# vssd1 0.61fF $ **FLOATING
C2432 a_10995_19899# vssd1 0.82fF $ **FLOATING
C2433 a_10402_19997# vssd1 0.63fF $ **FLOATING
C2434 a_10570_19743# vssd1 0.58fF $ **FLOATING
C2435 a_10129_19631# vssd1 1.43fF $ **FLOATING
C2436 a_9963_19631# vssd1 1.81fF $ **FLOATING
C2437 a_4903_19631# vssd1 0.18fF $ **FLOATING
C2438 a_7015_19881# vssd1 0.25fF $ **FLOATING
C2439 _1325_.X vssd1 1.88fF $ **FLOATING
C2440 a_5911_19881# vssd1 0.25fF $ **FLOATING
C2441 _1780_.X vssd1 7.37fF $ **FLOATING
C2442 a_2609_19881# vssd1 0.19fF $ **FLOATING
C2443 _1777_.X vssd1 6.68fF $ **FLOATING
C2444 a_9176_19881# vssd1 0.50fF $ **FLOATING
C2445 a_8027_19997# vssd1 0.51fF $ **FLOATING
C2446 a_7847_19997# vssd1 0.60fF $ **FLOATING
C2447 _1325_.A2 vssd1 11.87fF $ **FLOATING
C2448 _1325_.B1 vssd1 6.71fF $ **FLOATING
C2449 a_6797_19605# vssd1 0.55fF $ **FLOATING
C2450 _1780_.B1 vssd1 15.37fF $ **FLOATING
C2451 a_5693_19605# vssd1 0.55fF $ **FLOATING
C2452 _1234_.Y vssd1 2.51fF $ **FLOATING
C2453 _1234_.A2 vssd1 10.35fF $ **FLOATING
C2454 a_3983_19631# vssd1 1.20fF $ **FLOATING
C2455 _0929_.A vssd1 11.71fF $ **FLOATING
C2456 _1311_.B1 vssd1 4.06fF $ **FLOATING
C2457 _1311_.A1 vssd1 4.50fF $ **FLOATING
C2458 _1311_.A2 vssd1 2.49fF $ **FLOATING
C2459 a_2472_19605# vssd1 0.85fF $ **FLOATING
C2460 a_1823_19796# vssd1 0.52fF $ **FLOATING
C2461 _1970_.Q vssd1 5.28fF $ **FLOATING
C2462 a_25589_20175# vssd1 0.23fF $ **FLOATING
C2463 _1525_.X vssd1 2.94fF $ **FLOATING
C2464 _1822_.Q vssd1 5.22fF $ **FLOATING
C2465 a_19053_20175# vssd1 0.21fF $ **FLOATING
C2466 a_18969_20175# vssd1 0.17fF $ **FLOATING
C2467 a_22553_20175# vssd1 0.23fF $ **FLOATING
C2468 _0975_.X vssd1 2.44fF $ **FLOATING
C2469 _1187_.X vssd1 6.26fF $ **FLOATING
C2470 a_26099_20175# vssd1 0.61fF $ **FLOATING
C2471 a_26267_20149# vssd1 0.82fF $ **FLOATING
C2472 a_25674_20175# vssd1 0.63fF $ **FLOATING
C2473 a_25842_20149# vssd1 0.58fF $ **FLOATING
C2474 a_25401_20181# vssd1 1.43fF $ **FLOATING
C2475 _1970_.D vssd1 1.92fF $ **FLOATING
C2476 a_25235_20181# vssd1 1.81fF $ **FLOATING
C2477 _1525_.A vssd1 1.80fF $ **FLOATING
C2478 a_24087_20394# vssd1 0.52fF $ **FLOATING
C2479 a_23063_20175# vssd1 0.61fF $ **FLOATING
C2480 a_23231_20149# vssd1 0.82fF $ **FLOATING
C2481 a_22638_20175# vssd1 0.63fF $ **FLOATING
C2482 a_22806_20149# vssd1 0.58fF $ **FLOATING
C2483 a_22365_20181# vssd1 1.43fF $ **FLOATING
C2484 _1822_.D vssd1 5.00fF $ **FLOATING
C2485 a_22199_20181# vssd1 1.81fF $ **FLOATING
C2486 _1521_.A vssd1 0.91fF $ **FLOATING
C2487 a_21327_20394# vssd1 0.52fF $ **FLOATING
C2488 a_20492_20291# vssd1 0.50fF $ **FLOATING
C2489 a_18887_20175# vssd1 0.97fF $ **FLOATING
C2490 _0975_.C1 vssd1 3.55fF $ **FLOATING
C2491 a_17723_20513# vssd1 0.56fF $ **FLOATING
C2492 a_16904_20291# vssd1 0.50fF $ **FLOATING
C2493 a_15299_20291# vssd1 0.70fF $ **FLOATING
C2494 _1187_.A vssd1 3.40fF $ **FLOATING
C2495 _0981_.B vssd1 12.99fF $ **FLOATING
C2496 _1781_.Y vssd1 9.20fF $ **FLOATING
C2497 a_13257_20495# vssd1 0.21fF $ **FLOATING
C2498 a_14043_20513# vssd1 0.56fF $ **FLOATING
C2499 a_13019_20495# vssd1 0.71fF $ **FLOATING
C2500 a_12027_20495# vssd1 0.71fF $ **FLOATING
C2501 a_11907_20175# vssd1 0.77fF $ **FLOATING
C2502 a_11711_20175# vssd1 0.74fF $ **FLOATING
C2503 a_10344_20495# vssd1 0.24fF $ **FLOATING
C2504 a_10154_20495# vssd1 0.22fF $ **FLOATING
C2505 _1233_.X vssd1 2.22fF $ **FLOATING
C2506 a_4525_20175# vssd1 0.21fF $ **FLOATING
C2507 _0956_.C vssd1 14.04fF $ **FLOATING
C2508 _1781_.B vssd1 4.71fF $ **FLOATING
C2509 _1313_.X vssd1 8.19fF $ **FLOATING
C2510 _1257_.X vssd1 1.72fF $ **FLOATING
C2511 a_3276_20495# vssd1 0.22fF $ **FLOATING
C2512 a_3185_20495# vssd1 0.12fF $ **FLOATING
C2513 _0930_.Y vssd1 4.82fF $ **FLOATING
C2514 a_9963_20175# vssd1 0.89fF $ **FLOATING
C2515 a_8785_20473# vssd1 0.61fF $ **FLOATING
C2516 _1233_.A1 vssd1 3.96fF $ **FLOATING
C2517 _1232_.Y vssd1 12.02fF $ **FLOATING
C2518 a_8356_20407# vssd1 0.59fF $ **FLOATING
C2519 a_7571_20175# vssd1 0.70fF $ **FLOATING
C2520 a_5455_20541# vssd1 0.73fF $ **FLOATING
C2521 a_4443_20175# vssd1 0.80fF $ **FLOATING
C2522 _1302_.B1 vssd1 2.08fF $ **FLOATING
C2523 a_3087_20175# vssd1 0.87fF $ **FLOATING
C2524 _1257_.B2 vssd1 3.25fF $ **FLOATING
C2525 _1257_.B1 vssd1 1.41fF $ **FLOATING
C2526 a_2327_20183# vssd1 0.65fF $ **FLOATING
C2527 _1313_.A vssd1 9.44fF $ **FLOATING
C2528 _0930_.A vssd1 20.49fF $ **FLOATING
C2529 _0930_.B vssd1 14.49fF $ **FLOATING
C2530 _1823_.Q vssd1 5.68fF $ **FLOATING
C2531 a_27153_20719# vssd1 0.23fF $ **FLOATING
C2532 a_27663_21085# vssd1 0.61fF $ **FLOATING
C2533 a_27831_20987# vssd1 0.82fF $ **FLOATING
C2534 a_27238_21085# vssd1 0.63fF $ **FLOATING
C2535 a_27406_20831# vssd1 0.58fF $ **FLOATING
C2536 a_26965_20719# vssd1 1.43fF $ **FLOATING
C2537 _1823_.D vssd1 2.87fF $ **FLOATING
C2538 a_26799_20719# vssd1 1.81fF $ **FLOATING
C2539 _1823_.CLK vssd1 12.44fF $ **FLOATING
C2540 _1973_.Q vssd1 6.74fF $ **FLOATING
C2541 a_24945_20719# vssd1 0.23fF $ **FLOATING
C2542 a_25455_21085# vssd1 0.61fF $ **FLOATING
C2543 a_25623_20987# vssd1 0.82fF $ **FLOATING
C2544 a_25030_21085# vssd1 0.63fF $ **FLOATING
C2545 a_25198_20831# vssd1 0.58fF $ **FLOATING
C2546 a_24757_20719# vssd1 1.43fF $ **FLOATING
C2547 a_24591_20719# vssd1 1.81fF $ **FLOATING
C2548 _1184_.X vssd1 2.80fF $ **FLOATING
C2549 a_19605_20969# vssd1 0.21fF $ **FLOATING
C2550 a_19521_20969# vssd1 0.17fF $ **FLOATING
C2551 _1137_.X vssd1 2.25fF $ **FLOATING
C2552 _1022_.X vssd1 1.21fF $ **FLOATING
C2553 _0963_.B vssd1 17.30fF $ **FLOATING
C2554 _1018_.X vssd1 2.25fF $ **FLOATING
C2555 a_10073_20693# vssd1 0.61fF $ **FLOATING
C2556 _1334_.A1 vssd1 3.86fF $ **FLOATING
C2557 a_6469_20719# vssd1 0.19fF $ **FLOATING
C2558 _1433_.X vssd1 4.55fF $ **FLOATING
C2559 _1557_.X vssd1 2.70fF $ **FLOATING
C2560 a_4253_20719# vssd1 0.17fF $ **FLOATING
C2561 a_6186_21041# vssd1 0.54fF $ **FLOATING
C2562 _1327_.A2_N vssd1 2.28fF $ **FLOATING
C2563 _1327_.A1_N vssd1 2.79fF $ **FLOATING
C2564 a_23023_21085# vssd1 0.51fF $ **FLOATING
C2565 a_22843_21085# vssd1 0.60fF $ **FLOATING
C2566 _1502_.A vssd1 2.10fF $ **FLOATING
C2567 a_22247_20884# vssd1 0.52fF $ **FLOATING
C2568 a_21412_20969# vssd1 0.50fF $ **FLOATING
C2569 a_20584_20969# vssd1 0.50fF $ **FLOATING
C2570 a_19439_20719# vssd1 0.97fF $ **FLOATING
C2571 _1184_.A2 vssd1 1.90fF $ **FLOATING
C2572 _1184_.B1 vssd1 6.13fF $ **FLOATING
C2573 _1184_.C1 vssd1 4.00fF $ **FLOATING
C2574 a_18519_20719# vssd1 0.62fF $ **FLOATING
C2575 a_17415_20719# vssd1 0.62fF $ **FLOATING
C2576 a_16159_20747# vssd1 0.56fF $ **FLOATING
C2577 a_15207_20719# vssd1 0.70fF $ **FLOATING
C2578 _1459_.A vssd1 24.67fF $ **FLOATING
C2579 a_14379_20719# vssd1 0.62fF $ **FLOATING
C2580 a_13183_20719# vssd1 0.70fF $ **FLOATING
C2581 a_12295_20747# vssd1 0.56fF $ **FLOATING
C2582 a_11476_20969# vssd1 0.50fF $ **FLOATING
C2583 _1443_.A vssd1 2.06fF $ **FLOATING
C2584 a_10839_20884# vssd1 0.52fF $ **FLOATING
C2585 a_9644_20871# vssd1 0.59fF $ **FLOATING
C2586 _1433_.A vssd1 2.55fF $ **FLOATING
C2587 a_8447_20884# vssd1 0.52fF $ **FLOATING
C2588 _1445_.A vssd1 1.76fF $ **FLOATING
C2589 a_7803_20884# vssd1 0.52fF $ **FLOATING
C2590 _1557_.A vssd1 1.46fF $ **FLOATING
C2591 a_7159_20884# vssd1 0.52fF $ **FLOATING
C2592 a_6056_20871# vssd1 0.64fF $ **FLOATING
C2593 a_5271_20719# vssd1 0.65fF $ **FLOATING
C2594 _1322_.A vssd1 4.45fF $ **FLOATING
C2595 a_2953_20969# vssd1 0.21fF $ **FLOATING
C2596 a_2869_20969# vssd1 0.17fF $ **FLOATING
C2597 a_1757_20969# vssd1 0.21fF $ **FLOATING
C2598 a_1673_20969# vssd1 0.17fF $ **FLOATING
C2599 a_4035_20693# vssd1 0.55fF $ **FLOATING
C2600 a_2787_20719# vssd1 0.97fF $ **FLOATING
C2601 _1269_.A1 vssd1 14.08fF $ **FLOATING
C2602 _1269_.B1 vssd1 2.58fF $ **FLOATING
C2603 _1268_.X vssd1 0.99fF $ **FLOATING
C2604 a_1591_20719# vssd1 0.97fF $ **FLOATING
C2605 _1283_.B1 vssd1 2.46fF $ **FLOATING
C2606 _1699_.X vssd1 1.25fF $ **FLOATING
C2607 _1969_.Q vssd1 5.00fF $ **FLOATING
C2608 a_24025_21263# vssd1 0.23fF $ **FLOATING
C2609 _1048_.X vssd1 2.45fF $ **FLOATING
C2610 a_15696_21263# vssd1 0.26fF $ **FLOATING
C2611 _1077_.X vssd1 2.05fF $ **FLOATING
C2612 _1851_.Q vssd1 6.40fF $ **FLOATING
C2613 a_11793_21263# vssd1 0.21fF $ **FLOATING
C2614 a_13721_21263# vssd1 0.23fF $ **FLOATING
C2615 _1072_.X vssd1 2.68fF $ **FLOATING
C2616 a_2009_21263# vssd1 0.67fF $ **FLOATING
C2617 _1699_.A vssd1 1.86fF $ **FLOATING
C2618 a_25559_21482# vssd1 0.52fF $ **FLOATING
C2619 a_24535_21263# vssd1 0.61fF $ **FLOATING
C2620 a_24703_21237# vssd1 0.82fF $ **FLOATING
C2621 a_24110_21263# vssd1 0.63fF $ **FLOATING
C2622 a_24278_21237# vssd1 0.58fF $ **FLOATING
C2623 a_23837_21269# vssd1 1.43fF $ **FLOATING
C2624 a_23671_21269# vssd1 1.81fF $ **FLOATING
C2625 _1515_.A vssd1 1.49fF $ **FLOATING
C2626 a_22983_21482# vssd1 0.52fF $ **FLOATING
C2627 a_22195_21263# vssd1 0.51fF $ **FLOATING
C2628 a_22015_21263# vssd1 0.60fF $ **FLOATING
C2629 _1690_.A_N vssd1 14.62fF $ **FLOATING
C2630 _1529_.A vssd1 1.37fF $ **FLOATING
C2631 a_21143_21482# vssd1 0.52fF $ **FLOATING
C2632 a_20308_21379# vssd1 0.50fF $ **FLOATING
C2633 a_19388_21379# vssd1 0.50fF $ **FLOATING
C2634 a_18519_21376# vssd1 0.62fF $ **FLOATING
C2635 a_17691_21376# vssd1 0.62fF $ **FLOATING
C2636 _1075_.C vssd1 13.48fF $ **FLOATING
C2637 a_16863_21376# vssd1 0.62fF $ **FLOATING
C2638 _1074_.C vssd1 18.61fF $ **FLOATING
C2639 _1074_.X vssd1 1.29fF $ **FLOATING
C2640 _1075_.X vssd1 1.70fF $ **FLOATING
C2641 _1077_.D1 vssd1 3.47fF $ **FLOATING
C2642 a_15265_21237# vssd1 0.67fF $ **FLOATING
C2643 a_14231_21263# vssd1 0.61fF $ **FLOATING
C2644 a_14399_21237# vssd1 0.82fF $ **FLOATING
C2645 a_13806_21263# vssd1 0.63fF $ **FLOATING
C2646 a_13974_21237# vssd1 0.58fF $ **FLOATING
C2647 a_13533_21269# vssd1 1.43fF $ **FLOATING
C2648 _1851_.D vssd1 2.17fF $ **FLOATING
C2649 a_13367_21269# vssd1 1.81fF $ **FLOATING
C2650 _1549_.A vssd1 2.05fF $ **FLOATING
C2651 a_12771_21482# vssd1 0.52fF $ **FLOATING
C2652 a_11711_21263# vssd1 0.80fF $ **FLOATING
C2653 a_10883_21271# vssd1 0.65fF $ **FLOATING
C2654 a_10055_21376# vssd1 0.62fF $ **FLOATING
C2655 _1139_.C vssd1 15.83fF $ **FLOATING
C2656 a_9223_21263# vssd1 0.51fF $ **FLOATING
C2657 a_9043_21263# vssd1 0.60fF $ **FLOATING
C2658 _1776_.X vssd1 3.62fF $ **FLOATING
C2659 a_5183_21583# vssd1 0.21fF $ **FLOATING
C2660 a_4064_21583# vssd1 0.15fF $ **FLOATING
C2661 io_out[5] vssd1 4.70fF
C2662 a_2706_21583# vssd1 0.26fF $ **FLOATING
C2663 a_2199_21583# vssd1 0.19fF $ **FLOATING
C2664 a_2009_21583# vssd1 0.19fF $ **FLOATING
C2665 io_out[1] vssd1 1.95fF
C2666 a_7755_21263# vssd1 1.20fF $ **FLOATING
C2667 a_6968_21379# vssd1 0.50fF $ **FLOATING
C2668 _1292_.C1 vssd1 2.98fF $ **FLOATING
C2669 a_5047_21237# vssd1 0.79fF $ **FLOATING
C2670 _1312_.B1 vssd1 1.90fF $ **FLOATING
C2671 a_3759_21237# vssd1 0.72fF $ **FLOATING
C2672 _1260_.B1 vssd1 2.13fF $ **FLOATING
C2673 a_1643_21237# vssd1 1.57fF $ **FLOATING
C2674 _1878_.Q vssd1 9.07fF $ **FLOATING
C2675 a_27153_21807# vssd1 0.23fF $ **FLOATING
C2676 a_27663_22173# vssd1 0.61fF $ **FLOATING
C2677 a_27831_22075# vssd1 0.82fF $ **FLOATING
C2678 a_27238_22173# vssd1 0.63fF $ **FLOATING
C2679 a_27406_21919# vssd1 0.58fF $ **FLOATING
C2680 a_26965_21807# vssd1 1.43fF $ **FLOATING
C2681 _1878_.D vssd1 4.34fF $ **FLOATING
C2682 a_26799_21807# vssd1 1.81fF $ **FLOATING
C2683 _1877_.Q vssd1 7.40fF $ **FLOATING
C2684 a_25313_21807# vssd1 0.23fF $ **FLOATING
C2685 a_25823_22173# vssd1 0.61fF $ **FLOATING
C2686 a_25991_22075# vssd1 0.82fF $ **FLOATING
C2687 a_25398_22173# vssd1 0.63fF $ **FLOATING
C2688 a_25566_21919# vssd1 0.58fF $ **FLOATING
C2689 a_25125_21807# vssd1 1.43fF $ **FLOATING
C2690 a_24959_21807# vssd1 1.81fF $ **FLOATING
C2691 _1889_.Q vssd1 6.72fF $ **FLOATING
C2692 a_23013_21807# vssd1 0.23fF $ **FLOATING
C2693 a_23523_22173# vssd1 0.61fF $ **FLOATING
C2694 a_23691_22075# vssd1 0.82fF $ **FLOATING
C2695 a_23098_22173# vssd1 0.63fF $ **FLOATING
C2696 a_23266_21919# vssd1 0.58fF $ **FLOATING
C2697 a_22825_21807# vssd1 1.43fF $ **FLOATING
C2698 a_22659_21807# vssd1 1.81fF $ **FLOATING
C2699 _1889_.D vssd1 1.92fF $ **FLOATING
C2700 _1877_.D vssd1 3.60fF $ **FLOATING
C2701 _1113_.C vssd1 17.09fF $ **FLOATING
C2702 _1073_.X vssd1 2.86fF $ **FLOATING
C2703 a_16301_22057# vssd1 0.21fF $ **FLOATING
C2704 a_21827_22173# vssd1 0.51fF $ **FLOATING
C2705 a_21647_22173# vssd1 0.60fF $ **FLOATING
C2706 a_20768_22057# vssd1 0.50fF $ **FLOATING
C2707 _1523_.A vssd1 1.12fF $ **FLOATING
C2708 a_20131_21972# vssd1 0.52fF $ **FLOATING
C2709 _1395_.A vssd1 2.32fF $ **FLOATING
C2710 a_19487_21972# vssd1 0.52fF $ **FLOATING
C2711 a_18751_21972# vssd1 0.52fF $ **FLOATING
C2712 _1397_.A vssd1 1.73fF $ **FLOATING
C2713 a_18107_21972# vssd1 0.52fF $ **FLOATING
C2714 a_17231_21807# vssd1 0.62fF $ **FLOATING
C2715 a_16219_22057# vssd1 0.80fF $ **FLOATING
C2716 _1073_.A2 vssd1 6.10fF $ **FLOATING
C2717 a_15299_21807# vssd1 0.70fF $ **FLOATING
C2718 a_14563_21807# vssd1 0.65fF $ **FLOATING
C2719 a_10951_22057# vssd1 0.50fF $ **FLOATING
C2720 a_10593_22057# vssd1 0.42fF $ **FLOATING
C2721 a_9135_21807# vssd1 0.73fF $ **FLOATING
C2722 a_8395_22057# vssd1 0.25fF $ **FLOATING
C2723 a_5545_22057# vssd1 0.20fF $ **FLOATING
C2724 _1785_.X vssd1 2.62fF $ **FLOATING
C2725 a_4526_22057# vssd1 0.22fF $ **FLOATING
C2726 io_out[4] vssd1 3.85fF
C2727 a_2769_22057# vssd1 0.21fF $ **FLOATING
C2728 a_2685_22057# vssd1 0.17fF $ **FLOATING
C2729 a_1841_22057# vssd1 0.20fF $ **FLOATING
C2730 io_out[0] vssd1 2.69fF
C2731 a_13183_21807# vssd1 0.62fF $ **FLOATING
C2732 a_12396_22057# vssd1 0.50fF $ **FLOATING
C2733 a_10423_21807# vssd1 1.45fF $ **FLOATING
C2734 a_9284_21781# vssd1 0.72fF $ **FLOATING
C2735 _1293_.A1 vssd1 23.77fF $ **FLOATING
C2736 a_8177_21781# vssd1 0.55fF $ **FLOATING
C2737 a_6847_22057# vssd1 0.64fF $ **FLOATING
C2738 a_5416_21781# vssd1 0.65fF $ **FLOATING
C2739 a_4220_21959# vssd1 0.70fF $ **FLOATING
C2740 a_2603_21807# vssd1 0.97fF $ **FLOATING
C2741 _1237_.B2 vssd1 2.52fF $ **FLOATING
C2742 a_1643_21781# vssd1 0.80fF $ **FLOATING
C2743 _1879_.Q vssd1 4.94fF $ **FLOATING
C2744 a_25589_22351# vssd1 0.23fF $ **FLOATING
C2745 _1828_.Q vssd1 5.44fF $ **FLOATING
C2746 a_23105_22351# vssd1 0.23fF $ **FLOATING
C2747 _1497_.X vssd1 0.98fF $ **FLOATING
C2748 _1021_.X vssd1 1.96fF $ **FLOATING
C2749 a_15512_22351# vssd1 0.26fF $ **FLOATING
C2750 _1116_.X vssd1 4.89fF $ **FLOATING
C2751 a_12752_22351# vssd1 0.26fF $ **FLOATING
C2752 _1142_.X vssd1 3.43fF $ **FLOATING
C2753 a_9949_22351# vssd1 0.23fF $ **FLOATING
C2754 a_3435_22671# vssd1 0.21fF $ **FLOATING
C2755 _1240_.X vssd1 1.43fF $ **FLOATING
C2756 a_26099_22351# vssd1 0.61fF $ **FLOATING
C2757 a_26267_22325# vssd1 0.82fF $ **FLOATING
C2758 a_25674_22351# vssd1 0.63fF $ **FLOATING
C2759 a_25842_22325# vssd1 0.58fF $ **FLOATING
C2760 a_25401_22357# vssd1 1.43fF $ **FLOATING
C2761 _1879_.D vssd1 2.87fF $ **FLOATING
C2762 a_25235_22357# vssd1 1.81fF $ **FLOATING
C2763 a_23615_22351# vssd1 0.61fF $ **FLOATING
C2764 a_23783_22325# vssd1 0.82fF $ **FLOATING
C2765 a_23190_22351# vssd1 0.63fF $ **FLOATING
C2766 a_23358_22325# vssd1 0.58fF $ **FLOATING
C2767 a_22917_22357# vssd1 1.43fF $ **FLOATING
C2768 _1828_.D vssd1 2.60fF $ **FLOATING
C2769 a_22751_22357# vssd1 1.81fF $ **FLOATING
C2770 _1509_.A vssd1 1.78fF $ **FLOATING
C2771 a_22063_22570# vssd1 0.52fF $ **FLOATING
C2772 _1404_.A vssd1 2.24fF $ **FLOATING
C2773 a_21051_22570# vssd1 0.52fF $ **FLOATING
C2774 a_20216_22467# vssd1 0.50fF $ **FLOATING
C2775 a_19388_22467# vssd1 0.50fF $ **FLOATING
C2776 a_18560_22467# vssd1 0.50fF $ **FLOATING
C2777 a_17691_22464# vssd1 0.62fF $ **FLOATING
C2778 _1021_.A vssd1 13.08fF $ **FLOATING
C2779 a_16904_22467# vssd1 0.50fF $ **FLOATING
C2780 _1116_.B1 vssd1 1.79fF $ **FLOATING
C2781 _1116_.C1 vssd1 1.21fF $ **FLOATING
C2782 _1116_.D1 vssd1 1.75fF $ **FLOATING
C2783 a_15081_22325# vssd1 0.67fF $ **FLOATING
C2784 a_13643_22464# vssd1 0.62fF $ **FLOATING
C2785 _1142_.B1 vssd1 2.03fF $ **FLOATING
C2786 _1142_.D1 vssd1 1.78fF $ **FLOATING
C2787 a_12321_22325# vssd1 0.67fF $ **FLOATING
C2788 a_10459_22351# vssd1 0.61fF $ **FLOATING
C2789 a_10627_22325# vssd1 0.82fF $ **FLOATING
C2790 a_10034_22351# vssd1 0.63fF $ **FLOATING
C2791 a_10202_22325# vssd1 0.58fF $ **FLOATING
C2792 a_9761_22357# vssd1 1.43fF $ **FLOATING
C2793 _1817_.D vssd1 3.78fF $ **FLOATING
C2794 a_9595_22357# vssd1 1.81fF $ **FLOATING
C2795 a_8855_22351# vssd1 0.51fF $ **FLOATING
C2796 a_8675_22351# vssd1 0.60fF $ **FLOATING
C2797 a_7935_22351# vssd1 0.51fF $ **FLOATING
C2798 a_7755_22351# vssd1 0.60fF $ **FLOATING
C2799 a_7015_22351# vssd1 0.51fF $ **FLOATING
C2800 a_6835_22351# vssd1 0.60fF $ **FLOATING
C2801 _1374_.A_N vssd1 22.80fF $ **FLOATING
C2802 a_5565_22649# vssd1 0.61fF $ **FLOATING
C2803 _1303_.A1 vssd1 1.96fF $ **FLOATING
C2804 a_5136_22583# vssd1 0.59fF $ **FLOATING
C2805 a_4351_22359# vssd1 0.65fF $ **FLOATING
C2806 _1240_.B1 vssd1 0.96fF $ **FLOATING
C2807 a_3299_22325# vssd1 0.79fF $ **FLOATING
C2808 a_1779_22453# vssd1 0.75fF $ **FLOATING
C2809 a_1673_22453# vssd1 0.45fF $ **FLOATING
C2810 _1968_.Q vssd1 6.82fF $ **FLOATING
C2811 a_26417_22895# vssd1 0.23fF $ **FLOATING
C2812 a_26927_23261# vssd1 0.61fF $ **FLOATING
C2813 a_27095_23163# vssd1 0.82fF $ **FLOATING
C2814 a_26502_23261# vssd1 0.63fF $ **FLOATING
C2815 a_26670_23007# vssd1 0.58fF $ **FLOATING
C2816 a_26229_22895# vssd1 1.43fF $ **FLOATING
C2817 _1968_.D vssd1 3.88fF $ **FLOATING
C2818 a_26063_22895# vssd1 1.81fF $ **FLOATING
C2819 _1829_.Q vssd1 6.65fF $ **FLOATING
C2820 a_20897_22895# vssd1 0.23fF $ **FLOATING
C2821 _1517_.A vssd1 3.22fF $ **FLOATING
C2822 a_24639_23060# vssd1 0.52fF $ **FLOATING
C2823 _1697_.A vssd1 2.28fF $ **FLOATING
C2824 a_23535_23060# vssd1 0.52fF $ **FLOATING
C2825 a_22751_22895# vssd1 0.70fF $ **FLOATING
C2826 a_21407_23261# vssd1 0.61fF $ **FLOATING
C2827 a_21575_23163# vssd1 0.82fF $ **FLOATING
C2828 a_20982_23261# vssd1 0.63fF $ **FLOATING
C2829 a_21150_23007# vssd1 0.58fF $ **FLOATING
C2830 a_20709_22895# vssd1 1.43fF $ **FLOATING
C2831 _1829_.D vssd1 2.57fF $ **FLOATING
C2832 a_20543_22895# vssd1 1.81fF $ **FLOATING
C2833 _0964_.A vssd1 15.41fF $ **FLOATING
C2834 _1054_.C vssd1 5.59fF $ **FLOATING
C2835 _1055_.C vssd1 2.89fF $ **FLOATING
C2836 _0961_.A vssd1 16.06fF $ **FLOATING
C2837 _1186_.X vssd1 2.78fF $ **FLOATING
C2838 a_12153_23145# vssd1 0.21fF $ **FLOATING
C2839 a_12069_23145# vssd1 0.17fF $ **FLOATING
C2840 a_10413_23145# vssd1 0.21fF $ **FLOATING
C2841 a_6369_22895# vssd1 0.17fF $ **FLOATING
C2842 a_5449_22895# vssd1 0.17fF $ **FLOATING
C2843 a_4263_22895# vssd1 0.21fF $ **FLOATING
C2844 a_9613_22869# vssd1 0.61fF $ **FLOATING
C2845 _1238_.X vssd1 2.41fF $ **FLOATING
C2846 a_7561_22941# vssd1 0.43fF $ **FLOATING
C2847 _1282_.X vssd1 3.42fF $ **FLOATING
C2848 _1307_.X vssd1 1.60fF $ **FLOATING
C2849 a_1769_23145# vssd1 0.24fF $ **FLOATING
C2850 _0925_.Y vssd1 1.84fF $ **FLOATING
C2851 a_19619_23261# vssd1 0.51fF $ **FLOATING
C2852 a_19439_23261# vssd1 0.60fF $ **FLOATING
C2853 a_18560_23145# vssd1 0.50fF $ **FLOATING
C2854 a_17539_22923# vssd1 0.56fF $ **FLOATING
C2855 a_16711_22923# vssd1 0.56fF $ **FLOATING
C2856 a_15851_22895# vssd1 0.62fF $ **FLOATING
C2857 _1545_.A vssd1 0.88fF $ **FLOATING
C2858 a_15255_23060# vssd1 0.52fF $ **FLOATING
C2859 a_14467_23261# vssd1 0.51fF $ **FLOATING
C2860 a_14287_23261# vssd1 0.60fF $ **FLOATING
C2861 _1544_.A_N vssd1 22.04fF $ **FLOATING
C2862 a_13367_22895# vssd1 0.62fF $ **FLOATING
C2863 a_11987_22895# vssd1 0.97fF $ **FLOATING
C2864 _1186_.C1 vssd1 1.05fF $ **FLOATING
C2865 a_11391_23060# vssd1 0.52fF $ **FLOATING
C2866 a_10331_23145# vssd1 0.80fF $ **FLOATING
C2867 _1817_.Q vssd1 3.14fF $ **FLOATING
C2868 a_9184_23047# vssd1 0.59fF $ **FLOATING
C2869 a_7667_22901# vssd1 0.67fF $ **FLOATING
C2870 _1282_.A2 vssd1 7.99fF $ **FLOATING
C2871 a_6151_22869# vssd1 0.55fF $ **FLOATING
C2872 _1303_.X vssd1 1.06fF $ **FLOATING
C2873 a_5231_22869# vssd1 0.55fF $ **FLOATING
C2874 _1284_.B1 vssd1 2.57fF $ **FLOATING
C2875 a_4127_22869# vssd1 0.79fF $ **FLOATING
C2876 a_2649_23047# vssd1 0.77fF $ **FLOATING
C2877 a_2471_22869# vssd1 0.83fF $ **FLOATING
C2878 _0925_.A2 vssd1 14.19fF $ **FLOATING
C2879 _1888_.Q vssd1 7.83fF $ **FLOATING
C2880 a_25589_23439# vssd1 0.23fF $ **FLOATING
C2881 a_23565_23439# vssd1 0.23fF $ **FLOATING
C2882 _1691_.X vssd1 2.34fF $ **FLOATING
C2883 _1140_.X vssd1 1.73fF $ **FLOATING
C2884 a_6651_23439# vssd1 0.39fF $ **FLOATING
C2885 a_5061_23439# vssd1 0.20fF $ **FLOATING
C2886 a_1841_23439# vssd1 0.20fF $ **FLOATING
C2887 a_26099_23439# vssd1 0.61fF $ **FLOATING
C2888 a_26267_23413# vssd1 0.82fF $ **FLOATING
C2889 a_25674_23439# vssd1 0.63fF $ **FLOATING
C2890 a_25842_23413# vssd1 0.58fF $ **FLOATING
C2891 a_25401_23445# vssd1 1.43fF $ **FLOATING
C2892 _1888_.D vssd1 3.82fF $ **FLOATING
C2893 a_25235_23445# vssd1 1.81fF $ **FLOATING
C2894 a_24075_23439# vssd1 0.61fF $ **FLOATING
C2895 a_24243_23413# vssd1 0.82fF $ **FLOATING
C2896 a_23650_23439# vssd1 0.63fF $ **FLOATING
C2897 a_23818_23413# vssd1 0.58fF $ **FLOATING
C2898 a_23377_23445# vssd1 1.43fF $ **FLOATING
C2899 _1892_.D vssd1 2.78fF $ **FLOATING
C2900 a_23211_23445# vssd1 1.81fF $ **FLOATING
C2901 _1691_.A vssd1 1.56fF $ **FLOATING
C2902 a_22155_23658# vssd1 0.52fF $ **FLOATING
C2903 _1406_.A vssd1 1.57fF $ **FLOATING
C2904 a_21143_23658# vssd1 0.52fF $ **FLOATING
C2905 _1410_.A vssd1 1.51fF $ **FLOATING
C2906 a_20499_23658# vssd1 0.52fF $ **FLOATING
C2907 a_19664_23555# vssd1 0.50fF $ **FLOATING
C2908 _1506_.B vssd1 9.53fF $ **FLOATING
C2909 a_18836_23555# vssd1 0.50fF $ **FLOATING
C2910 _1405_.B vssd1 12.65fF $ **FLOATING
C2911 _1418_.A vssd1 1.35fF $ **FLOATING
C2912 a_17647_23658# vssd1 0.52fF $ **FLOATING
C2913 a_16863_23439# vssd1 0.70fF $ **FLOATING
C2914 a_15483_23552# vssd1 0.62fF $ **FLOATING
C2915 a_14655_23552# vssd1 0.62fF $ **FLOATING
C2916 _1053_.A vssd1 12.29fF $ **FLOATING
C2917 _1421_.A vssd1 1.94fF $ **FLOATING
C2918 a_13875_23658# vssd1 0.52fF $ **FLOATING
C2919 a_13040_23555# vssd1 0.50fF $ **FLOATING
C2920 a_12189_23737# vssd1 0.61fF $ **FLOATING
C2921 a_11760_23671# vssd1 0.59fF $ **FLOATING
C2922 a_10791_23552# vssd1 0.62fF $ **FLOATING
C2923 _1140_.C vssd1 20.83fF $ **FLOATING
C2924 a_10073_23737# vssd1 0.61fF $ **FLOATING
C2925 _1335_.A1 vssd1 2.14fF $ **FLOATING
C2926 a_9644_23671# vssd1 0.59fF $ **FLOATING
C2927 a_8399_23492# vssd1 0.79fF $ **FLOATING
C2928 a_8548_23413# vssd1 1.17fF $ **FLOATING
C2929 a_7481_23555# vssd1 0.66fF $ **FLOATING
C2930 _0922_.Y vssd1 8.26fF $ **FLOATING
C2931 io_out[3] vssd1 2.69fF
C2932 io_out[2] vssd1 1.73fF
C2933 _1375_.A vssd1 2.45fF $ **FLOATING
C2934 a_5871_23658# vssd1 0.52fF $ **FLOATING
C2935 _1285_.B1 vssd1 1.39fF $ **FLOATING
C2936 a_4863_23413# vssd1 0.80fF $ **FLOATING
C2937 a_2686_23439# vssd1 4.03fF $ **FLOATING
C2938 _1272_.B1 vssd1 1.17fF $ **FLOATING
C2939 _1272_.A2 vssd1 2.40fF $ **FLOATING
C2940 a_1643_23413# vssd1 0.80fF $ **FLOATING
C2941 _1885_.Q vssd1 6.65fF $ **FLOATING
C2942 a_26785_23983# vssd1 0.23fF $ **FLOATING
C2943 a_27295_24349# vssd1 0.61fF $ **FLOATING
C2944 a_27463_24251# vssd1 0.82fF $ **FLOATING
C2945 a_26870_24349# vssd1 0.63fF $ **FLOATING
C2946 a_27038_24095# vssd1 0.58fF $ **FLOATING
C2947 a_26597_23983# vssd1 1.43fF $ **FLOATING
C2948 _1885_.D vssd1 3.35fF $ **FLOATING
C2949 a_26431_23983# vssd1 1.81fF $ **FLOATING
C2950 _1972_.Q vssd1 7.40fF $ **FLOATING
C2951 a_24945_23983# vssd1 0.23fF $ **FLOATING
C2952 a_25455_24349# vssd1 0.61fF $ **FLOATING
C2953 a_25623_24251# vssd1 0.82fF $ **FLOATING
C2954 a_25030_24349# vssd1 0.63fF $ **FLOATING
C2955 a_25198_24095# vssd1 0.58fF $ **FLOATING
C2956 a_24757_23983# vssd1 1.43fF $ **FLOATING
C2957 _1972_.D vssd1 1.71fF $ **FLOATING
C2958 a_24591_23983# vssd1 1.81fF $ **FLOATING
C2959 _1832_.Q vssd1 6.10fF $ **FLOATING
C2960 a_22645_23983# vssd1 0.23fF $ **FLOATING
C2961 a_23155_24349# vssd1 0.61fF $ **FLOATING
C2962 a_23323_24251# vssd1 0.82fF $ **FLOATING
C2963 a_22730_24349# vssd1 0.63fF $ **FLOATING
C2964 a_22898_24095# vssd1 0.58fF $ **FLOATING
C2965 a_22457_23983# vssd1 1.43fF $ **FLOATING
C2966 _1832_.D vssd1 2.00fF $ **FLOATING
C2967 a_22291_23983# vssd1 1.81fF $ **FLOATING
C2968 a_17996_24233# vssd1 0.26fF $ **FLOATING
C2969 _1134_.X vssd1 4.29fF $ **FLOATING
C2970 _1845_.Q vssd1 6.76fF $ **FLOATING
C2971 a_16021_23983# vssd1 0.23fF $ **FLOATING
C2972 a_21091_24349# vssd1 0.51fF $ **FLOATING
C2973 a_20911_24349# vssd1 0.60fF $ **FLOATING
C2974 a_20171_24349# vssd1 0.51fF $ **FLOATING
C2975 a_19991_24349# vssd1 0.60fF $ **FLOATING
C2976 _1408_.A vssd1 1.09fF $ **FLOATING
C2977 a_18751_24148# vssd1 0.52fF $ **FLOATING
C2978 _1134_.B1 vssd1 1.76fF $ **FLOATING
C2979 a_17565_24129# vssd1 0.67fF $ **FLOATING
C2980 a_16531_24349# vssd1 0.61fF $ **FLOATING
C2981 a_16699_24251# vssd1 0.82fF $ **FLOATING
C2982 a_16106_24349# vssd1 0.63fF $ **FLOATING
C2983 a_16274_24095# vssd1 0.58fF $ **FLOATING
C2984 a_15833_23983# vssd1 1.43fF $ **FLOATING
C2985 a_15667_23983# vssd1 1.81fF $ **FLOATING
C2986 a_14776_24233# vssd1 0.26fF $ **FLOATING
C2987 _1056_.X vssd1 9.84fF $ **FLOATING
C2988 _0984_.X vssd1 3.62fF $ **FLOATING
C2989 a_12337_24233# vssd1 0.21fF $ **FLOATING
C2990 a_12253_24233# vssd1 0.17fF $ **FLOATING
C2991 a_10951_24233# vssd1 0.50fF $ **FLOATING
C2992 a_10593_24233# vssd1 0.42fF $ **FLOATING
C2993 a_5392_23983# vssd1 0.22fF $ **FLOATING
C2994 a_5301_23983# vssd1 0.12fF $ **FLOATING
C2995 _1294_.X vssd1 2.16fF $ **FLOATING
C2996 _2008_.Q vssd1 11.59fF $ **FLOATING
C2997 a_2405_23983# vssd1 0.23fF $ **FLOATING
C2998 _1056_.B1 vssd1 0.98fF $ **FLOATING
C2999 _1056_.C1 vssd1 1.80fF $ **FLOATING
C3000 _1056_.D1 vssd1 1.43fF $ **FLOATING
C3001 a_14345_24129# vssd1 0.67fF $ **FLOATING
C3002 a_13408_24233# vssd1 0.50fF $ **FLOATING
C3003 a_12171_23983# vssd1 0.97fF $ **FLOATING
C3004 _0984_.A2 vssd1 2.90fF $ **FLOATING
C3005 _0984_.B1 vssd1 7.28fF $ **FLOATING
C3006 a_10423_23983# vssd1 1.45fF $ **FLOATING
C3007 a_9268_24233# vssd1 0.50fF $ **FLOATING
C3008 a_8215_23983# vssd1 0.70fF $ **FLOATING
C3009 _1448_.A vssd1 21.64fF $ **FLOATING
C3010 a_7428_24233# vssd1 0.50fF $ **FLOATING
C3011 a_6600_24233# vssd1 0.50fF $ **FLOATING
C3012 a_5203_24233# vssd1 0.87fF $ **FLOATING
C3013 _1294_.B2 vssd1 2.73fF $ **FLOATING
C3014 _1294_.B1 vssd1 1.77fF $ **FLOATING
C3015 _1772_.A0 vssd1 8.28fF $ **FLOATING
C3016 a_4213_24135# vssd1 0.77fF $ **FLOATING
C3017 a_4035_23957# vssd1 0.83fF $ **FLOATING
C3018 a_2915_24349# vssd1 0.61fF $ **FLOATING
C3019 a_3083_24251# vssd1 0.82fF $ **FLOATING
C3020 a_2490_24349# vssd1 0.63fF $ **FLOATING
C3021 a_2658_24095# vssd1 0.58fF $ **FLOATING
C3022 a_2217_23983# vssd1 1.43fF $ **FLOATING
C3023 a_2051_23983# vssd1 1.81fF $ **FLOATING
C3024 _1884_.Q vssd1 5.95fF $ **FLOATING
C3025 a_25589_24527# vssd1 0.23fF $ **FLOATING
C3026 _1834_.Q vssd1 7.18fF $ **FLOATING
C3027 a_22369_24527# vssd1 0.23fF $ **FLOATING
C3028 _1133_.X vssd1 0.81fF $ **FLOATING
C3029 a_15833_24527# vssd1 0.21fF $ **FLOATING
C3030 a_15749_24527# vssd1 0.17fF $ **FLOATING
C3031 _1181_.X vssd1 2.83fF $ **FLOATING
C3032 _1819_.Q vssd1 4.92fF $ **FLOATING
C3033 a_13813_24527# vssd1 0.23fF $ **FLOATING
C3034 a_10399_24527# vssd1 0.50fF $ **FLOATING
C3035 a_10041_24527# vssd1 0.42fF $ **FLOATING
C3036 _1310_.Y vssd1 2.78fF $ **FLOATING
C3037 a_5731_24847# vssd1 0.18fF $ **FLOATING
C3038 _2006_.Q vssd1 14.27fF $ **FLOATING
C3039 a_1591_24527# vssd1 0.39fF $ **FLOATING
C3040 a_2957_24527# vssd1 0.23fF $ **FLOATING
C3041 a_26099_24527# vssd1 0.61fF $ **FLOATING
C3042 a_26267_24501# vssd1 0.82fF $ **FLOATING
C3043 a_25674_24527# vssd1 0.63fF $ **FLOATING
C3044 a_25842_24501# vssd1 0.58fF $ **FLOATING
C3045 a_25401_24533# vssd1 1.43fF $ **FLOATING
C3046 a_25235_24533# vssd1 1.81fF $ **FLOATING
C3047 _1504_.A vssd1 2.93fF $ **FLOATING
C3048 a_24547_24746# vssd1 0.52fF $ **FLOATING
C3049 _1507_.A vssd1 2.92fF $ **FLOATING
C3050 a_23903_24746# vssd1 0.52fF $ **FLOATING
C3051 a_22879_24527# vssd1 0.61fF $ **FLOATING
C3052 a_23047_24501# vssd1 0.82fF $ **FLOATING
C3053 a_22454_24527# vssd1 0.63fF $ **FLOATING
C3054 a_22622_24501# vssd1 0.58fF $ **FLOATING
C3055 a_22181_24533# vssd1 1.43fF $ **FLOATING
C3056 _1834_.D vssd1 2.49fF $ **FLOATING
C3057 a_22015_24533# vssd1 1.81fF $ **FLOATING
C3058 _1519_.A vssd1 1.05fF $ **FLOATING
C3059 a_21051_24746# vssd1 0.52fF $ **FLOATING
C3060 _1414_.A vssd1 1.55fF $ **FLOATING
C3061 a_20407_24746# vssd1 0.52fF $ **FLOATING
C3062 a_19619_24527# vssd1 0.51fF $ **FLOATING
C3063 _1530_.B vssd1 6.00fF $ **FLOATING
C3064 a_19439_24527# vssd1 0.60fF $ **FLOATING
C3065 a_18423_24527# vssd1 0.51fF $ **FLOATING
C3066 a_18243_24527# vssd1 0.60fF $ **FLOATING
C3067 a_17415_24640# vssd1 0.62fF $ **FLOATING
C3068 _1133_.C vssd1 13.78fF $ **FLOATING
C3069 a_15667_24527# vssd1 0.97fF $ **FLOATING
C3070 a_14323_24527# vssd1 0.61fF $ **FLOATING
C3071 a_14491_24501# vssd1 0.82fF $ **FLOATING
C3072 a_13898_24527# vssd1 0.63fF $ **FLOATING
C3073 a_14066_24501# vssd1 0.58fF $ **FLOATING
C3074 a_13625_24533# vssd1 1.43fF $ **FLOATING
C3075 _1819_.D vssd1 4.76fF $ **FLOATING
C3076 a_13459_24533# vssd1 1.81fF $ **FLOATING
C3077 a_12189_24825# vssd1 0.61fF $ **FLOATING
C3078 a_11760_24759# vssd1 0.59fF $ **FLOATING
C3079 a_9871_24527# vssd1 1.45fF $ **FLOATING
C3080 _0918_.A vssd1 12.97fF $ **FLOATING
C3081 _1547_.A vssd1 3.22fF $ **FLOATING
C3082 a_9275_24746# vssd1 0.52fF $ **FLOATING
C3083 a_8440_24643# vssd1 0.50fF $ **FLOATING
C3084 a_7479_24527# vssd1 1.20fF $ **FLOATING
C3085 a_6559_24640# vssd1 0.62fF $ **FLOATING
C3086 _1304_.B vssd1 18.63fF $ **FLOATING
C3087 _1310_.B1 vssd1 5.37fF $ **FLOATING
C3088 _1766_.A0 vssd1 8.68fF $ **FLOATING
C3089 a_4765_24759# vssd1 0.77fF $ **FLOATING
C3090 a_4587_24501# vssd1 0.83fF $ **FLOATING
C3091 a_3467_24527# vssd1 0.61fF $ **FLOATING
C3092 a_3635_24501# vssd1 0.97fF $ **FLOATING
C3093 a_3042_24527# vssd1 0.63fF $ **FLOATING
C3094 a_3210_24501# vssd1 0.58fF $ **FLOATING
C3095 a_2769_24533# vssd1 1.43fF $ **FLOATING
C3096 a_2603_24533# vssd1 1.81fF $ **FLOATING
C3097 _1771_.B vssd1 1.65fF $ **FLOATING
C3098 _1882_.Q vssd1 7.10fF $ **FLOATING
C3099 a_26417_25071# vssd1 0.23fF $ **FLOATING
C3100 a_26927_25437# vssd1 0.61fF $ **FLOATING
C3101 a_27095_25339# vssd1 0.82fF $ **FLOATING
C3102 a_26502_25437# vssd1 0.63fF $ **FLOATING
C3103 a_26670_25183# vssd1 0.58fF $ **FLOATING
C3104 a_26229_25071# vssd1 1.43fF $ **FLOATING
C3105 _1882_.D vssd1 4.09fF $ **FLOATING
C3106 a_26063_25071# vssd1 1.81fF $ **FLOATING
C3107 _1882_.CLK vssd1 10.18fF $ **FLOATING
C3108 _1270_.Y vssd1 11.17fF $ **FLOATING
C3109 _1270_.A vssd1 18.62fF $ **FLOATING
C3110 _1412_.A vssd1 2.38fF $ **FLOATING
C3111 a_23351_25236# vssd1 0.52fF $ **FLOATING
C3112 a_22567_25071# vssd1 0.65fF $ **FLOATING
C3113 _0958_.B vssd1 17.92fF $ **FLOATING
C3114 _0958_.A vssd1 28.77fF $ **FLOATING
C3115 a_16665_25071# vssd1 0.23fF $ **FLOATING
C3116 _1132_.X vssd1 2.24fF $ **FLOATING
C3117 _1132_.C vssd1 11.73fF $ **FLOATING
C3118 _1132_.A vssd1 19.97fF $ **FLOATING
C3119 _1852_.Q vssd1 6.61fF $ **FLOATING
C3120 a_11789_25071# vssd1 0.23fF $ **FLOATING
C3121 a_21831_25071# vssd1 0.70fF $ **FLOATING
C3122 _1511_.A vssd1 2.11fF $ **FLOATING
C3123 a_21235_25236# vssd1 0.52fF $ **FLOATING
C3124 _1416_.A vssd1 1.64fF $ **FLOATING
C3125 a_20315_25236# vssd1 0.52fF $ **FLOATING
C3126 a_19480_25321# vssd1 0.50fF $ **FLOATING
C3127 a_18367_25099# vssd1 0.56fF $ **FLOATING
C3128 a_17548_25321# vssd1 0.50fF $ **FLOATING
C3129 a_16488_25071# vssd1 0.50fF $ **FLOATING
C3130 a_16382_25071# vssd1 0.58fF $ **FLOATING
C3131 a_16205_25071# vssd1 0.50fF $ **FLOATING
C3132 a_15886_25071# vssd1 0.54fF $ **FLOATING
C3133 fanout37.A vssd1 12.94fF $ **FLOATING
C3134 a_14839_25071# vssd1 0.62fF $ **FLOATING
C3135 a_13316_25321# vssd1 0.50fF $ **FLOATING
C3136 a_12299_25437# vssd1 0.61fF $ **FLOATING
C3137 a_12467_25339# vssd1 0.82fF $ **FLOATING
C3138 a_11874_25437# vssd1 0.63fF $ **FLOATING
C3139 a_12042_25183# vssd1 0.58fF $ **FLOATING
C3140 a_11601_25071# vssd1 1.43fF $ **FLOATING
C3141 _1852_.D vssd1 4.60fF $ **FLOATING
C3142 a_11435_25071# vssd1 1.81fF $ **FLOATING
C3143 a_10349_25045# vssd1 0.61fF $ **FLOATING
C3144 _0906_.X vssd1 1.25fF $ **FLOATING
C3145 a_9920_25223# vssd1 0.59fF $ **FLOATING
C3146 a_9135_25071# vssd1 0.70fF $ **FLOATING
C3147 a_8213_25335# vssd1 0.60fF $ **FLOATING
C3148 a_8113_25117# vssd1 0.49fF $ **FLOATING
C3149 a_6230_25321# vssd1 0.33fF $ **FLOATING
C3150 _2007_.Q vssd1 6.33fF $ **FLOATING
C3151 a_4337_25071# vssd1 0.23fF $ **FLOATING
C3152 a_7111_25071# vssd1 1.20fF $ **FLOATING
C3153 a_6073_25045# vssd1 0.72fF $ **FLOATING
C3154 a_4847_25437# vssd1 0.61fF $ **FLOATING
C3155 a_5015_25339# vssd1 0.82fF $ **FLOATING
C3156 a_4422_25437# vssd1 0.63fF $ **FLOATING
C3157 a_4590_25183# vssd1 0.58fF $ **FLOATING
C3158 a_4149_25071# vssd1 1.43fF $ **FLOATING
C3159 _2007_.D vssd1 2.09fF $ **FLOATING
C3160 a_3983_25071# vssd1 1.81fF $ **FLOATING
C3161 _2005_.Q vssd1 16.17fF $ **FLOATING
C3162 a_2313_25071# vssd1 0.23fF $ **FLOATING
C3163 a_2823_25437# vssd1 0.61fF $ **FLOATING
C3164 a_2991_25339# vssd1 0.97fF $ **FLOATING
C3165 a_2398_25437# vssd1 0.63fF $ **FLOATING
C3166 a_2566_25183# vssd1 0.58fF $ **FLOATING
C3167 a_2125_25071# vssd1 1.43fF $ **FLOATING
C3168 a_1959_25071# vssd1 1.81fF $ **FLOATING
C3169 _1837_.Q vssd1 6.62fF $ **FLOATING
C3170 a_24209_25615# vssd1 0.23fF $ **FLOATING
C3171 _1833_.Q vssd1 7.46fF $ **FLOATING
C3172 a_22369_25615# vssd1 0.23fF $ **FLOATING
C3173 _1513_.X vssd1 3.08fF $ **FLOATING
C3174 _1900_.Q vssd1 7.55fF $ **FLOATING
C3175 a_15285_25615# vssd1 0.23fF $ **FLOATING
C3176 _1431_.X vssd1 2.11fF $ **FLOATING
C3177 _1901_.Q vssd1 4.80fF $ **FLOATING
C3178 a_12801_25615# vssd1 0.23fF $ **FLOATING
C3179 a_5639_25615# vssd1 0.39fF $ **FLOATING
C3180 a_2408_25615# vssd1 0.43fF $ **FLOATING
C3181 a_2153_25615# vssd1 0.32fF $ **FLOATING
C3182 _0911_.A vssd1 16.77fF $ **FLOATING
C3183 a_7755_25615# vssd1 0.53fF $ **FLOATING
C3184 a_2601_25935# vssd1 0.27fF $ **FLOATING
C3185 a_25695_25615# vssd1 0.52fF $ **FLOATING
C3186 a_24719_25615# vssd1 0.61fF $ **FLOATING
C3187 a_24887_25589# vssd1 0.82fF $ **FLOATING
C3188 a_24294_25615# vssd1 0.63fF $ **FLOATING
C3189 a_24462_25589# vssd1 0.58fF $ **FLOATING
C3190 a_24021_25621# vssd1 1.43fF $ **FLOATING
C3191 _1837_.D vssd1 2.94fF $ **FLOATING
C3192 a_23855_25621# vssd1 1.81fF $ **FLOATING
C3193 a_22879_25615# vssd1 0.61fF $ **FLOATING
C3194 a_23047_25589# vssd1 0.82fF $ **FLOATING
C3195 a_22454_25615# vssd1 0.63fF $ **FLOATING
C3196 a_22622_25589# vssd1 0.58fF $ **FLOATING
C3197 a_22181_25621# vssd1 1.43fF $ **FLOATING
C3198 _1833_.D vssd1 2.14fF $ **FLOATING
C3199 a_22015_25621# vssd1 1.81fF $ **FLOATING
C3200 _1513_.A vssd1 2.35fF $ **FLOATING
C3201 a_21235_25834# vssd1 0.52fF $ **FLOATING
C3202 _1531_.A vssd1 1.30fF $ **FLOATING
C3203 a_20315_25834# vssd1 0.52fF $ **FLOATING
C3204 _1496_.A vssd1 0.90fF $ **FLOATING
C3205 a_19671_25834# vssd1 0.52fF $ **FLOATING
C3206 _1534_.A vssd1 1.45fF $ **FLOATING
C3207 a_19027_25834# vssd1 0.52fF $ **FLOATING
C3208 a_18239_25615# vssd1 0.51fF $ **FLOATING
C3209 a_18059_25615# vssd1 0.60fF $ **FLOATING
C3210 a_16904_25731# vssd1 0.50fF $ **FLOATING
C3211 a_15795_25615# vssd1 0.61fF $ **FLOATING
C3212 a_15963_25589# vssd1 0.82fF $ **FLOATING
C3213 a_15370_25615# vssd1 0.63fF $ **FLOATING
C3214 a_15538_25589# vssd1 0.58fF $ **FLOATING
C3215 a_15097_25621# vssd1 1.43fF $ **FLOATING
C3216 _1900_.D vssd1 3.73fF $ **FLOATING
C3217 a_14931_25621# vssd1 1.81fF $ **FLOATING
C3218 _1431_.A vssd1 2.02fF $ **FLOATING
C3219 a_14335_25834# vssd1 0.52fF $ **FLOATING
C3220 a_13311_25615# vssd1 0.61fF $ **FLOATING
C3221 a_13479_25589# vssd1 0.82fF $ **FLOATING
C3222 a_12886_25615# vssd1 0.63fF $ **FLOATING
C3223 a_13054_25589# vssd1 0.58fF $ **FLOATING
C3224 a_12613_25621# vssd1 1.43fF $ **FLOATING
C3225 _1901_.D vssd1 2.45fF $ **FLOATING
C3226 a_12447_25621# vssd1 1.81fF $ **FLOATING
C3227 a_11711_25615# vssd1 0.70fF $ **FLOATING
C3228 a_10740_25731# vssd1 0.50fF $ **FLOATING
C3229 a_9889_25913# vssd1 0.61fF $ **FLOATING
C3230 _1336_.A1 vssd1 1.93fF $ **FLOATING
C3231 a_9460_25847# vssd1 0.59fF $ **FLOATING
C3232 a_8615_25953# vssd1 0.56fF $ **FLOATING
C3233 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 9.69fF $ **FLOATING
C3234 a_6968_25731# vssd1 0.50fF $ **FLOATING
C3235 _1305_.B vssd1 9.14fF $ **FLOATING
C3236 a_3514_25615# vssd1 4.03fF $ **FLOATING
C3237 _1763_.A2 vssd1 7.55fF $ **FLOATING
C3238 _1887_.Q vssd1 10.58fF $ **FLOATING
C3239 a_27337_26159# vssd1 0.23fF $ **FLOATING
C3240 a_27847_26525# vssd1 0.61fF $ **FLOATING
C3241 a_28015_26427# vssd1 0.82fF $ **FLOATING
C3242 a_27422_26525# vssd1 0.63fF $ **FLOATING
C3243 a_27590_26271# vssd1 0.58fF $ **FLOATING
C3244 a_27149_26159# vssd1 1.43fF $ **FLOATING
C3245 _1887_.D vssd1 4.30fF $ **FLOATING
C3246 a_26983_26159# vssd1 1.81fF $ **FLOATING
C3247 _1887_.CLK vssd1 11.64fF $ **FLOATING
C3248 _1881_.Q vssd1 8.73fF $ **FLOATING
C3249 a_25497_26159# vssd1 0.23fF $ **FLOATING
C3250 a_26007_26525# vssd1 0.61fF $ **FLOATING
C3251 a_26175_26427# vssd1 0.82fF $ **FLOATING
C3252 a_25582_26525# vssd1 0.63fF $ **FLOATING
C3253 a_25750_26271# vssd1 0.58fF $ **FLOATING
C3254 a_25309_26159# vssd1 1.43fF $ **FLOATING
C3255 _1881_.D vssd1 2.10fF $ **FLOATING
C3256 a_25143_26159# vssd1 1.81fF $ **FLOATING
C3257 _1308_.Y vssd1 9.19fF $ **FLOATING
C3258 _0921_.Y vssd1 10.28fF $ **FLOATING
C3259 _1838_.Q vssd1 5.67fF $ **FLOATING
C3260 a_21633_26159# vssd1 0.23fF $ **FLOATING
C3261 _1308_.B vssd1 17.37fF $ **FLOATING
C3262 _0921_.A vssd1 22.62fF $ **FLOATING
C3263 _0921_.B vssd1 21.47fF $ **FLOATING
C3264 a_22143_26525# vssd1 0.61fF $ **FLOATING
C3265 a_22311_26427# vssd1 0.82fF $ **FLOATING
C3266 a_21718_26525# vssd1 0.63fF $ **FLOATING
C3267 a_21886_26271# vssd1 0.58fF $ **FLOATING
C3268 a_21445_26159# vssd1 1.43fF $ **FLOATING
C3269 _1838_.D vssd1 1.66fF $ **FLOATING
C3270 a_21279_26159# vssd1 1.81fF $ **FLOATING
C3271 _1898_.Q vssd1 6.36fF $ **FLOATING
C3272 a_19793_26159# vssd1 0.23fF $ **FLOATING
C3273 a_20303_26525# vssd1 0.61fF $ **FLOATING
C3274 a_20471_26427# vssd1 0.82fF $ **FLOATING
C3275 a_19878_26525# vssd1 0.63fF $ **FLOATING
C3276 a_20046_26271# vssd1 0.58fF $ **FLOATING
C3277 a_19605_26159# vssd1 1.43fF $ **FLOATING
C3278 a_19439_26159# vssd1 1.81fF $ **FLOATING
C3279 a_16849_26159# vssd1 0.23fF $ **FLOATING
C3280 a_18607_26525# vssd1 0.51fF $ **FLOATING
C3281 a_18427_26525# vssd1 0.60fF $ **FLOATING
C3282 a_17359_26525# vssd1 0.61fF $ **FLOATING
C3283 a_17527_26427# vssd1 0.82fF $ **FLOATING
C3284 a_16934_26525# vssd1 0.63fF $ **FLOATING
C3285 a_17102_26271# vssd1 0.58fF $ **FLOATING
C3286 a_16661_26159# vssd1 1.43fF $ **FLOATING
C3287 _1840_.D vssd1 3.11fF $ **FLOATING
C3288 a_16495_26159# vssd1 1.81fF $ **FLOATING
C3289 _0966_.X vssd1 3.28fF $ **FLOATING
C3290 a_15005_26409# vssd1 0.21fF $ **FLOATING
C3291 a_14921_26409# vssd1 0.17fF $ **FLOATING
C3292 _1422_.X vssd1 2.61fF $ **FLOATING
C3293 _1840_.Q vssd1 7.58fF $ **FLOATING
C3294 _1422_.B vssd1 17.14fF $ **FLOATING
C3295 _0983_.X vssd1 2.16fF $ **FLOATING
C3296 a_10229_26409# vssd1 0.21fF $ **FLOATING
C3297 a_6921_26159# vssd1 0.17fF $ **FLOATING
C3298 a_4441_26159# vssd1 0.27fF $ **FLOATING
C3299 _1306_.X vssd1 2.43fF $ **FLOATING
C3300 a_5271_26409# vssd1 0.39fF $ **FLOATING
C3301 a_4248_26409# vssd1 0.43fF $ **FLOATING
C3302 _1769_.Y vssd1 2.11fF $ **FLOATING
C3303 a_3993_26409# vssd1 0.32fF $ **FLOATING
C3304 a_14839_26159# vssd1 0.97fF $ **FLOATING
C3305 _0966_.A2 vssd1 3.00fF $ **FLOATING
C3306 _0966_.B1 vssd1 4.37fF $ **FLOATING
C3307 a_13275_26159# vssd1 0.53fF $ **FLOATING
C3308 a_12488_26409# vssd1 0.50fF $ **FLOATING
C3309 a_11619_26159# vssd1 0.53fF $ **FLOATING
C3310 a_10147_26409# vssd1 0.80fF $ **FLOATING
C3311 _0983_.A2 vssd1 7.33fF $ **FLOATING
C3312 _0983_.B1 vssd1 8.65fF $ **FLOATING
C3313 a_9135_26159# vssd1 0.53fF $ **FLOATING
C3314 a_8215_26159# vssd1 0.53fF $ **FLOATING
C3315 _1373_.A vssd1 2.28fF $ **FLOATING
C3316 a_7619_26324# vssd1 0.52fF $ **FLOATING
C3317 _1306_.A2 vssd1 11.91fF $ **FLOATING
C3318 a_6703_26133# vssd1 0.55fF $ **FLOATING
C3319 a_1766_26159# vssd1 4.03fF $ **FLOATING
C3320 clkbuf_1_1__f__0380_.A vssd1 6.31fF $ **FLOATING
C3321 temp1.capload\[14\].cap.Y vssd1 0.28fF $ **FLOATING
C3322 temp1.capload\[3\].cap.Y vssd1 0.28fF $ **FLOATING
C3323 _1883_.Q vssd1 6.90fF $ **FLOATING
C3324 a_25589_26703# vssd1 0.23fF $ **FLOATING
C3325 _0923_.Y vssd1 14.25fF $ **FLOATING
C3326 _1839_.Q vssd1 10.58fF $ **FLOATING
C3327 a_22369_26703# vssd1 0.23fF $ **FLOATING
C3328 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.LO vssd1 0.48fF $ **FLOATING
C3329 a_13183_26703# vssd1 0.53fF $ **FLOATING
C3330 a_12355_26703# vssd1 0.53fF $ **FLOATING
C3331 a_26099_26703# vssd1 0.61fF $ **FLOATING
C3332 a_26267_26677# vssd1 0.82fF $ **FLOATING
C3333 a_25674_26703# vssd1 0.63fF $ **FLOATING
C3334 a_25842_26677# vssd1 0.58fF $ **FLOATING
C3335 a_25401_26709# vssd1 1.43fF $ **FLOATING
C3336 _1883_.D vssd1 3.28fF $ **FLOATING
C3337 a_25235_26709# vssd1 1.81fF $ **FLOATING
C3338 _1341_.A vssd1 9.01fF $ **FLOATING
C3339 a_23903_26922# vssd1 0.52fF $ **FLOATING
C3340 a_22879_26703# vssd1 0.61fF $ **FLOATING
C3341 a_23047_26677# vssd1 0.82fF $ **FLOATING
C3342 a_22454_26703# vssd1 0.63fF $ **FLOATING
C3343 a_22622_26677# vssd1 0.58fF $ **FLOATING
C3344 a_22181_26709# vssd1 1.43fF $ **FLOATING
C3345 _1839_.D vssd1 4.27fF $ **FLOATING
C3346 a_22015_26709# vssd1 1.81fF $ **FLOATING
C3347 _1553_.A vssd1 8.46fF $ **FLOATING
C3348 a_20959_26922# vssd1 0.52fF $ **FLOATING
C3349 _1536_.A vssd1 1.29fF $ **FLOATING
C3350 a_20315_26922# vssd1 0.52fF $ **FLOATING
C3351 _1494_.A vssd1 2.04fF $ **FLOATING
C3352 a_19487_26922# vssd1 0.52fF $ **FLOATING
C3353 a_18699_26703# vssd1 0.51fF $ **FLOATING
C3354 a_18519_26703# vssd1 0.60fF $ **FLOATING
C3355 _1461_.A vssd1 3.26fF $ **FLOATING
C3356 a_17923_26922# vssd1 0.52fF $ **FLOATING
C3357 a_17088_26819# vssd1 0.50fF $ **FLOATING
C3358 a_15800_26819# vssd1 0.50fF $ **FLOATING
C3359 _1537_.B vssd1 23.81fF $ **FLOATING
C3360 a_14972_26819# vssd1 0.50fF $ **FLOATING
C3361 a_14144_26819# vssd1 0.50fF $ **FLOATING
C3362 a_7843_26703# vssd1 0.25fF $ **FLOATING
C3363 a_6559_26703# vssd1 0.44fF $ **FLOATING
C3364 a_5639_26703# vssd1 0.39fF $ **FLOATING
C3365 a_4811_26703# vssd1 0.39fF $ **FLOATING
C3366 a_1775_26703# vssd1 0.39fF $ **FLOATING
C3367 a_8951_26703# vssd1 0.53fF $ **FLOATING
C3368 _1261_.X vssd1 1.96fF $ **FLOATING
C3369 _1762_.Y vssd1 2.86fF $ **FLOATING
C3370 _1769_.B1 vssd1 1.55fF $ **FLOATING
C3371 _1773_.Y vssd1 2.11fF $ **FLOATING
C3372 _1458_.A vssd1 1.16fF $ **FLOATING
C3373 a_11023_26922# vssd1 0.52fF $ **FLOATING
C3374 a_10257_27001# vssd1 0.61fF $ **FLOATING
C3375 _1328_.A1 vssd1 5.15fF $ **FLOATING
C3376 _1328_.S vssd1 11.49fF $ **FLOATING
C3377 a_9828_26935# vssd1 0.59fF $ **FLOATING
C3378 temp1.dac.vdac_single.einvp_batch\[0\].pupd_56.HI vssd1 1.82fF $ **FLOATING
C3379 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 5.76fF $ **FLOATING
C3380 _1261_.A2 vssd1 2.78fF $ **FLOATING
C3381 _1261_.A1 vssd1 16.63fF $ **FLOATING
C3382 a_7625_26677# vssd1 0.55fF $ **FLOATING
C3383 _1286_.A1 vssd1 18.51fF $ **FLOATING
C3384 _1762_.A vssd1 18.53fF $ **FLOATING
C3385 _1768_.A vssd1 17.34fF $ **FLOATING
C3386 a_2686_26703# vssd1 4.03fF $ **FLOATING
C3387 _1773_.B vssd1 2.67fF $ **FLOATING
C3388 _1836_.Q vssd1 8.38fF $ **FLOATING
C3389 a_27337_27247# vssd1 0.23fF $ **FLOATING
C3390 a_27847_27613# vssd1 0.61fF $ **FLOATING
C3391 a_28015_27515# vssd1 0.82fF $ **FLOATING
C3392 a_27422_27613# vssd1 0.63fF $ **FLOATING
C3393 a_27590_27359# vssd1 0.58fF $ **FLOATING
C3394 a_27149_27247# vssd1 1.43fF $ **FLOATING
C3395 _1836_.D vssd1 3.22fF $ **FLOATING
C3396 a_26983_27247# vssd1 1.81fF $ **FLOATING
C3397 _1835_.Q vssd1 6.55fF $ **FLOATING
C3398 a_24945_27247# vssd1 0.23fF $ **FLOATING
C3399 a_25455_27613# vssd1 0.61fF $ **FLOATING
C3400 a_25623_27515# vssd1 0.82fF $ **FLOATING
C3401 a_25030_27613# vssd1 0.63fF $ **FLOATING
C3402 a_25198_27359# vssd1 0.58fF $ **FLOATING
C3403 a_24757_27247# vssd1 1.43fF $ **FLOATING
C3404 _1835_.D vssd1 4.39fF $ **FLOATING
C3405 a_24591_27247# vssd1 1.81fF $ **FLOATING
C3406 _1893_.Q vssd1 6.33fF $ **FLOATING
C3407 a_23013_27247# vssd1 0.23fF $ **FLOATING
C3408 a_23523_27613# vssd1 0.61fF $ **FLOATING
C3409 a_23691_27515# vssd1 0.82fF $ **FLOATING
C3410 a_23098_27613# vssd1 0.63fF $ **FLOATING
C3411 a_23266_27359# vssd1 0.58fF $ **FLOATING
C3412 a_22825_27247# vssd1 1.43fF $ **FLOATING
C3413 _1893_.D vssd1 2.69fF $ **FLOATING
C3414 a_22659_27247# vssd1 1.81fF $ **FLOATING
C3415 _1332_.Y vssd1 14.13fF $ **FLOATING
C3416 io_out[6] vssd1 11.01fF
C3417 a_21371_27247# vssd1 0.52fF $ **FLOATING
C3418 _1492_.A vssd1 1.89fF $ **FLOATING
C3419 a_20775_27412# vssd1 0.52fF $ **FLOATING
C3420 a_20131_27412# vssd1 0.52fF $ **FLOATING
C3421 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.HI vssd1 0.42fF $ **FLOATING
C3422 _1427_.A vssd1 1.53fF $ **FLOATING
C3423 _1542_.X vssd1 2.68fF $ **FLOATING
C3424 _1904_.Q vssd1 5.51fF $ **FLOATING
C3425 a_10777_27247# vssd1 0.23fF $ **FLOATING
C3426 a_18239_27613# vssd1 0.51fF $ **FLOATING
C3427 a_18059_27613# vssd1 0.60fF $ **FLOATING
C3428 a_17139_27247# vssd1 0.53fF $ **FLOATING
C3429 temp1.dac.vdac_single.einvp_batch\[0\].vref_55.LO vssd1 2.10fF $ **FLOATING
C3430 _1542_.A vssd1 3.11fF $ **FLOATING
C3431 a_16267_27412# vssd1 0.52fF $ **FLOATING
C3432 a_15391_27247# vssd1 0.53fF $ **FLOATING
C3433 a_14604_27497# vssd1 0.50fF $ **FLOATING
C3434 a_13183_27247# vssd1 0.53fF $ **FLOATING
C3435 a_12355_27247# vssd1 0.53fF $ **FLOATING
C3436 a_11287_27613# vssd1 0.61fF $ **FLOATING
C3437 a_11455_27515# vssd1 0.82fF $ **FLOATING
C3438 a_10862_27613# vssd1 0.63fF $ **FLOATING
C3439 a_11030_27359# vssd1 0.58fF $ **FLOATING
C3440 a_10589_27247# vssd1 1.43fF $ **FLOATING
C3441 a_10423_27247# vssd1 1.81fF $ **FLOATING
C3442 a_6099_27247# vssd1 0.28fF $ **FLOATING
C3443 a_8569_27247# vssd1 0.23fF $ **FLOATING
C3444 a_4441_27247# vssd1 0.27fF $ **FLOATING
C3445 a_4248_27497# vssd1 0.43fF $ **FLOATING
C3446 a_3993_27497# vssd1 0.32fF $ **FLOATING
C3447 _2003_.Q vssd1 6.22fF $ **FLOATING
C3448 a_2405_27247# vssd1 0.23fF $ **FLOATING
C3449 a_9595_27247# vssd1 0.53fF $ **FLOATING
C3450 a_8392_27247# vssd1 0.50fF $ **FLOATING
C3451 a_8286_27247# vssd1 0.58fF $ **FLOATING
C3452 a_8109_27247# vssd1 0.50fF $ **FLOATING
C3453 a_7790_27247# vssd1 0.54fF $ **FLOATING
C3454 _1346_.A vssd1 3.98fF $ **FLOATING
C3455 a_6927_27247# vssd1 0.53fF $ **FLOATING
C3456 a_5271_27247# vssd1 0.53fF $ **FLOATING
C3457 a_2915_27613# vssd1 0.61fF $ **FLOATING
C3458 a_3083_27515# vssd1 0.82fF $ **FLOATING
C3459 a_2490_27613# vssd1 0.63fF $ **FLOATING
C3460 a_2658_27359# vssd1 0.58fF $ **FLOATING
C3461 a_2217_27247# vssd1 1.43fF $ **FLOATING
C3462 _2003_.D vssd1 1.58fF $ **FLOATING
C3463 a_2051_27247# vssd1 1.81fF $ **FLOATING
C3464 _1761_.X vssd1 12.43fF $ **FLOATING
C3465 a_27167_27791# vssd1 0.52fF $ **FLOATING
C3466 _1287_.A vssd1 14.09fF $ **FLOATING
C3467 a_25467_28010# vssd1 0.52fF $ **FLOATING
C3468 _1551_.A vssd1 9.73fF $ **FLOATING
C3469 a_24823_28010# vssd1 0.52fF $ **FLOATING
C3470 temp1.capload\[7\].cap_52.HI vssd1 0.42fF $ **FLOATING
C3471 _1876_.Q vssd1 6.92fF $ **FLOATING
C3472 a_22645_27791# vssd1 0.23fF $ **FLOATING
C3473 _1875_.Q vssd1 6.15fF $ **FLOATING
C3474 a_18785_27791# vssd1 0.21fF $ **FLOATING
C3475 a_20437_27791# vssd1 0.23fF $ **FLOATING
C3476 _0965_.X vssd1 3.46fF $ **FLOATING
C3477 _1899_.Q vssd1 7.19fF $ **FLOATING
C3478 a_15013_27791# vssd1 0.21fF $ **FLOATING
C3479 a_17217_27791# vssd1 0.23fF $ **FLOATING
C3480 a_15943_27791# vssd1 0.53fF $ **FLOATING
C3481 _1180_.X vssd1 1.90fF $ **FLOATING
C3482 a_13261_27791# vssd1 0.23fF $ **FLOATING
C3483 _1818_.Q vssd1 4.18fF $ **FLOATING
C3484 a_8120_27791# vssd1 0.24fF $ **FLOATING
C3485 a_9949_27791# vssd1 0.23fF $ **FLOATING
C3486 a_8767_27791# vssd1 0.53fF $ **FLOATING
C3487 a_5455_27791# vssd1 0.44fF $ **FLOATING
C3488 _0913_.Y vssd1 14.73fF $ **FLOATING
C3489 a_4627_27791# vssd1 0.53fF $ **FLOATING
C3490 _2004_.Q vssd1 17.45fF $ **FLOATING
C3491 a_1683_27791# vssd1 0.39fF $ **FLOATING
C3492 a_2957_27791# vssd1 0.23fF $ **FLOATING
C3493 _1767_.Y vssd1 2.11fF $ **FLOATING
C3494 a_23155_27791# vssd1 0.61fF $ **FLOATING
C3495 a_23323_27765# vssd1 0.82fF $ **FLOATING
C3496 a_22730_27791# vssd1 0.63fF $ **FLOATING
C3497 a_22898_27765# vssd1 0.58fF $ **FLOATING
C3498 a_22457_27797# vssd1 1.43fF $ **FLOATING
C3499 _1876_.D vssd1 2.96fF $ **FLOATING
C3500 a_22291_27797# vssd1 1.81fF $ **FLOATING
C3501 _1876_.CLK vssd1 11.37fF $ **FLOATING
C3502 a_20947_27791# vssd1 0.61fF $ **FLOATING
C3503 a_21115_27765# vssd1 0.82fF $ **FLOATING
C3504 a_20522_27791# vssd1 0.63fF $ **FLOATING
C3505 a_20690_27765# vssd1 0.58fF $ **FLOATING
C3506 a_20249_27797# vssd1 1.43fF $ **FLOATING
C3507 _1875_.D vssd1 1.56fF $ **FLOATING
C3508 a_20083_27797# vssd1 1.81fF $ **FLOATING
C3509 a_18703_27791# vssd1 0.80fF $ **FLOATING
C3510 a_17727_27791# vssd1 0.61fF $ **FLOATING
C3511 a_17895_27765# vssd1 0.82fF $ **FLOATING
C3512 a_17302_27791# vssd1 0.63fF $ **FLOATING
C3513 a_17470_27765# vssd1 0.58fF $ **FLOATING
C3514 a_17029_27797# vssd1 1.43fF $ **FLOATING
C3515 _1899_.D vssd1 3.56fF $ **FLOATING
C3516 a_16863_27797# vssd1 1.81fF $ **FLOATING
C3517 a_14931_27791# vssd1 0.80fF $ **FLOATING
C3518 _0965_.A2 vssd1 7.51fF $ **FLOATING
C3519 _0965_.B1 vssd1 6.18fF $ **FLOATING
C3520 a_14144_27907# vssd1 0.50fF $ **FLOATING
C3521 a_13084_27791# vssd1 0.50fF $ **FLOATING
C3522 a_12978_27791# vssd1 0.58fF $ **FLOATING
C3523 a_12801_27791# vssd1 0.50fF $ **FLOATING
C3524 a_12482_27791# vssd1 0.54fF $ **FLOATING
C3525 a_11711_27791# vssd1 0.70fF $ **FLOATING
C3526 a_10459_27791# vssd1 0.61fF $ **FLOATING
C3527 a_10627_27765# vssd1 0.82fF $ **FLOATING
C3528 a_10034_27791# vssd1 0.63fF $ **FLOATING
C3529 a_10202_27765# vssd1 0.58fF $ **FLOATING
C3530 a_9761_27797# vssd1 1.43fF $ **FLOATING
C3531 _1818_.D vssd1 2.48fF $ **FLOATING
C3532 a_9595_27797# vssd1 1.81fF $ **FLOATING
C3533 a_7847_27791# vssd1 0.57fF $ **FLOATING
C3534 a_6923_27791# vssd1 0.51fF $ **FLOATING
C3535 a_6743_27791# vssd1 0.60fF $ **FLOATING
C3536 _0913_.A1 vssd1 21.73fF $ **FLOATING
C3537 a_3467_27791# vssd1 0.61fF $ **FLOATING
C3538 a_3635_27765# vssd1 0.97fF $ **FLOATING
C3539 a_3042_27791# vssd1 0.63fF $ **FLOATING
C3540 a_3210_27765# vssd1 0.58fF $ **FLOATING
C3541 a_2769_27797# vssd1 1.43fF $ **FLOATING
C3542 _2004_.D vssd1 1.71fF $ **FLOATING
C3543 a_2603_27797# vssd1 1.81fF $ **FLOATING
C3544 _1767_.B vssd1 3.38fF $ **FLOATING
C3545 _1886_.Q vssd1 8.59fF $ **FLOATING
C3546 a_27245_28335# vssd1 0.23fF $ **FLOATING
C3547 a_27755_28701# vssd1 0.61fF $ **FLOATING
C3548 a_27923_28603# vssd1 0.82fF $ **FLOATING
C3549 a_27330_28701# vssd1 0.63fF $ **FLOATING
C3550 a_27498_28447# vssd1 0.58fF $ **FLOATING
C3551 a_27057_28335# vssd1 1.43fF $ **FLOATING
C3552 _1886_.D vssd1 4.09fF $ **FLOATING
C3553 a_26891_28335# vssd1 1.81fF $ **FLOATING
C3554 _1894_.Q vssd1 9.20fF $ **FLOATING
C3555 a_24945_28335# vssd1 0.23fF $ **FLOATING
C3556 a_25455_28701# vssd1 0.61fF $ **FLOATING
C3557 a_25623_28603# vssd1 0.82fF $ **FLOATING
C3558 a_25030_28701# vssd1 0.63fF $ **FLOATING
C3559 a_25198_28447# vssd1 0.58fF $ **FLOATING
C3560 a_24757_28335# vssd1 1.43fF $ **FLOATING
C3561 _1894_.D vssd1 4.60fF $ **FLOATING
C3562 a_24591_28335# vssd1 1.81fF $ **FLOATING
C3563 temp1.capload\[5\].cap_50.HI vssd1 0.42fF $ **FLOATING
C3564 temp1.capload\[3\].cap_48.LO vssd1 3.44fF $ **FLOATING
C3565 temp1.capload\[3\].cap_48.HI vssd1 0.42fF $ **FLOATING
C3566 temp1.capload\[9\].cap_54.HI vssd1 0.42fF $ **FLOATING
C3567 _1844_.Q vssd1 7.51fF $ **FLOATING
C3568 a_19977_28335# vssd1 0.23fF $ **FLOATING
C3569 _1483_.A vssd1 4.29fF $ **FLOATING
C3570 a_21511_28500# vssd1 0.52fF $ **FLOATING
C3571 a_20487_28701# vssd1 0.61fF $ **FLOATING
C3572 a_20655_28603# vssd1 0.82fF $ **FLOATING
C3573 a_20062_28701# vssd1 0.63fF $ **FLOATING
C3574 a_20230_28447# vssd1 0.58fF $ **FLOATING
C3575 a_19789_28335# vssd1 1.43fF $ **FLOATING
C3576 a_19623_28335# vssd1 1.81fF $ **FLOATING
C3577 a_7479_28585# vssd1 0.44fF $ **FLOATING
C3578 _1764_.Y vssd1 1.37fF $ **FLOATING
C3579 a_3983_28585# vssd1 0.39fF $ **FLOATING
C3580 a_2129_28335# vssd1 0.23fF $ **FLOATING
C3581 a_18607_28701# vssd1 0.51fF $ **FLOATING
C3582 a_18427_28701# vssd1 0.60fF $ **FLOATING
C3583 a_15750_28335# vssd1 4.03fF $ **FLOATING
C3584 a_14927_28701# vssd1 0.51fF $ **FLOATING
C3585 a_14747_28701# vssd1 0.60fF $ **FLOATING
C3586 _1489_.A_N vssd1 17.08fF $ **FLOATING
C3587 a_13183_28335# vssd1 0.53fF $ **FLOATING
C3588 a_12355_28335# vssd1 0.53fF $ **FLOATING
C3589 a_11527_28335# vssd1 0.53fF $ **FLOATING
C3590 a_10699_28335# vssd1 0.53fF $ **FLOATING
C3591 a_9871_28335# vssd1 0.53fF $ **FLOATING
C3592 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 8.92fF $ **FLOATING
C3593 _1274_.A vssd1 9.07fF $ **FLOATING
C3594 _1273_.A1 vssd1 16.51fF $ **FLOATING
C3595 a_5354_28335# vssd1 4.03fF $ **FLOATING
C3596 _1764_.B vssd1 6.90fF $ **FLOATING
C3597 _1764_.A vssd1 17.47fF $ **FLOATING
C3598 a_2639_28701# vssd1 0.61fF $ **FLOATING
C3599 a_2807_28603# vssd1 0.82fF $ **FLOATING
C3600 a_2214_28701# vssd1 0.63fF $ **FLOATING
C3601 a_2382_28447# vssd1 0.58fF $ **FLOATING
C3602 a_1941_28335# vssd1 1.43fF $ **FLOATING
C3603 a_1775_28335# vssd1 1.81fF $ **FLOATING
C3604 _2009_.CLK vssd1 16.96fF $ **FLOATING
C3605 _1344_.Y vssd1 10.35fF $ **FLOATING
C3606 _1342_.Y vssd1 10.12fF $ **FLOATING
C3607 _1895_.Q vssd1 7.07fF $ **FLOATING
C3608 a_24301_28879# vssd1 0.23fF $ **FLOATING
C3609 a_27859_29098# vssd1 0.52fF $ **FLOATING
C3610 _1344_.B vssd1 13.16fF $ **FLOATING
C3611 a_24811_28879# vssd1 0.61fF $ **FLOATING
C3612 a_24979_28853# vssd1 0.82fF $ **FLOATING
C3613 a_24386_28879# vssd1 0.63fF $ **FLOATING
C3614 a_24554_28853# vssd1 0.58fF $ **FLOATING
C3615 a_24113_28885# vssd1 1.43fF $ **FLOATING
C3616 _1895_.D vssd1 3.42fF $ **FLOATING
C3617 a_23947_28885# vssd1 1.81fF $ **FLOATING
C3618 temp1.capload\[12\].cap_42.HI vssd1 0.42fF $ **FLOATING
C3619 temp1.capload\[2\].cap.Y vssd1 0.28fF $ **FLOATING
C3620 a_20437_28879# vssd1 0.23fF $ **FLOATING
C3621 _1863_.Q vssd1 7.91fF $ **FLOATING
C3622 a_17677_28879# vssd1 0.23fF $ **FLOATING
C3623 a_13183_28879# vssd1 0.53fF $ **FLOATING
C3624 a_12355_28879# vssd1 0.53fF $ **FLOATING
C3625 _1429_.X vssd1 4.57fF $ **FLOATING
C3626 _1453_.X vssd1 7.89fF $ **FLOATING
C3627 a_9043_28879# vssd1 0.53fF $ **FLOATING
C3628 a_8215_28879# vssd1 0.53fF $ **FLOATING
C3629 a_6829_29199# vssd1 0.17fF $ **FLOATING
C3630 _1259_.X vssd1 5.48fF $ **FLOATING
C3631 a_5639_28879# vssd1 0.53fF $ **FLOATING
C3632 a_4719_28879# vssd1 0.53fF $ **FLOATING
C3633 _0909_.X vssd1 11.37fF $ **FLOATING
C3634 _1490_.A vssd1 2.39fF $ **FLOATING
C3635 a_22063_29098# vssd1 0.52fF $ **FLOATING
C3636 a_20947_28879# vssd1 0.61fF $ **FLOATING
C3637 a_21115_28853# vssd1 0.82fF $ **FLOATING
C3638 a_20522_28879# vssd1 0.63fF $ **FLOATING
C3639 a_20690_28853# vssd1 0.58fF $ **FLOATING
C3640 a_20249_28885# vssd1 1.43fF $ **FLOATING
C3641 _1870_.D vssd1 1.44fF $ **FLOATING
C3642 a_20083_28885# vssd1 1.81fF $ **FLOATING
C3643 a_19204_28995# vssd1 0.50fF $ **FLOATING
C3644 _1870_.Q vssd1 5.37fF $ **FLOATING
C3645 _1484_.B vssd1 14.26fF $ **FLOATING
C3646 a_18187_28879# vssd1 0.61fF $ **FLOATING
C3647 a_18355_28853# vssd1 0.82fF $ **FLOATING
C3648 a_17762_28879# vssd1 0.63fF $ **FLOATING
C3649 a_17930_28853# vssd1 0.58fF $ **FLOATING
C3650 a_17489_28885# vssd1 1.43fF $ **FLOATING
C3651 a_17323_28885# vssd1 1.81fF $ **FLOATING
C3652 a_15939_28879# vssd1 0.51fF $ **FLOATING
C3653 a_15759_28879# vssd1 0.60fF $ **FLOATING
C3654 _1424_.A_N vssd1 19.87fF $ **FLOATING
C3655 a_14467_28879# vssd1 0.51fF $ **FLOATING
C3656 a_14287_28879# vssd1 0.60fF $ **FLOATING
C3657 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref.TE vssd1 8.87fF $ **FLOATING
C3658 _1429_.A vssd1 4.97fF $ **FLOATING
C3659 a_11759_29098# vssd1 0.52fF $ **FLOATING
C3660 a_10419_28879# vssd1 0.51fF $ **FLOATING
C3661 a_10239_28879# vssd1 0.60fF $ **FLOATING
C3662 a_7479_28887# vssd1 0.65fF $ **FLOATING
C3663 a_6611_29111# vssd1 0.55fF $ **FLOATING
C3664 _1342_.B vssd1 11.81fF $ **FLOATING
C3665 a_3801_28981# vssd1 0.76fF $ **FLOATING
C3666 _0909_.C vssd1 2.65fF $ **FLOATING
C3667 _0909_.B vssd1 6.64fF $ **FLOATING
C3668 _0909_.A vssd1 20.45fF $ **FLOATING
C3669 a_1674_28879# vssd1 4.03fF $ **FLOATING
C3670 _1880_.Q vssd1 8.80fF $ **FLOATING
C3671 a_25497_29423# vssd1 0.23fF $ **FLOATING
C3672 a_27675_29588# vssd1 0.52fF $ **FLOATING
C3673 _1352_.A vssd1 9.78fF $ **FLOATING
C3674 a_27031_29588# vssd1 0.52fF $ **FLOATING
C3675 a_26007_29789# vssd1 0.61fF $ **FLOATING
C3676 a_26175_29691# vssd1 0.82fF $ **FLOATING
C3677 a_25582_29789# vssd1 0.63fF $ **FLOATING
C3678 a_25750_29535# vssd1 0.58fF $ **FLOATING
C3679 a_25309_29423# vssd1 1.43fF $ **FLOATING
C3680 _1880_.D vssd1 3.12fF $ **FLOATING
C3681 a_25143_29423# vssd1 1.81fF $ **FLOATING
C3682 _1880_.CLK vssd1 9.53fF $ **FLOATING
C3683 temp1.capload\[9\].cap.Y vssd1 0.28fF $ **FLOATING
C3684 _1869_.Q vssd1 8.93fF $ **FLOATING
C3685 a_22185_29423# vssd1 0.23fF $ **FLOATING
C3686 temp1.capload\[9\].cap.A vssd1 1.90fF $ **FLOATING
C3687 a_22695_29789# vssd1 0.61fF $ **FLOATING
C3688 a_22863_29691# vssd1 0.82fF $ **FLOATING
C3689 a_22270_29789# vssd1 0.63fF $ **FLOATING
C3690 a_22438_29535# vssd1 0.58fF $ **FLOATING
C3691 a_21997_29423# vssd1 1.43fF $ **FLOATING
C3692 a_21831_29423# vssd1 1.81fF $ **FLOATING
C3693 _1864_.Q vssd1 8.69fF $ **FLOATING
C3694 a_19793_29423# vssd1 0.23fF $ **FLOATING
C3695 a_20303_29789# vssd1 0.61fF $ **FLOATING
C3696 a_20471_29691# vssd1 0.82fF $ **FLOATING
C3697 a_19878_29789# vssd1 0.63fF $ **FLOATING
C3698 a_20046_29535# vssd1 0.58fF $ **FLOATING
C3699 a_19605_29423# vssd1 1.43fF $ **FLOATING
C3700 a_19439_29423# vssd1 1.81fF $ **FLOATING
C3701 a_17493_29423# vssd1 0.23fF $ **FLOATING
C3702 a_18003_29789# vssd1 0.61fF $ **FLOATING
C3703 a_18171_29691# vssd1 0.82fF $ **FLOATING
C3704 a_17578_29789# vssd1 0.63fF $ **FLOATING
C3705 a_17746_29535# vssd1 0.58fF $ **FLOATING
C3706 a_17305_29423# vssd1 1.43fF $ **FLOATING
C3707 a_17139_29423# vssd1 1.81fF $ **FLOATING
C3708 _1858_.Q vssd1 6.12fF $ **FLOATING
C3709 a_15377_29423# vssd1 0.23fF $ **FLOATING
C3710 a_15887_29789# vssd1 0.61fF $ **FLOATING
C3711 a_16055_29691# vssd1 0.82fF $ **FLOATING
C3712 a_15462_29789# vssd1 0.63fF $ **FLOATING
C3713 a_15630_29535# vssd1 0.58fF $ **FLOATING
C3714 a_15189_29423# vssd1 1.43fF $ **FLOATING
C3715 _1858_.D vssd1 3.80fF $ **FLOATING
C3716 a_15023_29423# vssd1 1.81fF $ **FLOATING
C3717 _1469_.X vssd1 2.76fF $ **FLOATING
C3718 _1902_.Q vssd1 6.24fF $ **FLOATING
C3719 a_12065_29423# vssd1 0.23fF $ **FLOATING
C3720 a_14287_29423# vssd1 0.70fF $ **FLOATING
C3721 _1469_.A vssd1 2.59fF $ **FLOATING
C3722 a_13599_29588# vssd1 0.52fF $ **FLOATING
C3723 a_12575_29789# vssd1 0.61fF $ **FLOATING
C3724 a_12743_29691# vssd1 0.82fF $ **FLOATING
C3725 a_12150_29789# vssd1 0.63fF $ **FLOATING
C3726 a_12318_29535# vssd1 0.58fF $ **FLOATING
C3727 a_11877_29423# vssd1 1.43fF $ **FLOATING
C3728 _1902_.D vssd1 6.95fF $ **FLOATING
C3729 a_11711_29423# vssd1 1.81fF $ **FLOATING
C3730 _1903_.Q vssd1 5.78fF $ **FLOATING
C3731 a_9949_29423# vssd1 0.23fF $ **FLOATING
C3732 a_10459_29789# vssd1 0.61fF $ **FLOATING
C3733 a_10627_29691# vssd1 0.82fF $ **FLOATING
C3734 a_10034_29789# vssd1 0.63fF $ **FLOATING
C3735 a_10202_29535# vssd1 0.58fF $ **FLOATING
C3736 a_9761_29423# vssd1 1.43fF $ **FLOATING
C3737 _1903_.D vssd1 7.41fF $ **FLOATING
C3738 a_9595_29423# vssd1 1.81fF $ **FLOATING
C3739 _1760_.X vssd1 12.67fF $ **FLOATING
C3740 a_8215_29423# vssd1 0.53fF $ **FLOATING
C3741 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 13.73fF $ **FLOATING
C3742 a_7387_29423# vssd1 0.53fF $ **FLOATING
C3743 a_6559_29423# vssd1 0.53fF $ **FLOATING
C3744 a_5731_29423# vssd1 0.53fF $ **FLOATING
C3745 a_4903_29423# vssd1 0.53fF $ **FLOATING
C3746 a_4075_29423# vssd1 0.53fF $ **FLOATING
C3747 a_2309_29789# vssd1 0.85fF $ **FLOATING
C3748 _1760_.B vssd1 11.75fF $ **FLOATING
C3749 a_2143_29789# vssd1 0.60fF $ **FLOATING
C3750 _1760_.A_N vssd1 4.38fF $ **FLOATING
C3751 temp1.capload\[5\].cap.Y vssd1 0.28fF $ **FLOATING
C3752 temp1.capload\[8\].cap.Y vssd1 0.28fF $ **FLOATING
C3753 temp1.capload\[7\].cap.Y vssd1 0.28fF $ **FLOATING
C3754 _1843_.Q vssd1 6.25fF $ **FLOATING
C3755 a_23197_29967# vssd1 0.23fF $ **FLOATING
C3756 temp1.capload\[12\].cap.Y vssd1 0.28fF $ **FLOATING
C3757 _1869_.D vssd1 1.82fF $ **FLOATING
C3758 a_19609_29967# vssd1 0.23fF $ **FLOATING
C3759 a_17217_29967# vssd1 0.23fF $ **FLOATING
C3760 a_15483_29967# vssd1 0.53fF $ **FLOATING
C3761 _1857_.Q vssd1 6.11fF $ **FLOATING
C3762 a_13077_29967# vssd1 0.23fF $ **FLOATING
C3763 a_11711_29967# vssd1 0.53fF $ **FLOATING
C3764 a_10133_29967# vssd1 0.23fF $ **FLOATING
C3765 a_8937_29967# vssd1 0.23fF $ **FLOATING
C3766 _1463_.A vssd1 9.64fF $ **FLOATING
C3767 a_5087_29967# vssd1 0.44fF $ **FLOATING
C3768 a_1975_29967# vssd1 0.22fF $ **FLOATING
C3769 _1555_.X vssd1 3.59fF $ **FLOATING
C3770 clkbuf_0_temp1.i_precharge_n.X vssd1 6.27fF $ **FLOATING
C3771 _1775_.X vssd1 1.50fF $ **FLOATING
C3772 _1456_.A vssd1 11.75fF $ **FLOATING
C3773 a_27859_30186# vssd1 0.52fF $ **FLOATING
C3774 temp1.inv2_2.A vssd1 14.25fF $ **FLOATING
C3775 temp1.capload\[5\].cap.A vssd1 2.60fF $ **FLOATING
C3776 temp1.capload\[7\].cap.A vssd1 1.97fF $ **FLOATING
C3777 a_23707_29967# vssd1 0.61fF $ **FLOATING
C3778 a_23875_29941# vssd1 0.82fF $ **FLOATING
C3779 a_23282_29967# vssd1 0.63fF $ **FLOATING
C3780 a_23450_29941# vssd1 0.58fF $ **FLOATING
C3781 a_23009_29973# vssd1 1.43fF $ **FLOATING
C3782 _1843_.D vssd1 3.13fF $ **FLOATING
C3783 a_22843_29973# vssd1 1.81fF $ **FLOATING
C3784 temp1.capload\[12\].cap.A vssd1 2.00fF $ **FLOATING
C3785 _1485_.A vssd1 1.70fF $ **FLOATING
C3786 a_20775_30186# vssd1 0.52fF $ **FLOATING
C3787 _1481_.A vssd1 4.05fF $ **FLOATING
C3788 a_20131_30186# vssd1 0.52fF $ **FLOATING
C3789 a_19432_29967# vssd1 0.50fF $ **FLOATING
C3790 a_19326_29967# vssd1 0.58fF $ **FLOATING
C3791 a_19149_29967# vssd1 0.50fF $ **FLOATING
C3792 a_18830_29967# vssd1 0.54fF $ **FLOATING
C3793 fanout33.A vssd1 13.78fF $ **FLOATING
C3794 a_17727_29967# vssd1 0.61fF $ **FLOATING
C3795 a_17895_29941# vssd1 0.82fF $ **FLOATING
C3796 a_17302_29967# vssd1 0.63fF $ **FLOATING
C3797 a_17470_29941# vssd1 0.58fF $ **FLOATING
C3798 a_17029_29973# vssd1 1.43fF $ **FLOATING
C3799 a_16863_29973# vssd1 1.81fF $ **FLOATING
C3800 temp1.dcdc.A vssd1 7.15fF $ **FLOATING
C3801 a_14743_29967# vssd1 0.51fF $ **FLOATING
C3802 _1867_.Q vssd1 5.68fF $ **FLOATING
C3803 a_14563_29967# vssd1 0.60fF $ **FLOATING
C3804 a_13587_29967# vssd1 0.61fF $ **FLOATING
C3805 a_13755_29941# vssd1 0.82fF $ **FLOATING
C3806 a_13162_29967# vssd1 0.63fF $ **FLOATING
C3807 a_13330_29941# vssd1 0.58fF $ **FLOATING
C3808 a_12889_29973# vssd1 1.43fF $ **FLOATING
C3809 _1456_.X vssd1 7.59fF $ **FLOATING
C3810 a_12723_29973# vssd1 1.81fF $ **FLOATING
C3811 a_10643_29967# vssd1 0.61fF $ **FLOATING
C3812 a_10811_29941# vssd1 0.82fF $ **FLOATING
C3813 a_10218_29967# vssd1 0.63fF $ **FLOATING
C3814 a_10386_29941# vssd1 0.58fF $ **FLOATING
C3815 a_9945_29973# vssd1 1.43fF $ **FLOATING
C3816 a_9779_29973# vssd1 1.81fF $ **FLOATING
C3817 a_8760_29967# vssd1 0.50fF $ **FLOATING
C3818 a_8654_29967# vssd1 0.58fF $ **FLOATING
C3819 a_8477_29967# vssd1 0.50fF $ **FLOATING
C3820 a_8158_29967# vssd1 0.54fF $ **FLOATING
C3821 a_7383_29967# vssd1 0.51fF $ **FLOATING
C3822 a_7203_29967# vssd1 0.60fF $ **FLOATING
C3823 _1555_.A vssd1 4.37fF $ **FLOATING
C3824 a_6607_30186# vssd1 0.52fF $ **FLOATING
C3825 _1242_.B1 vssd1 14.15fF $ **FLOATING
C3826 _1242_.A1 vssd1 15.27fF $ **FLOATING
C3827 a_2962_29967# vssd1 4.03fF $ **FLOATING
C3828 clkbuf_0_temp1.i_precharge_n.A vssd1 13.00fF $ **FLOATING
C3829 _1775_.C1 vssd1 23.08fF $ **FLOATING
C3830 _1775_.B1 vssd1 4.02fF $ **FLOATING
C3831 temp1.inv2_2.Y vssd1 11.56fF $ **FLOATING
C3832 _1775_.A2 vssd1 23.71fF $ **FLOATING
C3833 _1242_.A2 vssd1 15.90fF $ **FLOATING
C3834 a_1735_29941# vssd1 1.12fF $ **FLOATING
C3835 _1450_.X vssd1 9.11fF $ **FLOATING
C3836 _1450_.A vssd1 10.71fF $ **FLOATING
C3837 a_27859_30676# vssd1 0.52fF $ **FLOATING
C3838 temp1.capload\[4\].cap_49.HI vssd1 0.42fF $ **FLOATING
C3839 temp1.capload\[2\].cap_47.LO vssd1 2.98fF $ **FLOATING
C3840 temp1.capload\[2\].cap_47.HI vssd1 0.42fF $ **FLOATING
C3841 temp1.capload\[15\].cap_45.HI vssd1 0.42fF $ **FLOATING
C3842 temp1.capload\[1\].cap.Y vssd1 0.28fF $ **FLOATING
C3843 temp1.capload\[1\].cap.A vssd1 1.13fF $ **FLOATING
C3844 temp1.capload\[1\].cap_46.HI vssd1 0.42fF $ **FLOATING
C3845 temp1.capload\[13\].cap.Y vssd1 0.28fF $ **FLOATING
C3846 _1872_.Q vssd1 4.21fF $ **FLOATING
C3847 a_21725_30511# vssd1 0.23fF $ **FLOATING
C3848 a_22235_30877# vssd1 0.61fF $ **FLOATING
C3849 a_22403_30779# vssd1 0.82fF $ **FLOATING
C3850 a_21810_30877# vssd1 0.63fF $ **FLOATING
C3851 a_21978_30623# vssd1 0.58fF $ **FLOATING
C3852 a_21537_30511# vssd1 1.43fF $ **FLOATING
C3853 a_21371_30511# vssd1 1.81fF $ **FLOATING
C3854 a_19885_30511# vssd1 0.23fF $ **FLOATING
C3855 a_20395_30877# vssd1 0.61fF $ **FLOATING
C3856 a_20563_30779# vssd1 0.82fF $ **FLOATING
C3857 a_19970_30877# vssd1 0.63fF $ **FLOATING
C3858 a_20138_30623# vssd1 0.58fF $ **FLOATING
C3859 a_19697_30511# vssd1 1.43fF $ **FLOATING
C3860 _1871_.D vssd1 1.31fF $ **FLOATING
C3861 a_19531_30511# vssd1 1.81fF $ **FLOATING
C3862 _1471_.X vssd1 2.10fF $ **FLOATING
C3863 _1853_.Q vssd1 8.40fF $ **FLOATING
C3864 a_14641_30511# vssd1 0.23fF $ **FLOATING
C3865 _1425_.A vssd1 2.38fF $ **FLOATING
C3866 a_18475_30676# vssd1 0.52fF $ **FLOATING
C3867 _1471_.A vssd1 3.87fF $ **FLOATING
C3868 a_17831_30676# vssd1 0.52fF $ **FLOATING
C3869 a_16955_30511# vssd1 0.53fF $ **FLOATING
C3870 a_16127_30511# vssd1 0.53fF $ **FLOATING
C3871 a_15151_30877# vssd1 0.61fF $ **FLOATING
C3872 a_15319_30779# vssd1 0.82fF $ **FLOATING
C3873 a_14726_30877# vssd1 0.63fF $ **FLOATING
C3874 a_14894_30623# vssd1 0.58fF $ **FLOATING
C3875 a_14453_30511# vssd1 1.43fF $ **FLOATING
C3876 a_14287_30511# vssd1 1.81fF $ **FLOATING
C3877 a_13367_30511# vssd1 0.53fF $ **FLOATING
C3878 a_12631_30511# vssd1 0.65fF $ **FLOATING
C3879 _1349_.A vssd1 3.94fF $ **FLOATING
C3880 a_8385_30511# vssd1 0.23fF $ **FLOATING
C3881 _1330_.X vssd1 9.85fF $ **FLOATING
C3882 clkbuf_1_1__f_net57.X vssd1 14.26fF $ **FLOATING
C3883 a_10506_30511# vssd1 4.03fF $ **FLOATING
C3884 a_9595_30511# vssd1 0.53fF $ **FLOATING
C3885 a_8208_30511# vssd1 0.50fF $ **FLOATING
C3886 a_8102_30511# vssd1 0.58fF $ **FLOATING
C3887 a_7925_30511# vssd1 0.50fF $ **FLOATING
C3888 a_7606_30511# vssd1 0.54fF $ **FLOATING
C3889 a_6559_30511# vssd1 0.53fF $ **FLOATING
C3890 a_5731_30511# vssd1 0.53fF $ **FLOATING
C3891 a_4213_30663# vssd1 0.77fF $ **FLOATING
C3892 a_4035_30485# vssd1 0.83fF $ **FLOATING
C3893 a_1674_30511# vssd1 4.03fF $ **FLOATING
C3894 temp1.capload\[0\].cap_39.HI vssd1 0.42fF $ **FLOATING
C3895 temp1.capload\[0\].cap.Y vssd1 0.28fF $ **FLOATING
C3896 a_27215_31274# vssd1 0.52fF $ **FLOATING
C3897 temp1.capload\[0\].cap.A vssd1 1.40fF $ **FLOATING
C3898 temp1.capload\[11\].cap_41.HI vssd1 0.42fF $ **FLOATING
C3899 temp1.capload\[10\].cap_40.HI vssd1 0.42fF $ **FLOATING
C3900 _1447_.X vssd1 5.89fF $ **FLOATING
C3901 temp1.capload\[4\].cap.Y vssd1 0.28fF $ **FLOATING
C3902 _1874_.Q vssd1 8.22fF $ **FLOATING
C3903 a_22369_31055# vssd1 0.23fF $ **FLOATING
C3904 _1487_.X vssd1 1.16fF $ **FLOATING
C3905 a_19701_31055# vssd1 0.23fF $ **FLOATING
C3906 _1862_.Q vssd1 6.22fF $ **FLOATING
C3907 a_17861_31055# vssd1 0.23fF $ **FLOATING
C3908 _1861_.Q vssd1 6.31fF $ **FLOATING
C3909 a_15285_31055# vssd1 0.23fF $ **FLOATING
C3910 _1856_.Q vssd1 8.88fF $ **FLOATING
C3911 a_13445_31055# vssd1 0.23fF $ **FLOATING
C3912 a_12263_31055# vssd1 0.53fF $ **FLOATING
C3913 a_9489_31055# vssd1 0.23fF $ **FLOATING
C3914 a_8307_31055# vssd1 0.53fF $ **FLOATING
C3915 a_7479_31055# vssd1 0.53fF $ **FLOATING
C3916 a_6651_31055# vssd1 0.53fF $ **FLOATING
C3917 a_5639_31055# vssd1 0.53fF $ **FLOATING
C3918 a_4811_31055# vssd1 0.53fF $ **FLOATING
C3919 clkbuf_0_net57.X vssd1 6.77fF $ **FLOATING
C3920 a_1683_31055# vssd1 0.53fF $ **FLOATING
C3921 _1447_.A vssd1 10.67fF $ **FLOATING
C3922 a_24547_31274# vssd1 0.52fF $ **FLOATING
C3923 temp1.capload\[4\].cap.A vssd1 2.19fF $ **FLOATING
C3924 a_22879_31055# vssd1 0.61fF $ **FLOATING
C3925 a_23047_31029# vssd1 0.82fF $ **FLOATING
C3926 a_22454_31055# vssd1 0.63fF $ **FLOATING
C3927 a_22622_31029# vssd1 0.58fF $ **FLOATING
C3928 a_22181_31061# vssd1 1.43fF $ **FLOATING
C3929 _1874_.D vssd1 3.04fF $ **FLOATING
C3930 a_22015_31061# vssd1 1.81fF $ **FLOATING
C3931 a_21235_31274# vssd1 0.52fF $ **FLOATING
C3932 a_20211_31055# vssd1 0.61fF $ **FLOATING
C3933 a_20379_31029# vssd1 0.82fF $ **FLOATING
C3934 a_19786_31055# vssd1 0.63fF $ **FLOATING
C3935 a_19954_31029# vssd1 0.58fF $ **FLOATING
C3936 a_19513_31061# vssd1 1.43fF $ **FLOATING
C3937 a_19347_31061# vssd1 1.81fF $ **FLOATING
C3938 a_18371_31055# vssd1 0.61fF $ **FLOATING
C3939 a_18539_31029# vssd1 0.82fF $ **FLOATING
C3940 a_17946_31055# vssd1 0.63fF $ **FLOATING
C3941 a_18114_31029# vssd1 0.58fF $ **FLOATING
C3942 a_17673_31061# vssd1 1.43fF $ **FLOATING
C3943 a_17507_31061# vssd1 1.81fF $ **FLOATING
C3944 _1538_.A vssd1 2.79fF $ **FLOATING
C3945 a_16911_31274# vssd1 0.52fF $ **FLOATING
C3946 a_15795_31055# vssd1 0.61fF $ **FLOATING
C3947 a_15963_31029# vssd1 0.82fF $ **FLOATING
C3948 a_15370_31055# vssd1 0.63fF $ **FLOATING
C3949 a_15538_31029# vssd1 0.58fF $ **FLOATING
C3950 a_15097_31061# vssd1 1.43fF $ **FLOATING
C3951 _1465_.X vssd1 5.92fF $ **FLOATING
C3952 a_14931_31061# vssd1 1.81fF $ **FLOATING
C3953 a_13955_31055# vssd1 0.61fF $ **FLOATING
C3954 a_14123_31029# vssd1 0.82fF $ **FLOATING
C3955 a_13530_31055# vssd1 0.63fF $ **FLOATING
C3956 a_13698_31029# vssd1 0.58fF $ **FLOATING
C3957 a_13257_31061# vssd1 1.43fF $ **FLOATING
C3958 _1856_.D vssd1 7.73fF $ **FLOATING
C3959 a_13091_31061# vssd1 1.81fF $ **FLOATING
C3960 _1479_.A vssd1 2.84fF $ **FLOATING
C3961 a_11023_31274# vssd1 0.52fF $ **FLOATING
C3962 a_9999_31055# vssd1 0.61fF $ **FLOATING
C3963 a_10167_31029# vssd1 0.82fF $ **FLOATING
C3964 a_9574_31055# vssd1 0.63fF $ **FLOATING
C3965 a_9742_31029# vssd1 0.58fF $ **FLOATING
C3966 a_9301_31061# vssd1 1.43fF $ **FLOATING
C3967 _1860_.D vssd1 9.31fF $ **FLOATING
C3968 a_9135_31061# vssd1 1.81fF $ **FLOATING
C3969 _1860_.CLK vssd1 12.00fF $ **FLOATING
C3970 a_2594_31055# vssd1 4.03fF $ **FLOATING
C3971 clkbuf_0_net57.A vssd1 12.22fF $ **FLOATING
C3972 _1347_.Y vssd1 14.58fF $ **FLOATING
C3973 temp1.capload\[8\].cap_53.LO vssd1 2.71fF $ **FLOATING
C3974 temp1.capload\[8\].cap_53.HI vssd1 0.42fF $ **FLOATING
C3975 _1353_.Y vssd1 11.97fF $ **FLOATING
C3976 _1873_.Q vssd1 8.52fF $ **FLOATING
C3977 a_24945_31599# vssd1 0.23fF $ **FLOATING
C3978 _1353_.A vssd1 20.21fF $ **FLOATING
C3979 _1353_.B vssd1 9.67fF $ **FLOATING
C3980 a_25455_31965# vssd1 0.61fF $ **FLOATING
C3981 a_25623_31867# vssd1 0.82fF $ **FLOATING
C3982 a_25030_31965# vssd1 0.63fF $ **FLOATING
C3983 a_25198_31711# vssd1 0.58fF $ **FLOATING
C3984 a_24757_31599# vssd1 1.43fF $ **FLOATING
C3985 _1873_.D vssd1 3.08fF $ **FLOATING
C3986 a_24591_31599# vssd1 1.81fF $ **FLOATING
C3987 _1475_.X vssd1 6.05fF $ **FLOATING
C3988 _1842_.Q vssd1 5.84fF $ **FLOATING
C3989 a_21909_31599# vssd1 0.23fF $ **FLOATING
C3990 a_23443_31764# vssd1 0.52fF $ **FLOATING
C3991 a_22419_31965# vssd1 0.61fF $ **FLOATING
C3992 a_22587_31867# vssd1 0.82fF $ **FLOATING
C3993 a_21994_31965# vssd1 0.63fF $ **FLOATING
C3994 a_22162_31711# vssd1 0.58fF $ **FLOATING
C3995 a_21721_31599# vssd1 1.43fF $ **FLOATING
C3996 _1842_.D vssd1 2.62fF $ **FLOATING
C3997 a_21555_31599# vssd1 1.81fF $ **FLOATING
C3998 _1873_.CLK vssd1 14.51fF $ **FLOATING
C3999 _1897_.Q vssd1 7.61fF $ **FLOATING
C4000 a_19793_31599# vssd1 0.23fF $ **FLOATING
C4001 a_20303_31965# vssd1 0.61fF $ **FLOATING
C4002 a_20471_31867# vssd1 0.82fF $ **FLOATING
C4003 a_19878_31965# vssd1 0.63fF $ **FLOATING
C4004 a_20046_31711# vssd1 0.58fF $ **FLOATING
C4005 a_19605_31599# vssd1 1.43fF $ **FLOATING
C4006 a_19439_31599# vssd1 1.81fF $ **FLOATING
C4007 _1859_.Q vssd1 9.78fF $ **FLOATING
C4008 a_16849_31599# vssd1 0.23fF $ **FLOATING
C4009 a_18335_31599# vssd1 0.53fF $ **FLOATING
C4010 a_17359_31965# vssd1 0.61fF $ **FLOATING
C4011 a_17527_31867# vssd1 0.82fF $ **FLOATING
C4012 a_16934_31965# vssd1 0.63fF $ **FLOATING
C4013 a_17102_31711# vssd1 0.58fF $ **FLOATING
C4014 a_16661_31599# vssd1 1.43fF $ **FLOATING
C4015 _1859_.D vssd1 3.09fF $ **FLOATING
C4016 a_16495_31599# vssd1 1.81fF $ **FLOATING
C4017 clkbuf_0_temp1.dcdel_capnode_notouch_.X vssd1 7.58fF $ **FLOATING
C4018 _1486_.X vssd1 5.22fF $ **FLOATING
C4019 _1473_.X vssd1 5.10fF $ **FLOATING
C4020 _1855_.Q vssd1 5.59fF $ **FLOATING
C4021 a_11053_31599# vssd1 0.23fF $ **FLOATING
C4022 a_14370_31599# vssd1 4.03fF $ **FLOATING
C4023 clkbuf_0_temp1.dcdel_capnode_notouch_.A vssd1 2.52fF $ **FLOATING
C4024 a_13455_31965# vssd1 0.51fF $ **FLOATING
C4025 _1486_.B vssd1 6.77fF $ **FLOATING
C4026 a_13275_31965# vssd1 0.60fF $ **FLOATING
C4027 _1473_.A vssd1 2.98fF $ **FLOATING
C4028 a_12679_31764# vssd1 0.52fF $ **FLOATING
C4029 a_11563_31965# vssd1 0.61fF $ **FLOATING
C4030 a_11731_31867# vssd1 0.82fF $ **FLOATING
C4031 a_11138_31965# vssd1 0.63fF $ **FLOATING
C4032 a_11306_31711# vssd1 0.58fF $ **FLOATING
C4033 a_10865_31599# vssd1 1.43fF $ **FLOATING
C4034 _1855_.D vssd1 11.38fF $ **FLOATING
C4035 a_10699_31599# vssd1 1.81fF $ **FLOATING
C4036 _1855_.CLK vssd1 12.45fF $ **FLOATING
C4037 _1464_.X vssd1 9.50fF $ **FLOATING
C4038 a_9775_31965# vssd1 0.51fF $ **FLOATING
C4039 _1464_.B vssd1 3.75fF $ **FLOATING
C4040 a_9595_31965# vssd1 0.60fF $ **FLOATING
C4041 a_8307_31599# vssd1 0.65fF $ **FLOATING
C4042 fanout12.A vssd1 11.34fF $ **FLOATING
C4043 _1451_.X vssd1 11.55fF $ **FLOATING
C4044 _1243_.Y vssd1 6.36fF $ **FLOATING
C4045 _1329_.X vssd1 2.34fF $ **FLOATING
C4046 a_7567_31965# vssd1 0.51fF $ **FLOATING
C4047 _1451_.B vssd1 6.83fF $ **FLOATING
C4048 a_7387_31965# vssd1 0.60fF $ **FLOATING
C4049 a_6559_31599# vssd1 0.53fF $ **FLOATING
C4050 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.A vssd1 4.79fF $ **FLOATING
C4051 a_5731_31599# vssd1 0.53fF $ **FLOATING
C4052 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd.TE vssd1 6.83fF $ **FLOATING
C4053 a_4903_31599# vssd1 0.53fF $ **FLOATING
C4054 a_4075_31599# vssd1 0.53fF $ **FLOATING
C4055 _1243_.A vssd1 5.91fF $ **FLOATING
C4056 _1329_.S vssd1 14.72fF $ **FLOATING
C4057 _1329_.A0 vssd1 3.82fF $ **FLOATING
C4058 _1329_.A1 vssd1 6.12fF $ **FLOATING
C4059 a_2281_31751# vssd1 0.77fF $ **FLOATING
C4060 a_2103_31573# vssd1 0.83fF $ **FLOATING
C4061 io_out[7] vssd1 12.61fF
C4062 a_27811_32143# vssd1 0.52fF $ **FLOATING
C4063 temp1.capload\[13\].cap_43.LO vssd1 2.39fF $ **FLOATING
C4064 temp1.capload\[6\].cap_51.HI vssd1 0.42fF $ **FLOATING
C4065 temp1.capload\[6\].cap.Y vssd1 0.28fF $ **FLOATING
C4066 temp1.capload\[6\].cap_51.LO vssd1 1.33fF $ **FLOATING
C4067 temp1.capload\[6\].cap.B vssd1 12.23fF $ **FLOATING
C4068 temp1.capload\[14\].cap_44.LO vssd1 4.44fF $ **FLOATING
C4069 temp1.capload\[13\].cap_43.HI vssd1 0.42fF $ **FLOATING
C4070 temp1.capload\[14\].cap_44.HI vssd1 0.42fF $ **FLOATING
C4071 _1477_.X vssd1 4.88fF $ **FLOATING
C4072 temp1.capload\[15\].cap.Y vssd1 0.28fF $ **FLOATING
C4073 temp1.capload\[11\].cap.Y vssd1 0.28fF $ **FLOATING
C4074 _1896_.Q vssd1 8.27fF $ **FLOATING
C4075 a_20161_32143# vssd1 0.23fF $ **FLOATING
C4076 _1841_.Q vssd1 4.95fF $ **FLOATING
C4077 a_17861_32143# vssd1 0.23fF $ **FLOATING
C4078 _1540_.X vssd1 2.35fF $ **FLOATING
C4079 _1868_.Q vssd1 6.39fF $ **FLOATING
C4080 a_15285_32143# vssd1 0.23fF $ **FLOATING
C4081 temp1.capload\[10\].cap.Y vssd1 0.28fF $ **FLOATING
C4082 _1474_.X vssd1 5.85fF $ **FLOATING
C4083 _1467_.X vssd1 3.89fF $ **FLOATING
C4084 a_10791_32143# vssd1 0.53fF $ **FLOATING
C4085 a_9963_32143# vssd1 0.53fF $ **FLOATING
C4086 a_9135_32143# vssd1 0.53fF $ **FLOATING
C4087 a_8215_32143# vssd1 0.53fF $ **FLOATING
C4088 a_7387_32143# vssd1 0.53fF $ **FLOATING
C4089 a_6559_32143# vssd1 0.53fF $ **FLOATING
C4090 a_5639_32143# vssd1 0.53fF $ **FLOATING
C4091 a_4811_32143# vssd1 0.53fF $ **FLOATING
C4092 a_3983_32143# vssd1 0.53fF $ **FLOATING
C4093 a_3063_32143# vssd1 0.53fF $ **FLOATING
C4094 _1477_.A vssd1 6.41fF $ **FLOATING
C4095 a_23351_32362# vssd1 0.52fF $ **FLOATING
C4096 temp1.capload\[15\].cap.A vssd1 2.63fF $ **FLOATING
C4097 temp1.capload\[11\].cap.A vssd1 3.35fF $ **FLOATING
C4098 a_20671_32143# vssd1 0.61fF $ **FLOATING
C4099 a_20839_32117# vssd1 0.82fF $ **FLOATING
C4100 a_20246_32143# vssd1 0.63fF $ **FLOATING
C4101 a_20414_32117# vssd1 0.58fF $ **FLOATING
C4102 a_19973_32149# vssd1 1.43fF $ **FLOATING
C4103 _1896_.D vssd1 2.66fF $ **FLOATING
C4104 a_19807_32149# vssd1 1.81fF $ **FLOATING
C4105 _1896_.CLK vssd1 5.29fF $ **FLOATING
C4106 a_18371_32143# vssd1 0.61fF $ **FLOATING
C4107 a_18539_32117# vssd1 0.82fF $ **FLOATING
C4108 a_17946_32143# vssd1 0.63fF $ **FLOATING
C4109 a_18114_32117# vssd1 0.58fF $ **FLOATING
C4110 a_17673_32149# vssd1 1.43fF $ **FLOATING
C4111 _1841_.D vssd1 7.29fF $ **FLOATING
C4112 a_17507_32149# vssd1 1.81fF $ **FLOATING
C4113 _1540_.A vssd1 2.90fF $ **FLOATING
C4114 a_16911_32362# vssd1 0.52fF $ **FLOATING
C4115 a_15795_32143# vssd1 0.61fF $ **FLOATING
C4116 a_15963_32117# vssd1 0.82fF $ **FLOATING
C4117 a_15370_32143# vssd1 0.63fF $ **FLOATING
C4118 a_15538_32117# vssd1 0.58fF $ **FLOATING
C4119 a_15097_32149# vssd1 1.43fF $ **FLOATING
C4120 _1868_.D vssd1 3.35fF $ **FLOATING
C4121 a_14931_32149# vssd1 1.81fF $ **FLOATING
C4122 _1841_.CLK vssd1 11.55fF $ **FLOATING
C4123 temp1.capload\[10\].cap.A vssd1 6.83fF $ **FLOATING
C4124 temp1.capload\[15\].cap.B vssd1 14.71fF $ **FLOATING
C4125 a_13455_32143# vssd1 0.51fF $ **FLOATING
C4126 _1474_.B vssd1 7.75fF $ **FLOATING
C4127 a_13275_32143# vssd1 0.60fF $ **FLOATING
C4128 a_12535_32143# vssd1 0.51fF $ **FLOATING
C4129 _1476_.B vssd1 7.30fF $ **FLOATING
C4130 a_12355_32143# vssd1 0.60fF $ **FLOATING
C4131 _1474_.A_N vssd1 16.12fF $ **FLOATING
C4132 _1467_.A vssd1 3.11fF $ **FLOATING
C4133 a_11759_32362# vssd1 0.52fF $ **FLOATING
C4134 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref.TE vssd1 12.35fF $ **FLOATING
C4135 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 9.21fF $ **FLOATING
C4136 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 12.31fF $ **FLOATING
C4137 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd.Z vssd1 66.42fF $ **FLOATING
C4138 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 17.53fF $ **FLOATING
C4139 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.A vssd1 15.87fF $ **FLOATING
C4140 temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd.TE vssd1 16.37fF $ **FLOATING
C4141 _1338_.A vssd1 12.04fF $ **FLOATING
C4142 _1337_.S vssd1 12.63fF $ **FLOATING
C4143 _1337_.A1 vssd1 6.80fF $ **FLOATING
C4144 _1337_.A0 vssd1 14.44fF $ **FLOATING
C4145 a_2005_32375# vssd1 0.77fF $ **FLOATING
C4146 a_1827_32117# vssd1 0.83fF $ **FLOATING
C4147 vccd1 vssd1 3429.07fF
.ends
