magic
tech sky130A
magscale 1 2
timestamp 1681905124
<< viali >>
rect 4353 32521 4387 32555
rect 5181 32521 5215 32555
rect 8585 32521 8619 32555
rect 9505 32521 9539 32555
rect 11069 32521 11103 32555
rect 3341 32453 3375 32487
rect 1593 32385 1627 32419
rect 3985 32385 4019 32419
rect 12357 32385 12391 32419
rect 12541 32385 12575 32419
rect 14289 32385 14323 32419
rect 14473 32385 14507 32419
rect 14933 32385 14967 32419
rect 15117 32385 15151 32419
rect 15577 32385 15611 32419
rect 15761 32385 15795 32419
rect 4813 32317 4847 32351
rect 8217 32317 8251 32351
rect 9137 32317 9171 32351
rect 9505 32317 9539 32351
rect 10701 32317 10735 32351
rect 4353 32249 4387 32283
rect 5181 32249 5215 32283
rect 6009 32249 6043 32283
rect 8585 32249 8619 32283
rect 11069 32249 11103 32283
rect 11897 32249 11931 32283
rect 6745 32181 6779 32215
rect 7389 32181 7423 32215
rect 10149 32181 10183 32215
rect 13185 32181 13219 32215
rect 4537 31977 4571 32011
rect 6745 31977 6779 32011
rect 7389 31977 7423 32011
rect 5917 31909 5951 31943
rect 9321 31909 9355 31943
rect 13277 31909 13311 31943
rect 3341 31841 3375 31875
rect 9873 31841 9907 31875
rect 11069 31841 11103 31875
rect 1593 31773 1627 31807
rect 3985 31773 4019 31807
rect 4261 31773 4295 31807
rect 4405 31773 4439 31807
rect 5549 31773 5583 31807
rect 8217 31773 8251 31807
rect 8585 31773 8619 31807
rect 10241 31773 10275 31807
rect 10701 31773 10735 31807
rect 11529 31773 11563 31807
rect 11897 31773 11931 31807
rect 12357 31773 12391 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 14933 31773 14967 31807
rect 15117 31773 15151 31807
rect 15577 31773 15611 31807
rect 15761 31773 15795 31807
rect 16221 31773 16255 31807
rect 16405 31773 16439 31807
rect 4169 31705 4203 31739
rect 5917 31637 5951 31671
rect 8585 31637 8619 31671
rect 10241 31637 10275 31671
rect 11069 31637 11103 31671
rect 11897 31637 11931 31671
rect 12541 31637 12575 31671
rect 5181 31433 5215 31467
rect 6009 31433 6043 31467
rect 7481 31433 7515 31467
rect 8309 31433 8343 31467
rect 9137 31433 9171 31467
rect 10333 31433 10367 31467
rect 11161 31433 11195 31467
rect 12081 31433 12115 31467
rect 14105 31433 14139 31467
rect 14933 31433 14967 31467
rect 1777 31297 1811 31331
rect 2053 31297 2087 31331
rect 2605 31297 2639 31331
rect 4813 31297 4847 31331
rect 5641 31297 5675 31331
rect 7481 31297 7515 31331
rect 8309 31297 8343 31331
rect 9137 31297 9171 31331
rect 10333 31297 10367 31331
rect 10793 31297 10827 31331
rect 11161 31297 11195 31331
rect 13093 31297 13127 31331
rect 2145 31229 2179 31263
rect 7113 31229 7147 31263
rect 7941 31229 7975 31263
rect 8769 31229 8803 31263
rect 9965 31229 9999 31263
rect 11713 31229 11747 31263
rect 13737 31229 13771 31263
rect 14565 31229 14599 31263
rect 5181 31161 5215 31195
rect 6009 31161 6043 31195
rect 12081 31161 12115 31195
rect 14105 31161 14139 31195
rect 14933 31161 14967 31195
rect 3893 31093 3927 31127
rect 13185 31093 13219 31127
rect 6285 30889 6319 30923
rect 7665 30889 7699 30923
rect 8585 30889 8619 30923
rect 12173 30889 12207 30923
rect 9689 30821 9723 30855
rect 10517 30821 10551 30855
rect 11345 30821 11379 30855
rect 3433 30753 3467 30787
rect 4077 30753 4111 30787
rect 8217 30753 8251 30787
rect 8585 30753 8619 30787
rect 9321 30753 9355 30787
rect 10149 30753 10183 30787
rect 10977 30753 11011 30787
rect 11805 30753 11839 30787
rect 12173 30753 12207 30787
rect 13737 30753 13771 30787
rect 15945 30753 15979 30787
rect 1685 30685 1719 30719
rect 4261 30685 4295 30719
rect 4997 30685 5031 30719
rect 7297 30685 7331 30719
rect 7665 30685 7699 30719
rect 12633 30685 12667 30719
rect 13369 30685 13403 30719
rect 14841 30685 14875 30719
rect 15209 30685 15243 30719
rect 4537 30617 4571 30651
rect 15761 30617 15795 30651
rect 4445 30549 4479 30583
rect 9689 30549 9723 30583
rect 10517 30549 10551 30583
rect 11345 30549 11379 30583
rect 12817 30549 12851 30583
rect 13737 30549 13771 30583
rect 15209 30549 15243 30583
rect 6929 30345 6963 30379
rect 7757 30345 7791 30379
rect 9137 30345 9171 30379
rect 10333 30345 10367 30379
rect 11161 30345 11195 30379
rect 12725 30345 12759 30379
rect 13553 30345 13587 30379
rect 14381 30345 14415 30379
rect 15209 30345 15243 30379
rect 16037 30345 16071 30379
rect 2053 30277 2087 30311
rect 5181 30277 5215 30311
rect 1961 30209 1995 30243
rect 2145 30209 2179 30243
rect 2237 30209 2271 30243
rect 2421 30209 2455 30243
rect 2881 30209 2915 30243
rect 5365 30209 5399 30243
rect 5457 30209 5491 30243
rect 6561 30209 6595 30243
rect 7389 30209 7423 30243
rect 8769 30209 8803 30243
rect 9137 30209 9171 30243
rect 9965 30209 9999 30243
rect 10333 30209 10367 30243
rect 10793 30209 10827 30243
rect 11161 30209 11195 30243
rect 11713 30209 11747 30243
rect 11897 30209 11931 30243
rect 14013 30209 14047 30243
rect 14841 30209 14875 30243
rect 15669 30209 15703 30243
rect 5641 30141 5675 30175
rect 5733 30141 5767 30175
rect 12357 30141 12391 30175
rect 13185 30141 13219 30175
rect 14381 30141 14415 30175
rect 1777 30073 1811 30107
rect 6929 30073 6963 30107
rect 7757 30073 7791 30107
rect 12725 30073 12759 30107
rect 13553 30073 13587 30107
rect 15209 30073 15243 30107
rect 16037 30073 16071 30107
rect 4169 30005 4203 30039
rect 5457 29801 5491 29835
rect 9321 29801 9355 29835
rect 6561 29733 6595 29767
rect 11897 29733 11931 29767
rect 12909 29733 12943 29767
rect 8447 29665 8481 29699
rect 9965 29665 9999 29699
rect 10793 29665 10827 29699
rect 14841 29665 14875 29699
rect 16037 29665 16071 29699
rect 1685 29597 1719 29631
rect 3985 29597 4019 29631
rect 4261 29597 4295 29631
rect 4537 29597 4571 29631
rect 4813 29597 4847 29631
rect 6193 29597 6227 29631
rect 7481 29597 7515 29631
rect 7665 29597 7699 29631
rect 8344 29597 8378 29631
rect 10333 29597 10367 29631
rect 11161 29597 11195 29631
rect 12541 29597 12575 29631
rect 13369 29597 13403 29631
rect 13737 29597 13771 29631
rect 15209 29597 15243 29631
rect 15669 29597 15703 29631
rect 5273 29529 5307 29563
rect 11713 29529 11747 29563
rect 2973 29461 3007 29495
rect 4077 29461 4111 29495
rect 5457 29461 5491 29495
rect 5641 29461 5675 29495
rect 6561 29461 6595 29495
rect 7573 29461 7607 29495
rect 10333 29461 10367 29495
rect 11161 29461 11195 29495
rect 12909 29461 12943 29495
rect 13737 29461 13771 29495
rect 15209 29461 15243 29495
rect 16037 29461 16071 29495
rect 9965 29257 9999 29291
rect 11069 29257 11103 29291
rect 5273 29189 5307 29223
rect 1869 29121 1903 29155
rect 2053 29121 2087 29155
rect 2605 29121 2639 29155
rect 5457 29121 5491 29155
rect 6929 29121 6963 29155
rect 9781 29121 9815 29155
rect 10701 29121 10735 29155
rect 11069 29121 11103 29155
rect 11713 29121 11747 29155
rect 11897 29121 11931 29155
rect 13737 29121 13771 29155
rect 14565 29121 14599 29155
rect 15025 29121 15059 29155
rect 2145 29053 2179 29087
rect 4353 29053 4387 29087
rect 5733 29053 5767 29087
rect 7021 29053 7055 29087
rect 7205 29053 7239 29087
rect 8677 29053 8711 29087
rect 12357 29053 12391 29087
rect 12725 29053 12759 29087
rect 13369 29053 13403 29087
rect 14197 29053 14231 29087
rect 8033 28985 8067 29019
rect 9321 28985 9355 29019
rect 15209 28985 15243 29019
rect 5641 28917 5675 28951
rect 6561 28917 6595 28951
rect 12725 28917 12759 28951
rect 13737 28917 13771 28951
rect 14565 28917 14599 28951
rect 6837 28713 6871 28747
rect 9321 28713 9355 28747
rect 14657 28645 14691 28679
rect 11897 28577 11931 28611
rect 12725 28577 12759 28611
rect 13553 28577 13587 28611
rect 14289 28577 14323 28611
rect 2053 28509 2087 28543
rect 2320 28509 2354 28543
rect 3985 28509 4019 28543
rect 5917 28509 5951 28543
rect 6101 28509 6135 28543
rect 6653 28509 6687 28543
rect 7389 28509 7423 28543
rect 7573 28509 7607 28543
rect 8217 28509 8251 28543
rect 9781 28509 9815 28543
rect 9965 28509 9999 28543
rect 10425 28509 10459 28543
rect 10609 28509 10643 28543
rect 11529 28509 11563 28543
rect 12357 28509 12391 28543
rect 13185 28509 13219 28543
rect 4252 28441 4286 28475
rect 3433 28373 3467 28407
rect 5365 28373 5399 28407
rect 5917 28373 5951 28407
rect 7481 28373 7515 28407
rect 8033 28373 8067 28407
rect 11897 28373 11931 28407
rect 12725 28373 12759 28407
rect 13553 28373 13587 28407
rect 14657 28373 14691 28407
rect 4077 28169 4111 28203
rect 4905 28169 4939 28203
rect 8125 28169 8159 28203
rect 8953 28169 8987 28203
rect 10241 28169 10275 28203
rect 5917 28101 5951 28135
rect 6561 28101 6595 28135
rect 1777 28033 1811 28067
rect 2053 28033 2087 28067
rect 2605 28033 2639 28067
rect 4905 28033 4939 28067
rect 4997 28033 5031 28067
rect 5733 28033 5767 28067
rect 6745 28033 6779 28067
rect 7757 28033 7791 28067
rect 8585 28033 8619 28067
rect 10241 28033 10275 28067
rect 10977 28033 11011 28067
rect 11989 28033 12023 28067
rect 13001 28033 13035 28067
rect 13185 28033 13219 28067
rect 15200 28033 15234 28067
rect 2145 27965 2179 27999
rect 9873 27965 9907 27999
rect 11713 27965 11747 27999
rect 14933 27965 14967 27999
rect 8125 27897 8159 27931
rect 8953 27897 8987 27931
rect 11069 27897 11103 27931
rect 6929 27829 6963 27863
rect 13001 27829 13035 27863
rect 16313 27829 16347 27863
rect 10609 27625 10643 27659
rect 11437 27625 11471 27659
rect 6009 27557 6043 27591
rect 9275 27557 9309 27591
rect 7021 27489 7055 27523
rect 7757 27489 7791 27523
rect 10241 27489 10275 27523
rect 11069 27489 11103 27523
rect 11437 27489 11471 27523
rect 11989 27489 12023 27523
rect 1961 27421 1995 27455
rect 2228 27421 2262 27455
rect 4077 27421 4111 27455
rect 6929 27421 6963 27455
rect 7113 27421 7147 27455
rect 7481 27421 7515 27455
rect 8217 27421 8251 27455
rect 8401 27421 8435 27455
rect 9172 27421 9206 27455
rect 10609 27421 10643 27455
rect 11897 27421 11931 27455
rect 12081 27421 12115 27455
rect 18061 27421 18095 27455
rect 18429 27421 18463 27455
rect 20729 27421 20763 27455
rect 4721 27353 4755 27387
rect 20974 27353 21008 27387
rect 3341 27285 3375 27319
rect 4261 27285 4295 27319
rect 14289 27285 14323 27319
rect 18429 27285 18463 27319
rect 22109 27285 22143 27319
rect 1961 27081 1995 27115
rect 2237 27081 2271 27115
rect 11713 27081 11747 27115
rect 13553 27081 13587 27115
rect 14381 27081 14415 27115
rect 2789 26945 2823 26979
rect 3056 26945 3090 26979
rect 4813 26945 4847 26979
rect 4997 26945 5031 26979
rect 5273 26945 5307 26979
rect 5549 26945 5583 26979
rect 6561 26945 6595 26979
rect 6745 26945 6779 26979
rect 7389 26945 7423 26979
rect 7573 26945 7607 26979
rect 8033 26945 8067 26979
rect 8217 26945 8251 26979
rect 12081 26945 12115 26979
rect 13185 26945 13219 26979
rect 14013 26945 14047 26979
rect 14381 26945 14415 26979
rect 18337 26945 18371 26979
rect 19165 26945 19199 26979
rect 19432 26945 19466 26979
rect 23285 26945 23319 26979
rect 1593 26877 1627 26911
rect 1869 26877 1903 26911
rect 2053 26877 2087 26911
rect 4721 26877 4755 26911
rect 12173 26877 12207 26911
rect 12357 26877 12391 26911
rect 13553 26877 13587 26911
rect 23029 26877 23063 26911
rect 4169 26741 4203 26775
rect 6653 26741 6687 26775
rect 7389 26741 7423 26775
rect 20545 26741 20579 26775
rect 24409 26741 24443 26775
rect 7389 26537 7423 26571
rect 8585 26537 8619 26571
rect 9597 26537 9631 26571
rect 12725 26537 12759 26571
rect 13553 26537 13587 26571
rect 17601 26537 17635 26571
rect 26985 26537 27019 26571
rect 5365 26469 5399 26503
rect 3985 26401 4019 26435
rect 6929 26401 6963 26435
rect 8217 26401 8251 26435
rect 10149 26401 10183 26435
rect 12357 26401 12391 26435
rect 13185 26401 13219 26435
rect 21833 26401 21867 26435
rect 1593 26333 1627 26367
rect 4252 26333 4286 26367
rect 5825 26333 5859 26367
rect 6009 26333 6043 26367
rect 6561 26333 6595 26367
rect 7573 26333 7607 26367
rect 8585 26333 8619 26367
rect 9965 26333 9999 26367
rect 12725 26333 12759 26367
rect 13553 26333 13587 26367
rect 16221 26333 16255 26367
rect 25605 26333 25639 26367
rect 5917 26265 5951 26299
rect 6745 26265 6779 26299
rect 16488 26265 16522 26299
rect 22100 26265 22134 26299
rect 25850 26265 25884 26299
rect 2881 26197 2915 26231
rect 10057 26197 10091 26231
rect 23213 26197 23247 26231
rect 4427 25993 4461 26027
rect 4905 25993 4939 26027
rect 6837 25993 6871 26027
rect 6929 25993 6963 26027
rect 8953 25993 8987 26027
rect 13553 25993 13587 26027
rect 26617 25993 26651 26027
rect 6561 25925 6595 25959
rect 10885 25925 10919 25959
rect 16221 25925 16255 25959
rect 18604 25925 18638 25959
rect 25504 25925 25538 25959
rect 1685 25857 1719 25891
rect 1869 25857 1903 25891
rect 1961 25857 1995 25891
rect 2677 25857 2711 25891
rect 5641 25857 5675 25891
rect 5733 25857 5767 25891
rect 6745 25857 6779 25891
rect 7113 25857 7147 25891
rect 8861 25857 8895 25891
rect 10701 25857 10735 25891
rect 10977 25857 11011 25891
rect 12265 25857 12299 25891
rect 13185 25857 13219 25891
rect 16037 25857 16071 25891
rect 16313 25857 16347 25891
rect 18337 25857 18371 25891
rect 2421 25789 2455 25823
rect 4813 25789 4847 25823
rect 4997 25789 5031 25823
rect 10517 25789 10551 25823
rect 25237 25789 25271 25823
rect 5825 25721 5859 25755
rect 13553 25721 13587 25755
rect 3801 25653 3835 25687
rect 12357 25653 12391 25687
rect 15853 25653 15887 25687
rect 19717 25653 19751 25687
rect 4077 25449 4111 25483
rect 6101 25449 6135 25483
rect 6285 25449 6319 25483
rect 7573 25449 7607 25483
rect 8401 25449 8435 25483
rect 11621 25449 11655 25483
rect 25329 25449 25363 25483
rect 25973 25449 26007 25483
rect 7757 25381 7791 25415
rect 9137 25381 9171 25415
rect 4629 25313 4663 25347
rect 5733 25313 5767 25347
rect 9689 25313 9723 25347
rect 12265 25313 12299 25347
rect 2053 25245 2087 25279
rect 2320 25245 2354 25279
rect 4353 25245 4387 25279
rect 8309 25245 8343 25279
rect 11805 25245 11839 25279
rect 11989 25245 12023 25279
rect 12817 25245 12851 25279
rect 13001 25245 13035 25279
rect 25881 25245 25915 25279
rect 26985 25245 27019 25279
rect 4537 25177 4571 25211
rect 6101 25177 6135 25211
rect 7389 25177 7423 25211
rect 7573 25177 7607 25211
rect 9505 25177 9539 25211
rect 11897 25177 11931 25211
rect 12107 25177 12141 25211
rect 13185 25177 13219 25211
rect 25697 25177 25731 25211
rect 27252 25177 27286 25211
rect 3433 25109 3467 25143
rect 9597 25109 9631 25143
rect 28365 25109 28399 25143
rect 5457 24905 5491 24939
rect 10241 24905 10275 24939
rect 11897 24905 11931 24939
rect 3157 24837 3191 24871
rect 2012 24769 2046 24803
rect 2973 24769 3007 24803
rect 3801 24769 3835 24803
rect 3985 24769 4019 24803
rect 4445 24769 4479 24803
rect 4629 24769 4663 24803
rect 5365 24769 5399 24803
rect 5549 24769 5583 24803
rect 10241 24769 10275 24803
rect 11897 24769 11931 24803
rect 12265 24769 12299 24803
rect 12909 24769 12943 24803
rect 13093 24769 13127 24803
rect 13185 24769 13219 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 16865 24769 16899 24803
rect 17049 24769 17083 24803
rect 17233 24769 17267 24803
rect 2099 24701 2133 24735
rect 3249 24701 3283 24735
rect 10057 24701 10091 24735
rect 10609 24701 10643 24735
rect 11713 24701 11747 24735
rect 2697 24633 2731 24667
rect 14381 24633 14415 24667
rect 12725 24565 12759 24599
rect 2927 24361 2961 24395
rect 10241 24361 10275 24395
rect 16589 24361 16623 24395
rect 5181 24293 5215 24327
rect 11621 24225 11655 24259
rect 21005 24225 21039 24259
rect 1777 24157 1811 24191
rect 2033 24157 2067 24191
rect 2329 24157 2363 24191
rect 2824 24157 2858 24191
rect 4537 24157 4571 24191
rect 4905 24157 4939 24191
rect 5273 24157 5307 24191
rect 6561 24157 6595 24191
rect 10149 24157 10183 24191
rect 11253 24157 11287 24191
rect 11529 24157 11563 24191
rect 12541 24157 12575 24191
rect 12817 24157 12851 24191
rect 16497 24157 16531 24191
rect 16681 24157 16715 24191
rect 26985 24157 27019 24191
rect 1593 24089 1627 24123
rect 6377 24089 6411 24123
rect 12357 24089 12391 24123
rect 12725 24089 12759 24123
rect 21250 24089 21284 24123
rect 27252 24089 27286 24123
rect 2145 24021 2179 24055
rect 2237 24021 2271 24055
rect 6745 24021 6779 24055
rect 22385 24021 22419 24055
rect 28365 24021 28399 24055
rect 4077 23817 4111 23851
rect 6761 23817 6795 23851
rect 7849 23817 7883 23851
rect 9873 23817 9907 23851
rect 2605 23749 2639 23783
rect 4813 23749 4847 23783
rect 6561 23749 6595 23783
rect 7481 23749 7515 23783
rect 25022 23749 25056 23783
rect 5089 23681 5123 23715
rect 5181 23681 5215 23715
rect 5273 23681 5307 23715
rect 5457 23681 5491 23715
rect 7665 23681 7699 23715
rect 9873 23681 9907 23715
rect 11897 23681 11931 23715
rect 14565 23681 14599 23715
rect 14832 23681 14866 23715
rect 9689 23613 9723 23647
rect 10241 23613 10275 23647
rect 12173 23613 12207 23647
rect 24777 23613 24811 23647
rect 1777 23477 1811 23511
rect 6745 23477 6779 23511
rect 6929 23477 6963 23511
rect 15945 23477 15979 23511
rect 26157 23477 26191 23511
rect 11805 23273 11839 23307
rect 12541 23273 12575 23307
rect 10149 23205 10183 23239
rect 5641 23137 5675 23171
rect 5733 23137 5767 23171
rect 9781 23137 9815 23171
rect 25881 23137 25915 23171
rect 4905 23069 4939 23103
rect 5089 23069 5123 23103
rect 5273 23069 5307 23103
rect 9965 23069 9999 23103
rect 11529 23069 11563 23103
rect 12357 23069 12391 23103
rect 13277 23069 13311 23103
rect 17233 23069 17267 23103
rect 21281 23069 21315 23103
rect 4353 23001 4387 23035
rect 17500 23001 17534 23035
rect 26148 23001 26182 23035
rect 12817 22933 12851 22967
rect 13369 22933 13403 22967
rect 18613 22933 18647 22967
rect 21465 22933 21499 22967
rect 27261 22933 27295 22967
rect 11713 22729 11747 22763
rect 12081 22729 12115 22763
rect 21373 22729 21407 22763
rect 6929 22661 6963 22695
rect 7573 22661 7607 22695
rect 9956 22661 9990 22695
rect 24124 22661 24158 22695
rect 6745 22593 6779 22627
rect 7021 22593 7055 22627
rect 7481 22593 7515 22627
rect 7665 22593 7699 22627
rect 9689 22593 9723 22627
rect 11897 22593 11931 22627
rect 12173 22593 12207 22627
rect 12909 22593 12943 22627
rect 13176 22593 13210 22627
rect 19993 22593 20027 22627
rect 20249 22593 20283 22627
rect 22017 22593 22051 22627
rect 22284 22593 22318 22627
rect 23857 22593 23891 22627
rect 11069 22457 11103 22491
rect 6561 22389 6595 22423
rect 14289 22389 14323 22423
rect 23397 22389 23431 22423
rect 25237 22389 25271 22423
rect 7573 22185 7607 22219
rect 10977 22185 11011 22219
rect 10609 22117 10643 22151
rect 1961 22049 1995 22083
rect 6101 22049 6135 22083
rect 12081 22049 12115 22083
rect 24593 22049 24627 22083
rect 1685 21981 1719 22015
rect 1869 21981 1903 22015
rect 2145 21981 2179 22015
rect 2329 21981 2363 22015
rect 5181 21981 5215 22015
rect 6377 21981 6411 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 6745 21981 6779 22015
rect 12357 21981 12391 22015
rect 15669 21981 15703 22015
rect 16405 21981 16439 22015
rect 21557 21981 21591 22015
rect 26985 21981 27019 22015
rect 4997 21913 5031 21947
rect 5549 21913 5583 21947
rect 7205 21913 7239 21947
rect 7389 21913 7423 21947
rect 10977 21913 11011 21947
rect 16672 21913 16706 21947
rect 21802 21913 21836 21947
rect 24838 21913 24872 21947
rect 27230 21913 27264 21947
rect 5273 21845 5307 21879
rect 5365 21845 5399 21879
rect 11161 21845 11195 21879
rect 15853 21845 15887 21879
rect 17785 21845 17819 21879
rect 22937 21845 22971 21879
rect 25973 21845 26007 21879
rect 28365 21845 28399 21879
rect 4077 21641 4111 21675
rect 7205 21641 7239 21675
rect 9045 21641 9079 21675
rect 7932 21573 7966 21607
rect 12440 21573 12474 21607
rect 18512 21573 18546 21607
rect 3157 21505 3191 21539
rect 3985 21505 4019 21539
rect 6837 21505 6871 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 9772 21505 9806 21539
rect 12173 21505 12207 21539
rect 14013 21505 14047 21539
rect 14197 21505 14231 21539
rect 15577 21505 15611 21539
rect 15945 21505 15979 21539
rect 16221 21505 16255 21539
rect 18245 21505 18279 21539
rect 20352 21505 20386 21539
rect 23480 21505 23514 21539
rect 25237 21505 25271 21539
rect 25493 21505 25527 21539
rect 9505 21437 9539 21471
rect 15853 21437 15887 21471
rect 20085 21437 20119 21471
rect 23213 21437 23247 21471
rect 3341 21369 3375 21403
rect 10885 21301 10919 21335
rect 13553 21301 13587 21335
rect 14013 21301 14047 21335
rect 19625 21301 19659 21335
rect 21465 21301 21499 21335
rect 24593 21301 24627 21335
rect 26617 21301 26651 21335
rect 6469 21097 6503 21131
rect 7113 21029 7147 21063
rect 12725 21029 12759 21063
rect 14289 20961 14323 20995
rect 4905 20893 4939 20927
rect 5181 20893 5215 20927
rect 5365 20893 5399 20927
rect 7389 20893 7423 20927
rect 8585 20893 8619 20927
rect 11345 20893 11379 20927
rect 14473 20893 14507 20927
rect 15485 20893 15519 20927
rect 20637 20893 20671 20927
rect 20904 20893 20938 20927
rect 22477 20893 22511 20927
rect 26065 20893 26099 20927
rect 6285 20825 6319 20859
rect 6501 20825 6535 20859
rect 7113 20825 7147 20859
rect 8217 20825 8251 20859
rect 9597 20825 9631 20859
rect 9781 20825 9815 20859
rect 11612 20825 11646 20859
rect 15730 20825 15764 20859
rect 22722 20825 22756 20859
rect 26310 20825 26344 20859
rect 5089 20757 5123 20791
rect 6653 20757 6687 20791
rect 7297 20757 7331 20791
rect 9965 20757 9999 20791
rect 14657 20757 14691 20791
rect 16865 20757 16899 20791
rect 22017 20757 22051 20791
rect 23857 20757 23891 20791
rect 27445 20757 27479 20791
rect 5365 20553 5399 20587
rect 5733 20553 5767 20587
rect 7021 20553 7055 20587
rect 7389 20553 7423 20587
rect 10517 20553 10551 20587
rect 11713 20553 11747 20587
rect 16129 20553 16163 20587
rect 8401 20485 8435 20519
rect 11069 20485 11103 20519
rect 14350 20485 14384 20519
rect 4169 20417 4203 20451
rect 5549 20417 5583 20451
rect 5825 20417 5859 20451
rect 7205 20417 7239 20451
rect 7481 20417 7515 20451
rect 8217 20417 8251 20451
rect 9229 20417 9263 20451
rect 9505 20417 9539 20451
rect 10793 20417 10827 20451
rect 15945 20417 15979 20451
rect 16221 20417 16255 20451
rect 18409 20417 18443 20451
rect 20249 20417 20283 20451
rect 22017 20417 22051 20451
rect 22284 20417 22318 20451
rect 23857 20417 23891 20451
rect 24124 20417 24158 20451
rect 4261 20349 4295 20383
rect 10701 20349 10735 20383
rect 11161 20349 11195 20383
rect 11897 20349 11931 20383
rect 11989 20349 12023 20383
rect 12081 20349 12115 20383
rect 12173 20349 12207 20383
rect 14105 20349 14139 20383
rect 18153 20349 18187 20383
rect 19993 20349 20027 20383
rect 4537 20281 4571 20315
rect 9045 20281 9079 20315
rect 15945 20281 15979 20315
rect 4353 20213 4387 20247
rect 8585 20213 8619 20247
rect 9413 20213 9447 20247
rect 15485 20213 15519 20247
rect 19533 20213 19567 20247
rect 21373 20213 21407 20247
rect 23397 20213 23431 20247
rect 25237 20213 25271 20247
rect 5733 20009 5767 20043
rect 6745 20009 6779 20043
rect 6929 20009 6963 20043
rect 8309 20009 8343 20043
rect 10241 20009 10275 20043
rect 18153 20009 18187 20043
rect 22845 20009 22879 20043
rect 26617 20009 26651 20043
rect 5733 19873 5767 19907
rect 11069 19873 11103 19907
rect 16773 19873 16807 19907
rect 4169 19805 4203 19839
rect 4353 19805 4387 19839
rect 4905 19805 4939 19839
rect 4997 19805 5031 19839
rect 5641 19805 5675 19839
rect 8033 19805 8067 19839
rect 9689 19805 9723 19839
rect 10057 19805 10091 19839
rect 11253 19805 11287 19839
rect 20821 19805 20855 19839
rect 22661 19805 22695 19839
rect 25237 19805 25271 19839
rect 6561 19737 6595 19771
rect 9873 19737 9907 19771
rect 9965 19737 9999 19771
rect 11437 19737 11471 19771
rect 17018 19737 17052 19771
rect 21066 19737 21100 19771
rect 25504 19737 25538 19771
rect 4261 19669 4295 19703
rect 5181 19669 5215 19703
rect 6009 19669 6043 19703
rect 6761 19669 6795 19703
rect 11345 19669 11379 19703
rect 11621 19669 11655 19703
rect 22201 19669 22235 19703
rect 3249 19465 3283 19499
rect 8125 19465 8159 19499
rect 9873 19465 9907 19499
rect 10517 19465 10551 19499
rect 15117 19465 15151 19499
rect 15777 19465 15811 19499
rect 15945 19465 15979 19499
rect 17601 19465 17635 19499
rect 20285 19465 20319 19499
rect 23765 19465 23799 19499
rect 7205 19397 7239 19431
rect 9597 19397 9631 19431
rect 15577 19397 15611 19431
rect 17233 19397 17267 19431
rect 17433 19397 17467 19431
rect 20085 19397 20119 19431
rect 22652 19397 22686 19431
rect 3341 19329 3375 19363
rect 3525 19329 3559 19363
rect 4353 19329 4387 19363
rect 6561 19329 6595 19363
rect 6837 19329 6871 19363
rect 8493 19329 8527 19363
rect 10793 19329 10827 19363
rect 10885 19329 10919 19363
rect 10977 19329 11011 19363
rect 11161 19329 11195 19363
rect 12357 19329 12391 19363
rect 12817 19329 12851 19363
rect 13001 19329 13035 19363
rect 13737 19329 13771 19363
rect 13993 19329 14027 19363
rect 22385 19329 22419 19363
rect 25493 19329 25527 19363
rect 4629 19261 4663 19295
rect 7021 19261 7055 19295
rect 8309 19261 8343 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 25237 19261 25271 19295
rect 12817 19193 12851 19227
rect 3065 19125 3099 19159
rect 15761 19125 15795 19159
rect 17417 19125 17451 19159
rect 20269 19125 20303 19159
rect 20453 19125 20487 19159
rect 26617 19125 26651 19159
rect 4169 18921 4203 18955
rect 4353 18921 4387 18955
rect 6469 18921 6503 18955
rect 7021 18921 7055 18955
rect 8585 18921 8619 18955
rect 17325 18921 17359 18955
rect 19993 18921 20027 18955
rect 9137 18853 9171 18887
rect 14381 18853 14415 18887
rect 18061 18853 18095 18887
rect 22753 18853 22787 18887
rect 10241 18785 10275 18819
rect 16037 18785 16071 18819
rect 16681 18785 16715 18819
rect 18705 18785 18739 18819
rect 20177 18785 20211 18819
rect 23397 18785 23431 18819
rect 26249 18785 26283 18819
rect 5733 18717 5767 18751
rect 6009 18717 6043 18751
rect 6594 18717 6628 18751
rect 7113 18717 7147 18751
rect 7941 18717 7975 18751
rect 8034 18717 8068 18751
rect 8406 18717 8440 18751
rect 9321 18717 9355 18751
rect 9597 18717 9631 18751
rect 10057 18717 10091 18751
rect 11345 18717 11379 18751
rect 14841 18717 14875 18751
rect 16221 18717 16255 18751
rect 18245 18717 18279 18751
rect 18429 18717 18463 18751
rect 20085 18717 20119 18751
rect 20269 18717 20303 18751
rect 20453 18717 20487 18751
rect 20913 18717 20947 18751
rect 22937 18717 22971 18751
rect 23029 18717 23063 18751
rect 17371 18683 17405 18717
rect 3985 18649 4019 18683
rect 5549 18649 5583 18683
rect 8217 18649 8251 18683
rect 8309 18649 8343 18683
rect 10793 18649 10827 18683
rect 11612 18649 11646 18683
rect 14381 18649 14415 18683
rect 15117 18649 15151 18683
rect 16313 18649 16347 18683
rect 16405 18649 16439 18683
rect 16543 18649 16577 18683
rect 17141 18649 17175 18683
rect 18337 18649 18371 18683
rect 18547 18649 18581 18683
rect 21180 18649 21214 18683
rect 23121 18649 23155 18683
rect 23259 18649 23293 18683
rect 26494 18649 26528 18683
rect 4195 18581 4229 18615
rect 5917 18581 5951 18615
rect 6653 18581 6687 18615
rect 9505 18581 9539 18615
rect 10609 18581 10643 18615
rect 10701 18581 10735 18615
rect 12725 18581 12759 18615
rect 14933 18581 14967 18615
rect 17509 18581 17543 18615
rect 19717 18581 19751 18615
rect 22293 18581 22327 18615
rect 27629 18581 27663 18615
rect 5273 18377 5307 18411
rect 7297 18377 7331 18411
rect 10977 18377 11011 18411
rect 13553 18377 13587 18411
rect 22385 18377 22419 18411
rect 25421 18377 25455 18411
rect 6745 18309 6779 18343
rect 8953 18309 8987 18343
rect 13461 18309 13495 18343
rect 14718 18309 14752 18343
rect 17233 18309 17267 18343
rect 18429 18309 18463 18343
rect 22017 18309 22051 18343
rect 22217 18309 22251 18343
rect 23296 18309 23330 18343
rect 25053 18309 25087 18343
rect 25145 18309 25179 18343
rect 2973 18241 3007 18275
rect 3157 18241 3191 18275
rect 4261 18241 4295 18275
rect 4813 18241 4847 18275
rect 4997 18241 5031 18275
rect 6653 18241 6687 18275
rect 7573 18241 7607 18275
rect 7665 18241 7699 18275
rect 10333 18241 10367 18275
rect 10426 18241 10460 18275
rect 10609 18241 10643 18275
rect 10701 18241 10735 18275
rect 10839 18241 10873 18275
rect 14473 18241 14507 18275
rect 17049 18241 17083 18275
rect 17141 18241 17175 18275
rect 17351 18241 17385 18275
rect 18061 18241 18095 18275
rect 18154 18241 18188 18275
rect 18337 18241 18371 18275
rect 18567 18241 18601 18275
rect 19257 18241 19291 18275
rect 19349 18241 19383 18275
rect 24869 18241 24903 18275
rect 25237 18241 25271 18275
rect 7481 18173 7515 18207
rect 7757 18173 7791 18207
rect 17509 18173 17543 18207
rect 23029 18173 23063 18207
rect 3065 18037 3099 18071
rect 9229 18037 9263 18071
rect 15853 18037 15887 18071
rect 16865 18037 16899 18071
rect 18705 18037 18739 18071
rect 19533 18037 19567 18071
rect 22201 18037 22235 18071
rect 24409 18037 24443 18071
rect 2881 17833 2915 17867
rect 3341 17833 3375 17867
rect 5733 17833 5767 17867
rect 5917 17833 5951 17867
rect 7205 17833 7239 17867
rect 10149 17833 10183 17867
rect 12357 17833 12391 17867
rect 14289 17833 14323 17867
rect 18429 17833 18463 17867
rect 22937 17833 22971 17867
rect 6469 17765 6503 17799
rect 13737 17765 13771 17799
rect 20821 17765 20855 17799
rect 3065 17697 3099 17731
rect 4445 17697 4479 17731
rect 4537 17697 4571 17731
rect 11529 17697 11563 17731
rect 11805 17697 11839 17731
rect 13461 17697 13495 17731
rect 26985 17697 27019 17731
rect 2789 17629 2823 17663
rect 3985 17629 4019 17663
rect 6653 17629 6687 17663
rect 6745 17629 6779 17663
rect 7389 17629 7423 17663
rect 7481 17629 7515 17663
rect 7665 17629 7699 17663
rect 7757 17629 7791 17663
rect 8309 17629 8343 17663
rect 9965 17629 9999 17663
rect 10793 17629 10827 17663
rect 11069 17629 11103 17663
rect 11345 17629 11379 17663
rect 12633 17629 12667 17663
rect 13093 17629 13127 17663
rect 14473 17629 14507 17663
rect 14749 17629 14783 17663
rect 17049 17629 17083 17663
rect 19441 17629 19475 17663
rect 25053 17629 25087 17663
rect 5549 17561 5583 17595
rect 5733 17561 5767 17595
rect 6469 17561 6503 17595
rect 9321 17561 9355 17595
rect 9505 17561 9539 17595
rect 12357 17561 12391 17595
rect 13578 17561 13612 17595
rect 17294 17561 17328 17595
rect 19686 17561 19720 17595
rect 22753 17561 22787 17595
rect 25298 17561 25332 17595
rect 27230 17561 27264 17595
rect 4169 17493 4203 17527
rect 8493 17493 8527 17527
rect 12541 17493 12575 17527
rect 13369 17493 13403 17527
rect 14657 17493 14691 17527
rect 22953 17493 22987 17527
rect 23121 17493 23155 17527
rect 26433 17493 26467 17527
rect 28365 17493 28399 17527
rect 2697 17289 2731 17323
rect 3249 17289 3283 17323
rect 6009 17289 6043 17323
rect 8217 17289 8251 17323
rect 12265 17289 12299 17323
rect 12725 17289 12759 17323
rect 14841 17289 14875 17323
rect 19257 17289 19291 17323
rect 4629 17221 4663 17255
rect 5549 17221 5583 17255
rect 8125 17221 8159 17255
rect 9220 17221 9254 17255
rect 11897 17221 11931 17255
rect 13093 17221 13127 17255
rect 15025 17221 15059 17255
rect 18061 17221 18095 17255
rect 18261 17221 18295 17255
rect 18889 17221 18923 17255
rect 19089 17221 19123 17255
rect 20269 17221 20303 17255
rect 25504 17221 25538 17255
rect 1685 17153 1719 17187
rect 2513 17153 2547 17187
rect 2789 17153 2823 17187
rect 3433 17153 3467 17187
rect 3526 17153 3560 17187
rect 3801 17153 3835 17187
rect 4261 17153 4295 17187
rect 4445 17153 4479 17187
rect 5825 17153 5859 17187
rect 6561 17153 6595 17187
rect 6929 17153 6963 17187
rect 7205 17153 7239 17187
rect 10793 17153 10827 17187
rect 12081 17153 12115 17187
rect 12909 17153 12943 17187
rect 13185 17153 13219 17187
rect 20177 17153 20211 17187
rect 20361 17153 20395 17187
rect 20479 17153 20513 17187
rect 20637 17153 20671 17187
rect 21281 17153 21315 17187
rect 22284 17153 22318 17187
rect 25237 17153 25271 17187
rect 1777 17085 1811 17119
rect 5733 17085 5767 17119
rect 7297 17085 7331 17119
rect 7573 17085 7607 17119
rect 8953 17085 8987 17119
rect 14565 17085 14599 17119
rect 14933 17085 14967 17119
rect 21097 17085 21131 17119
rect 22017 17085 22051 17119
rect 3709 17017 3743 17051
rect 10333 17017 10367 17051
rect 18429 17017 18463 17051
rect 2329 16949 2363 16983
rect 5549 16949 5583 16983
rect 10977 16949 11011 16983
rect 15209 16949 15243 16983
rect 18245 16949 18279 16983
rect 19073 16949 19107 16983
rect 19993 16949 20027 16983
rect 21465 16949 21499 16983
rect 23397 16949 23431 16983
rect 26617 16949 26651 16983
rect 1777 16745 1811 16779
rect 5825 16745 5859 16779
rect 6009 16745 6043 16779
rect 20821 16745 20855 16779
rect 7297 16677 7331 16711
rect 9505 16677 9539 16711
rect 20177 16677 20211 16711
rect 23857 16677 23891 16711
rect 2697 16609 2731 16643
rect 4353 16609 4387 16643
rect 11529 16609 11563 16643
rect 15025 16609 15059 16643
rect 17877 16609 17911 16643
rect 18245 16609 18279 16643
rect 20913 16609 20947 16643
rect 26985 16609 27019 16643
rect 1593 16541 1627 16575
rect 2421 16541 2455 16575
rect 3341 16541 3375 16575
rect 3433 16541 3467 16575
rect 4629 16541 4663 16575
rect 4813 16541 4847 16575
rect 6469 16541 6503 16575
rect 7481 16541 7515 16575
rect 8585 16541 8619 16575
rect 9229 16541 9263 16575
rect 9505 16541 9539 16575
rect 9689 16541 9723 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 11069 16541 11103 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 16865 16541 16899 16575
rect 17049 16541 17083 16575
rect 18061 16541 18095 16575
rect 19540 16541 19574 16575
rect 19626 16541 19660 16575
rect 20039 16541 20073 16575
rect 21097 16541 21131 16575
rect 22293 16541 22327 16575
rect 22477 16541 22511 16575
rect 22569 16541 22603 16575
rect 22661 16541 22695 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 24593 16541 24627 16575
rect 3157 16473 3191 16507
rect 5641 16473 5675 16507
rect 8309 16473 8343 16507
rect 15292 16473 15326 16507
rect 19809 16473 19843 16507
rect 19901 16473 19935 16507
rect 20821 16473 20855 16507
rect 23581 16473 23615 16507
rect 24860 16473 24894 16507
rect 27230 16473 27264 16507
rect 3255 16405 3289 16439
rect 4537 16405 4571 16439
rect 5841 16405 5875 16439
rect 6653 16405 6687 16439
rect 8407 16405 8441 16439
rect 8493 16405 8527 16439
rect 16405 16405 16439 16439
rect 17233 16405 17267 16439
rect 21281 16405 21315 16439
rect 22845 16405 22879 16439
rect 25973 16405 26007 16439
rect 28365 16405 28399 16439
rect 3893 16201 3927 16235
rect 4813 16201 4847 16235
rect 5917 16201 5951 16235
rect 8493 16201 8527 16235
rect 9321 16133 9355 16167
rect 9413 16133 9447 16167
rect 11805 16133 11839 16167
rect 14289 16133 14323 16167
rect 15669 16133 15703 16167
rect 19257 16133 19291 16167
rect 19350 16133 19384 16167
rect 20085 16133 20119 16167
rect 20285 16133 20319 16167
rect 20913 16133 20947 16167
rect 21113 16133 21147 16167
rect 25504 16133 25538 16167
rect 15899 16099 15933 16133
rect 1869 16065 1903 16099
rect 2605 16065 2639 16099
rect 4997 16065 5031 16099
rect 5089 16065 5123 16099
rect 5273 16065 5307 16099
rect 5365 16065 5399 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6561 16065 6595 16099
rect 6709 16065 6743 16099
rect 6837 16065 6871 16099
rect 6929 16065 6963 16099
rect 7067 16065 7101 16099
rect 8309 16065 8343 16099
rect 9229 16065 9263 16099
rect 9689 16065 9723 16099
rect 10149 16065 10183 16099
rect 10425 16065 10459 16099
rect 10701 16065 10735 16099
rect 11713 16065 11747 16099
rect 11897 16065 11931 16099
rect 12449 16065 12483 16099
rect 12716 16065 12750 16099
rect 14473 16065 14507 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 17693 16065 17727 16099
rect 19166 16055 19200 16089
rect 19467 16065 19501 16099
rect 19625 16065 19659 16099
rect 22017 16065 22051 16099
rect 22273 16065 22307 16099
rect 23857 16065 23891 16099
rect 25237 16065 25271 16099
rect 8125 15997 8159 16031
rect 10885 15997 10919 16031
rect 17509 15997 17543 16031
rect 2053 15929 2087 15963
rect 9597 15929 9631 15963
rect 11161 15929 11195 15963
rect 20453 15929 20487 15963
rect 7205 15861 7239 15895
rect 8953 15861 8987 15895
rect 13829 15861 13863 15895
rect 15853 15861 15887 15895
rect 16037 15861 16071 15895
rect 17877 15861 17911 15895
rect 18981 15861 19015 15895
rect 20269 15861 20303 15895
rect 21097 15861 21131 15895
rect 21281 15861 21315 15895
rect 23397 15861 23431 15895
rect 24041 15861 24075 15895
rect 26617 15861 26651 15895
rect 2881 15657 2915 15691
rect 4169 15657 4203 15691
rect 5549 15657 5583 15691
rect 8309 15657 8343 15691
rect 10149 15657 10183 15691
rect 12725 15657 12759 15691
rect 16773 15657 16807 15691
rect 16957 15657 16991 15691
rect 20821 15657 20855 15691
rect 22385 15657 22419 15691
rect 1961 15589 1995 15623
rect 4353 15589 4387 15623
rect 9597 15589 9631 15623
rect 14381 15589 14415 15623
rect 5733 15521 5767 15555
rect 10333 15521 10367 15555
rect 19441 15521 19475 15555
rect 21925 15521 21959 15555
rect 23029 15521 23063 15555
rect 24593 15521 24627 15555
rect 1777 15453 1811 15487
rect 2513 15453 2547 15487
rect 5457 15453 5491 15487
rect 6469 15453 6503 15487
rect 6561 15453 6595 15487
rect 6745 15453 6779 15487
rect 6837 15453 6871 15487
rect 7665 15453 7699 15487
rect 7813 15453 7847 15487
rect 8171 15453 8205 15487
rect 9413 15453 9447 15487
rect 10425 15453 10459 15487
rect 11345 15453 11379 15487
rect 11601 15453 11635 15487
rect 14933 15453 14967 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16865 15453 16899 15487
rect 17049 15453 17083 15487
rect 17233 15453 17267 15487
rect 17693 15453 17727 15487
rect 17786 15453 17820 15487
rect 18158 15453 18192 15487
rect 21465 15453 21499 15487
rect 21557 15453 21591 15487
rect 22569 15453 22603 15487
rect 22661 15453 22695 15487
rect 26985 15453 27019 15487
rect 3985 15385 4019 15419
rect 4185 15385 4219 15419
rect 6285 15385 6319 15419
rect 7941 15385 7975 15419
rect 8033 15385 8067 15419
rect 10149 15385 10183 15419
rect 14381 15385 14415 15419
rect 15945 15385 15979 15419
rect 17969 15385 18003 15419
rect 18061 15385 18095 15419
rect 19708 15385 19742 15419
rect 21281 15385 21315 15419
rect 21649 15385 21683 15419
rect 21767 15385 21801 15419
rect 22753 15385 22787 15419
rect 22891 15385 22925 15419
rect 23581 15385 23615 15419
rect 23765 15385 23799 15419
rect 24860 15385 24894 15419
rect 27230 15385 27264 15419
rect 2881 15317 2915 15351
rect 3065 15317 3099 15351
rect 5733 15317 5767 15351
rect 10609 15317 10643 15351
rect 14841 15317 14875 15351
rect 15117 15317 15151 15351
rect 16497 15317 16531 15351
rect 18337 15317 18371 15351
rect 25973 15317 26007 15351
rect 28365 15317 28399 15351
rect 2253 15113 2287 15147
rect 6561 15113 6595 15147
rect 10793 15113 10827 15147
rect 11897 15113 11931 15147
rect 17065 15113 17099 15147
rect 22585 15113 22619 15147
rect 2053 15045 2087 15079
rect 9413 15045 9447 15079
rect 14994 15045 15028 15079
rect 16865 15045 16899 15079
rect 18705 15045 18739 15079
rect 20076 15045 20110 15079
rect 22385 15045 22419 15079
rect 23857 15045 23891 15079
rect 23949 15045 23983 15079
rect 25504 15045 25538 15079
rect 2881 14977 2915 15011
rect 5089 14977 5123 15011
rect 6837 14977 6871 15011
rect 7757 14977 7791 15011
rect 7941 14977 7975 15011
rect 8033 14977 8067 15011
rect 8696 14977 8730 15011
rect 8861 14977 8895 15011
rect 8953 14977 8987 15011
rect 9597 14977 9631 15011
rect 9689 14977 9723 15011
rect 10149 14977 10183 15011
rect 10242 14977 10276 15011
rect 10425 14977 10459 15011
rect 10517 14977 10551 15011
rect 10655 14977 10689 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 14749 14977 14783 15011
rect 17877 14977 17911 15011
rect 23581 14977 23615 15011
rect 23729 14977 23763 15011
rect 24087 14977 24121 15011
rect 25237 14977 25271 15011
rect 5181 14909 5215 14943
rect 6745 14909 6779 14943
rect 6929 14909 6963 14943
rect 7021 14909 7055 14943
rect 7573 14909 7607 14943
rect 9485 14909 9519 14943
rect 17693 14909 17727 14943
rect 19809 14909 19843 14943
rect 5457 14841 5491 14875
rect 18061 14841 18095 14875
rect 24225 14841 24259 14875
rect 2237 14773 2271 14807
rect 2421 14773 2455 14807
rect 4169 14773 4203 14807
rect 5089 14773 5123 14807
rect 8493 14773 8527 14807
rect 16129 14773 16163 14807
rect 17049 14773 17083 14807
rect 17233 14773 17267 14807
rect 18797 14773 18831 14807
rect 21189 14773 21223 14807
rect 22569 14773 22603 14807
rect 22753 14773 22787 14807
rect 26617 14773 26651 14807
rect 1777 14569 1811 14603
rect 3433 14569 3467 14603
rect 4353 14569 4387 14603
rect 5549 14569 5583 14603
rect 7849 14569 7883 14603
rect 11713 14569 11747 14603
rect 12541 14569 12575 14603
rect 16957 14569 16991 14603
rect 17785 14569 17819 14603
rect 17877 14569 17911 14603
rect 9137 14501 9171 14535
rect 17693 14501 17727 14535
rect 18797 14501 18831 14535
rect 19717 14501 19751 14535
rect 23765 14501 23799 14535
rect 2881 14433 2915 14467
rect 3985 14433 4019 14467
rect 14749 14433 14783 14467
rect 26985 14433 27019 14467
rect 1593 14365 1627 14399
rect 3249 14365 3283 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 6009 14365 6043 14399
rect 6101 14365 6135 14399
rect 6929 14365 6963 14399
rect 7205 14365 7239 14399
rect 7389 14365 7423 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 8401 14365 8435 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9413 14365 9447 14399
rect 9505 14365 9539 14399
rect 9625 14365 9659 14399
rect 11069 14365 11103 14399
rect 11217 14365 11251 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 11573 14365 11607 14399
rect 12817 14365 12851 14399
rect 14565 14365 14599 14399
rect 15577 14365 15611 14399
rect 18153 14365 18187 14399
rect 18613 14365 18647 14399
rect 21465 14365 21499 14399
rect 21649 14365 21683 14399
rect 22385 14365 22419 14399
rect 25145 14365 25179 14399
rect 25513 14365 25547 14399
rect 4353 14297 4387 14331
rect 12541 14297 12575 14331
rect 14289 14297 14323 14331
rect 15844 14297 15878 14331
rect 19533 14297 19567 14331
rect 22652 14297 22686 14331
rect 25329 14297 25363 14331
rect 25421 14297 25455 14331
rect 27230 14297 27264 14331
rect 3065 14229 3099 14263
rect 4537 14229 4571 14263
rect 6745 14229 6779 14263
rect 12725 14229 12759 14263
rect 14657 14229 14691 14263
rect 14933 14229 14967 14263
rect 17417 14229 17451 14263
rect 18061 14229 18095 14263
rect 21833 14229 21867 14263
rect 25697 14229 25731 14263
rect 28365 14229 28399 14263
rect 4721 14025 4755 14059
rect 6009 14025 6043 14059
rect 10977 14025 11011 14059
rect 13093 14025 13127 14059
rect 16313 14025 16347 14059
rect 18245 14025 18279 14059
rect 20821 14025 20855 14059
rect 22385 14025 22419 14059
rect 25513 14025 25547 14059
rect 26525 14025 26559 14059
rect 8401 13957 8435 13991
rect 9864 13957 9898 13991
rect 13553 13957 13587 13991
rect 13769 13957 13803 13991
rect 14958 13957 14992 13991
rect 15945 13957 15979 13991
rect 16161 13957 16195 13991
rect 22017 13957 22051 13991
rect 22217 13957 22251 13991
rect 23305 13957 23339 13991
rect 26157 13957 26191 13991
rect 26249 13957 26283 13991
rect 23535 13923 23569 13957
rect 3525 13889 3559 13923
rect 5089 13889 5123 13923
rect 5733 13889 5767 13923
rect 7113 13889 7147 13923
rect 8125 13889 8159 13923
rect 8309 13889 8343 13923
rect 8545 13889 8579 13923
rect 11980 13889 12014 13923
rect 18061 13889 18095 13923
rect 18337 13889 18371 13923
rect 18797 13889 18831 13923
rect 19064 13889 19098 13923
rect 20637 13889 20671 13923
rect 24133 13889 24167 13923
rect 24389 13889 24423 13923
rect 25973 13889 26007 13923
rect 26341 13889 26375 13923
rect 4905 13821 4939 13855
rect 4997 13821 5031 13855
rect 5181 13821 5215 13855
rect 6009 13821 6043 13855
rect 9597 13821 9631 13855
rect 11713 13821 11747 13855
rect 14473 13821 14507 13855
rect 14749 13821 14783 13855
rect 14841 13821 14875 13855
rect 5825 13753 5859 13787
rect 7297 13753 7331 13787
rect 8677 13753 8711 13787
rect 15117 13753 15151 13787
rect 17877 13753 17911 13787
rect 3709 13685 3743 13719
rect 13737 13685 13771 13719
rect 13921 13685 13955 13719
rect 16129 13685 16163 13719
rect 17601 13685 17635 13719
rect 17969 13685 18003 13719
rect 20177 13685 20211 13719
rect 22201 13685 22235 13719
rect 23489 13685 23523 13719
rect 23673 13685 23707 13719
rect 3985 13481 4019 13515
rect 6653 13481 6687 13515
rect 10609 13481 10643 13515
rect 14473 13481 14507 13515
rect 16313 13481 16347 13515
rect 16497 13481 16531 13515
rect 17693 13481 17727 13515
rect 23673 13481 23707 13515
rect 26065 13481 26099 13515
rect 5641 13413 5675 13447
rect 9413 13413 9447 13447
rect 15117 13413 15151 13447
rect 23765 13413 23799 13447
rect 4629 13345 4663 13379
rect 5825 13345 5859 13379
rect 6837 13345 6871 13379
rect 6929 13345 6963 13379
rect 11437 13345 11471 13379
rect 15669 13345 15703 13379
rect 26525 13345 26559 13379
rect 4261 13277 4295 13311
rect 4721 13277 4755 13311
rect 5917 13277 5951 13311
rect 6009 13277 6043 13311
rect 6101 13277 6135 13311
rect 7021 13277 7055 13311
rect 7113 13277 7147 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 8401 13277 8435 13311
rect 8585 13277 8619 13311
rect 9597 13277 9631 13311
rect 9689 13277 9723 13311
rect 10885 13277 10919 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 15301 13277 15335 13311
rect 17509 13277 17543 13311
rect 17601 13277 17635 13311
rect 17969 13277 18003 13311
rect 19533 13277 19567 13311
rect 21005 13277 21039 13311
rect 23581 13277 23615 13311
rect 24041 13277 24075 13311
rect 24685 13277 24719 13311
rect 4445 13209 4479 13243
rect 9413 13209 9447 13243
rect 10609 13209 10643 13243
rect 12173 13209 12207 13243
rect 14289 13209 14323 13243
rect 15393 13209 15427 13243
rect 16129 13209 16163 13243
rect 21250 13209 21284 13243
rect 24952 13209 24986 13243
rect 26792 13209 26826 13243
rect 4353 13141 4387 13175
rect 8493 13141 8527 13175
rect 10793 13141 10827 13175
rect 11621 13141 11655 13175
rect 14489 13141 14523 13175
rect 14657 13141 14691 13175
rect 15485 13141 15519 13175
rect 16329 13141 16363 13175
rect 17233 13141 17267 13175
rect 17877 13141 17911 13175
rect 19625 13141 19659 13175
rect 22385 13141 22419 13175
rect 23305 13141 23339 13175
rect 23949 13141 23983 13175
rect 27905 13141 27939 13175
rect 4721 12937 4755 12971
rect 5917 12937 5951 12971
rect 7941 12937 7975 12971
rect 13093 12937 13127 12971
rect 13921 12937 13955 12971
rect 14289 12937 14323 12971
rect 18153 12937 18187 12971
rect 18889 12937 18923 12971
rect 6653 12869 6687 12903
rect 6853 12869 6887 12903
rect 12541 12869 12575 12903
rect 14105 12869 14139 12903
rect 15945 12869 15979 12903
rect 17785 12869 17819 12903
rect 18001 12869 18035 12903
rect 19441 12869 19475 12903
rect 22661 12869 22695 12903
rect 4905 12801 4939 12835
rect 5641 12801 5675 12835
rect 7665 12801 7699 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 9045 12801 9079 12835
rect 9781 12801 9815 12835
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 15669 12801 15703 12835
rect 15817 12801 15851 12835
rect 16037 12801 16071 12835
rect 16134 12801 16168 12835
rect 17049 12801 17083 12835
rect 18705 12801 18739 12835
rect 19717 12801 19751 12835
rect 22293 12801 22327 12835
rect 22386 12801 22420 12835
rect 22569 12801 22603 12835
rect 22758 12801 22792 12835
rect 24041 12801 24075 12835
rect 24133 12801 24167 12835
rect 24317 12801 24351 12835
rect 25044 12801 25078 12835
rect 5181 12733 5215 12767
rect 5917 12733 5951 12767
rect 7941 12733 7975 12767
rect 13001 12733 13035 12767
rect 16865 12733 16899 12767
rect 19533 12733 19567 12767
rect 23581 12733 23615 12767
rect 23949 12733 23983 12767
rect 24777 12733 24811 12767
rect 7757 12665 7791 12699
rect 12541 12665 12575 12699
rect 23857 12665 23891 12699
rect 5089 12597 5123 12631
rect 5733 12597 5767 12631
rect 6837 12597 6871 12631
rect 7021 12597 7055 12631
rect 8493 12597 8527 12631
rect 9229 12597 9263 12631
rect 9873 12597 9907 12631
rect 13277 12597 13311 12631
rect 16313 12597 16347 12631
rect 17233 12597 17267 12631
rect 17969 12597 18003 12631
rect 19717 12597 19751 12631
rect 19901 12597 19935 12631
rect 22937 12597 22971 12631
rect 26157 12597 26191 12631
rect 3985 12393 4019 12427
rect 5273 12393 5307 12427
rect 5457 12393 5491 12427
rect 6377 12393 6411 12427
rect 7481 12393 7515 12427
rect 12081 12393 12115 12427
rect 17049 12393 17083 12427
rect 17141 12393 17175 12427
rect 19625 12393 19659 12427
rect 21465 12393 21499 12427
rect 23489 12393 23523 12427
rect 23673 12393 23707 12427
rect 9689 12325 9723 12359
rect 20637 12325 20671 12359
rect 1869 12257 1903 12291
rect 8493 12257 8527 12291
rect 10241 12257 10275 12291
rect 18337 12257 18371 12291
rect 20269 12257 20303 12291
rect 21097 12257 21131 12291
rect 1593 12189 1627 12223
rect 4169 12189 4203 12223
rect 4353 12189 4387 12223
rect 4445 12189 4479 12223
rect 4905 12189 4939 12223
rect 5273 12189 5307 12223
rect 6653 12189 6687 12223
rect 6745 12189 6779 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 7481 12189 7515 12223
rect 7665 12189 7699 12223
rect 8309 12189 8343 12223
rect 8585 12189 8619 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 14289 12189 14323 12223
rect 17233 12189 17267 12223
rect 17509 12189 17543 12223
rect 18061 12189 18095 12223
rect 18153 12189 18187 12223
rect 20453 12189 20487 12223
rect 21281 12189 21315 12223
rect 22201 12189 22235 12223
rect 22349 12189 22383 12223
rect 22477 12189 22511 12223
rect 22569 12189 22603 12223
rect 22666 12189 22700 12223
rect 25145 12189 25179 12223
rect 26985 12189 27019 12223
rect 19671 12155 19705 12189
rect 9689 12121 9723 12155
rect 14556 12121 14590 12155
rect 19441 12121 19475 12155
rect 23305 12121 23339 12155
rect 23505 12121 23539 12155
rect 25412 12121 25446 12155
rect 27230 12121 27264 12155
rect 8125 12053 8159 12087
rect 10149 12053 10183 12087
rect 10425 12053 10459 12087
rect 15669 12053 15703 12087
rect 16773 12053 16807 12087
rect 17417 12053 17451 12087
rect 19809 12053 19843 12087
rect 22845 12053 22879 12087
rect 26525 12053 26559 12087
rect 28365 12053 28399 12087
rect 6009 11849 6043 11883
rect 6929 11849 6963 11883
rect 8217 11849 8251 11883
rect 15577 11849 15611 11883
rect 25053 11849 25087 11883
rect 4261 11781 4295 11815
rect 6561 11781 6595 11815
rect 6745 11781 6779 11815
rect 9772 11781 9806 11815
rect 15209 11781 15243 11815
rect 19901 11781 19935 11815
rect 22845 11781 22879 11815
rect 22937 11781 22971 11815
rect 23940 11781 23974 11815
rect 25789 11781 25823 11815
rect 27445 11781 27479 11815
rect 3893 11713 3927 11747
rect 5181 11713 5215 11747
rect 5825 11713 5859 11747
rect 6009 11713 6043 11747
rect 8309 11713 8343 11747
rect 9505 11713 9539 11747
rect 11969 11713 12003 11747
rect 14197 11713 14231 11747
rect 14381 11713 14415 11747
rect 15025 11713 15059 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 16865 11713 16899 11747
rect 17693 11713 17727 11747
rect 17960 11713 17994 11747
rect 19533 11713 19567 11747
rect 19626 11713 19660 11747
rect 19809 11713 19843 11747
rect 19998 11713 20032 11747
rect 21097 11713 21131 11747
rect 21281 11713 21315 11747
rect 22661 11713 22695 11747
rect 23029 11713 23063 11747
rect 25513 11713 25547 11747
rect 25697 11713 25731 11747
rect 25881 11713 25915 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 27537 11713 27571 11747
rect 4997 11645 5031 11679
rect 5089 11645 5123 11679
rect 5273 11645 5307 11679
rect 8401 11645 8435 11679
rect 11713 11645 11747 11679
rect 23673 11645 23707 11679
rect 7849 11577 7883 11611
rect 14473 11577 14507 11611
rect 4813 11509 4847 11543
rect 10885 11509 10919 11543
rect 13093 11509 13127 11543
rect 17049 11509 17083 11543
rect 19073 11509 19107 11543
rect 20177 11509 20211 11543
rect 21465 11509 21499 11543
rect 23213 11509 23247 11543
rect 26065 11509 26099 11543
rect 27721 11509 27755 11543
rect 4077 11305 4111 11339
rect 5917 11305 5951 11339
rect 6837 11305 6871 11339
rect 9873 11305 9907 11339
rect 15761 11305 15795 11339
rect 15945 11305 15979 11339
rect 20361 11305 20395 11339
rect 25145 11305 25179 11339
rect 4629 11237 4663 11271
rect 7021 11237 7055 11271
rect 7665 11237 7699 11271
rect 9321 11237 9355 11271
rect 11805 11237 11839 11271
rect 18889 11237 18923 11271
rect 24041 11237 24075 11271
rect 27353 11237 27387 11271
rect 5365 11169 5399 11203
rect 9965 11169 9999 11203
rect 10425 11169 10459 11203
rect 15669 11169 15703 11203
rect 17509 11169 17543 11203
rect 19993 11169 20027 11203
rect 21557 11169 21591 11203
rect 4199 11101 4233 11135
rect 4721 11101 4755 11135
rect 5273 11101 5307 11135
rect 5457 11101 5491 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 6653 11101 6687 11135
rect 6837 11101 6871 11135
rect 9503 11101 9537 11135
rect 10692 11101 10726 11135
rect 14749 11101 14783 11135
rect 14841 11101 14875 11135
rect 15761 11101 15795 11135
rect 16681 11101 16715 11135
rect 16773 11101 16807 11135
rect 16957 11101 16991 11135
rect 17049 11101 17083 11135
rect 17776 11101 17810 11135
rect 20177 11101 20211 11135
rect 20913 11101 20947 11135
rect 21097 11101 21131 11135
rect 21189 11101 21223 11135
rect 21281 11101 21315 11135
rect 22661 11101 22695 11135
rect 22809 11101 22843 11135
rect 23165 11101 23199 11135
rect 23857 11101 23891 11135
rect 24593 11101 24627 11135
rect 24777 11101 24811 11135
rect 24961 11101 24995 11135
rect 25973 11101 26007 11135
rect 26229 11101 26263 11135
rect 5917 11033 5951 11067
rect 7941 11033 7975 11067
rect 8217 11033 8251 11067
rect 15485 11033 15519 11067
rect 16497 11033 16531 11067
rect 21419 11033 21453 11067
rect 22937 11033 22971 11067
rect 23029 11033 23063 11067
rect 24869 11033 24903 11067
rect 4261 10965 4295 10999
rect 8125 10965 8159 10999
rect 9505 10965 9539 10999
rect 14933 10965 14967 10999
rect 23305 10965 23339 10999
rect 6009 10761 6043 10795
rect 9045 10761 9079 10795
rect 14749 10761 14783 10795
rect 16313 10761 16347 10795
rect 18245 10761 18279 10795
rect 19809 10761 19843 10795
rect 24685 10761 24719 10795
rect 26617 10761 26651 10795
rect 27721 10761 27755 10795
rect 2605 10693 2639 10727
rect 5089 10693 5123 10727
rect 8585 10693 8619 10727
rect 10057 10693 10091 10727
rect 13176 10693 13210 10727
rect 19441 10693 19475 10727
rect 19657 10693 19691 10727
rect 20821 10693 20855 10727
rect 22201 10693 22235 10727
rect 24317 10693 24351 10727
rect 24517 10693 24551 10727
rect 4813 10625 4847 10659
rect 5733 10625 5767 10659
rect 6561 10625 6595 10659
rect 6745 10625 6779 10659
rect 7113 10625 7147 10659
rect 8217 10625 8251 10659
rect 9229 10625 9263 10659
rect 10241 10625 10275 10659
rect 10425 10625 10459 10659
rect 12909 10625 12943 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 15945 10625 15979 10659
rect 16129 10625 16163 10659
rect 16865 10625 16899 10659
rect 17132 10625 17166 10659
rect 20637 10625 20671 10659
rect 20913 10625 20947 10659
rect 21005 10625 21039 10659
rect 22477 10625 22511 10659
rect 23305 10625 23339 10659
rect 23489 10625 23523 10659
rect 23581 10625 23615 10659
rect 23673 10625 23707 10659
rect 25237 10625 25271 10659
rect 25493 10625 25527 10659
rect 27169 10625 27203 10659
rect 27353 10625 27387 10659
rect 27445 10625 27479 10659
rect 27537 10625 27571 10659
rect 6009 10557 6043 10591
rect 8401 10557 8435 10591
rect 8493 10557 8527 10591
rect 9505 10557 9539 10591
rect 10517 10557 10551 10591
rect 15209 10557 15243 10591
rect 22385 10557 22419 10591
rect 7021 10489 7055 10523
rect 15117 10489 15151 10523
rect 3893 10421 3927 10455
rect 5825 10421 5859 10455
rect 9413 10421 9447 10455
rect 14289 10421 14323 10455
rect 15025 10421 15059 10455
rect 19625 10421 19659 10455
rect 21189 10421 21223 10455
rect 22201 10421 22235 10455
rect 22661 10421 22695 10455
rect 23857 10421 23891 10455
rect 24501 10421 24535 10455
rect 1777 10217 1811 10251
rect 2697 10217 2731 10251
rect 3985 10217 4019 10251
rect 5273 10217 5307 10251
rect 9229 10217 9263 10251
rect 9321 10217 9355 10251
rect 10609 10217 10643 10251
rect 16129 10217 16163 10251
rect 17969 10217 18003 10251
rect 18429 10217 18463 10251
rect 20729 10217 20763 10251
rect 21833 10217 21867 10251
rect 28365 10217 28399 10251
rect 3341 10149 3375 10183
rect 4353 10149 4387 10183
rect 12817 10149 12851 10183
rect 22293 10149 22327 10183
rect 23673 10149 23707 10183
rect 7665 10081 7699 10115
rect 9413 10081 9447 10115
rect 10149 10081 10183 10115
rect 10241 10081 10275 10115
rect 11437 10081 11471 10115
rect 14289 10081 14323 10115
rect 18153 10081 18187 10115
rect 21925 10081 21959 10115
rect 25145 10081 25179 10115
rect 1593 10013 1627 10047
rect 2605 10013 2639 10047
rect 2789 10013 2823 10047
rect 3249 10013 3283 10047
rect 3433 10013 3467 10047
rect 4169 10013 4203 10047
rect 4445 10013 4479 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 6377 10013 6411 10047
rect 6561 10013 6595 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 8309 10013 8343 10047
rect 9137 10013 9171 10047
rect 9861 10013 9895 10047
rect 10057 10013 10091 10047
rect 10425 10013 10459 10047
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 18245 10013 18279 10047
rect 19441 10013 19475 10047
rect 19534 10013 19568 10047
rect 19906 10013 19940 10047
rect 22109 10013 22143 10047
rect 23121 10013 23155 10047
rect 23305 10013 23339 10047
rect 23489 10013 23523 10047
rect 25412 10013 25446 10047
rect 26985 10013 27019 10047
rect 8401 9945 8435 9979
rect 11693 9945 11727 9979
rect 14534 9945 14568 9979
rect 17785 9945 17819 9979
rect 19717 9945 19751 9979
rect 19809 9945 19843 9979
rect 20545 9945 20579 9979
rect 20761 9945 20795 9979
rect 21833 9945 21867 9979
rect 23397 9945 23431 9979
rect 27230 9945 27264 9979
rect 6745 9877 6779 9911
rect 7297 9877 7331 9911
rect 15669 9877 15703 9911
rect 20085 9877 20119 9911
rect 20913 9877 20947 9911
rect 26525 9877 26559 9911
rect 7405 9673 7439 9707
rect 15209 9673 15243 9707
rect 22477 9673 22511 9707
rect 25789 9673 25823 9707
rect 3249 9605 3283 9639
rect 4905 9605 4939 9639
rect 7205 9605 7239 9639
rect 9588 9605 9622 9639
rect 12265 9605 12299 9639
rect 13084 9605 13118 9639
rect 19901 9605 19935 9639
rect 20111 9605 20145 9639
rect 1593 9537 1627 9571
rect 4261 9537 4295 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 5641 9537 5675 9571
rect 5769 9537 5803 9571
rect 6561 9537 6595 9571
rect 8309 9537 8343 9571
rect 9321 9537 9355 9571
rect 11897 9537 11931 9571
rect 12081 9537 12115 9571
rect 12817 9537 12851 9571
rect 15209 9537 15243 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 15853 9537 15887 9571
rect 19809 9537 19843 9571
rect 20018 9537 20052 9571
rect 20269 9537 20303 9571
rect 20913 9537 20947 9571
rect 22385 9537 22419 9571
rect 22753 9537 22787 9571
rect 23305 9537 23339 9571
rect 23572 9537 23606 9571
rect 25145 9537 25179 9571
rect 25238 9537 25272 9571
rect 25421 9537 25455 9571
rect 25513 9537 25547 9571
rect 25651 9537 25685 9571
rect 1869 9469 1903 9503
rect 4629 9469 4663 9503
rect 4721 9469 4755 9503
rect 8585 9469 8619 9503
rect 20729 9469 20763 9503
rect 22569 9469 22603 9503
rect 5365 9401 5399 9435
rect 7573 9401 7607 9435
rect 8493 9401 8527 9435
rect 22661 9401 22695 9435
rect 6653 9333 6687 9367
rect 7389 9333 7423 9367
rect 8125 9333 8159 9367
rect 10701 9333 10735 9367
rect 14197 9333 14231 9367
rect 19625 9333 19659 9367
rect 21097 9333 21131 9367
rect 24685 9333 24719 9367
rect 2973 9129 3007 9163
rect 4169 9129 4203 9163
rect 6377 9129 6411 9163
rect 7573 9129 7607 9163
rect 9597 9129 9631 9163
rect 16037 9129 16071 9163
rect 17325 9129 17359 9163
rect 19533 9129 19567 9163
rect 24041 9129 24075 9163
rect 26433 9129 26467 9163
rect 28273 9129 28307 9163
rect 13645 9061 13679 9095
rect 14933 9061 14967 9095
rect 16221 9061 16255 9095
rect 18889 9061 18923 9095
rect 1593 8993 1627 9027
rect 11805 8993 11839 9027
rect 15025 8993 15059 9027
rect 15945 8993 15979 9027
rect 19533 8993 19567 9027
rect 4353 8925 4387 8959
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 6929 8925 6963 8959
rect 7021 8925 7055 8959
rect 7573 8925 7607 8959
rect 7757 8925 7791 8959
rect 9413 8925 9447 8959
rect 11529 8925 11563 8959
rect 12633 8925 12667 8959
rect 12725 8925 12759 8959
rect 13461 8925 13495 8959
rect 14841 8925 14875 8959
rect 15117 8925 15151 8959
rect 15301 8925 15335 8959
rect 16037 8925 16071 8959
rect 16773 8925 16807 8959
rect 17141 8925 17175 8959
rect 18245 8925 18279 8959
rect 18338 8925 18372 8959
rect 18521 8925 18555 8959
rect 18613 8925 18647 8959
rect 18710 8925 18744 8959
rect 19717 8925 19751 8959
rect 20821 8925 20855 8959
rect 22661 8925 22695 8959
rect 25053 8925 25087 8959
rect 26893 8925 26927 8959
rect 1860 8857 1894 8891
rect 5273 8857 5307 8891
rect 6653 8857 6687 8891
rect 12357 8857 12391 8891
rect 15761 8857 15795 8891
rect 16957 8857 16991 8891
rect 17049 8857 17083 8891
rect 19441 8857 19475 8891
rect 21088 8857 21122 8891
rect 22928 8857 22962 8891
rect 25320 8857 25354 8891
rect 27138 8857 27172 8891
rect 4537 8789 4571 8823
rect 5457 8789 5491 8823
rect 12541 8789 12575 8823
rect 12909 8789 12943 8823
rect 14565 8789 14599 8823
rect 19901 8789 19935 8823
rect 22201 8789 22235 8823
rect 5273 8585 5307 8619
rect 7941 8585 7975 8619
rect 13093 8585 13127 8619
rect 15853 8585 15887 8619
rect 17877 8585 17911 8619
rect 26157 8585 26191 8619
rect 6561 8517 6595 8551
rect 11958 8517 11992 8551
rect 15393 8517 15427 8551
rect 19533 8517 19567 8551
rect 20729 8517 20763 8551
rect 22998 8517 23032 8551
rect 5457 8449 5491 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7021 8449 7055 8483
rect 7113 8449 7147 8483
rect 7665 8449 7699 8483
rect 11713 8449 11747 8483
rect 13553 8449 13587 8483
rect 15669 8449 15703 8483
rect 18061 8449 18095 8483
rect 18153 8449 18187 8483
rect 18322 8449 18356 8483
rect 18439 8439 18473 8473
rect 19349 8449 19383 8483
rect 19625 8449 19659 8483
rect 19717 8449 19751 8483
rect 20453 8449 20487 8483
rect 20545 8449 20579 8483
rect 22017 8449 22051 8483
rect 22753 8449 22787 8483
rect 25044 8449 25078 8483
rect 7941 8381 7975 8415
rect 15577 8381 15611 8415
rect 24777 8381 24811 8415
rect 5549 8313 5583 8347
rect 5641 8313 5675 8347
rect 7757 8313 7791 8347
rect 24133 8313 24167 8347
rect 13737 8245 13771 8279
rect 15669 8245 15703 8279
rect 19901 8245 19935 8279
rect 22201 8245 22235 8279
rect 4537 8041 4571 8075
rect 4721 8041 4755 8075
rect 18245 8041 18279 8075
rect 21189 8041 21223 8075
rect 22293 8041 22327 8075
rect 23397 8041 23431 8075
rect 28365 8041 28399 8075
rect 13277 7973 13311 8007
rect 7113 7905 7147 7939
rect 18429 7905 18463 7939
rect 1777 7837 1811 7871
rect 4261 7837 4295 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 7205 7837 7239 7871
rect 9229 7837 9263 7871
rect 9496 7837 9530 7871
rect 12633 7837 12667 7871
rect 12781 7837 12815 7871
rect 13001 7837 13035 7871
rect 13098 7837 13132 7871
rect 14289 7837 14323 7871
rect 14545 7837 14579 7871
rect 16129 7837 16163 7871
rect 16222 7837 16256 7871
rect 16405 7837 16439 7871
rect 16497 7837 16531 7871
rect 16635 7837 16669 7871
rect 18337 7837 18371 7871
rect 18705 7837 18739 7871
rect 19809 7837 19843 7871
rect 21649 7837 21683 7871
rect 21797 7837 21831 7871
rect 22114 7837 22148 7871
rect 22753 7837 22787 7871
rect 22901 7837 22935 7871
rect 23218 7837 23252 7871
rect 25053 7837 25087 7871
rect 25320 7837 25354 7871
rect 26985 7837 27019 7871
rect 12909 7769 12943 7803
rect 20076 7769 20110 7803
rect 21925 7769 21959 7803
rect 22017 7769 22051 7803
rect 23029 7769 23063 7803
rect 23121 7769 23155 7803
rect 27230 7769 27264 7803
rect 1593 7701 1627 7735
rect 6377 7701 6411 7735
rect 10609 7701 10643 7735
rect 15669 7701 15703 7735
rect 16773 7701 16807 7735
rect 17969 7701 18003 7735
rect 18613 7701 18647 7735
rect 26433 7701 26467 7735
rect 5825 7497 5859 7531
rect 12725 7497 12759 7531
rect 16129 7497 16163 7531
rect 17509 7497 17543 7531
rect 20729 7497 20763 7531
rect 23949 7497 23983 7531
rect 26617 7497 26651 7531
rect 8576 7429 8610 7463
rect 10149 7429 10183 7463
rect 12357 7429 12391 7463
rect 13185 7429 13219 7463
rect 13385 7429 13419 7463
rect 14013 7429 14047 7463
rect 17141 7429 17175 7463
rect 17233 7429 17267 7463
rect 20361 7429 20395 7463
rect 20453 7429 20487 7463
rect 1777 7361 1811 7395
rect 2881 7361 2915 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 10333 7361 10367 7395
rect 10425 7361 10459 7395
rect 10701 7361 10735 7395
rect 12081 7361 12115 7395
rect 12229 7361 12263 7395
rect 12449 7361 12483 7395
rect 12587 7361 12621 7395
rect 14289 7361 14323 7395
rect 15485 7361 15519 7395
rect 15761 7361 15795 7395
rect 15945 7361 15979 7395
rect 16865 7361 16899 7395
rect 17013 7361 17047 7395
rect 17330 7361 17364 7395
rect 18797 7361 18831 7395
rect 20177 7361 20211 7395
rect 20545 7361 20579 7395
rect 22825 7361 22859 7395
rect 25504 7361 25538 7395
rect 8309 7293 8343 7327
rect 14197 7293 14231 7327
rect 18613 7293 18647 7327
rect 22569 7293 22603 7327
rect 25237 7293 25271 7327
rect 9689 7225 9723 7259
rect 13553 7225 13587 7259
rect 1593 7157 1627 7191
rect 2973 7157 3007 7191
rect 5457 7157 5491 7191
rect 10609 7157 10643 7191
rect 13369 7157 13403 7191
rect 14289 7157 14323 7191
rect 14473 7157 14507 7191
rect 15945 7157 15979 7191
rect 18981 7157 19015 7191
rect 9321 6953 9355 6987
rect 13553 6953 13587 6987
rect 14473 6953 14507 6987
rect 16681 6953 16715 6987
rect 20821 6953 20855 6987
rect 24041 6953 24075 6987
rect 26249 6953 26283 6987
rect 28089 6953 28123 6987
rect 1593 6817 1627 6851
rect 6469 6817 6503 6851
rect 17325 6817 17359 6851
rect 19441 6817 19475 6851
rect 26709 6817 26743 6851
rect 1860 6749 1894 6783
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 9137 6749 9171 6783
rect 10057 6749 10091 6783
rect 11529 6749 11563 6783
rect 11677 6749 11711 6783
rect 11805 6749 11839 6783
rect 12035 6749 12069 6783
rect 14657 6749 14691 6783
rect 14749 6749 14783 6783
rect 14933 6749 14967 6783
rect 15025 6749 15059 6783
rect 15853 6749 15887 6783
rect 15945 6749 15979 6783
rect 16865 6749 16899 6783
rect 16957 6749 16991 6783
rect 17049 6749 17083 6783
rect 19625 6749 19659 6783
rect 20269 6749 20303 6783
rect 20661 6749 20695 6783
rect 21281 6749 21315 6783
rect 21557 6749 21591 6783
rect 21649 6749 21683 6783
rect 22293 6749 22327 6783
rect 22477 6749 22511 6783
rect 23489 6749 23523 6783
rect 23857 6749 23891 6783
rect 24869 6749 24903 6783
rect 25136 6749 25170 6783
rect 5641 6681 5675 6715
rect 6736 6681 6770 6715
rect 11897 6681 11931 6715
rect 13369 6681 13403 6715
rect 17167 6681 17201 6715
rect 20453 6681 20487 6715
rect 20545 6681 20579 6715
rect 21465 6681 21499 6715
rect 22661 6681 22695 6715
rect 23673 6681 23707 6715
rect 23765 6681 23799 6715
rect 26954 6681 26988 6715
rect 2973 6613 3007 6647
rect 5549 6613 5583 6647
rect 7849 6613 7883 6647
rect 9873 6613 9907 6647
rect 12173 6613 12207 6647
rect 13574 6613 13608 6647
rect 13737 6613 13771 6647
rect 16129 6613 16163 6647
rect 19809 6613 19843 6647
rect 21833 6613 21867 6647
rect 2973 6409 3007 6443
rect 5549 6409 5583 6443
rect 6653 6409 6687 6443
rect 15301 6409 15335 6443
rect 15761 6409 15795 6443
rect 20545 6409 20579 6443
rect 22385 6409 22419 6443
rect 24685 6409 24719 6443
rect 26525 6409 26559 6443
rect 1860 6341 1894 6375
rect 7564 6341 7598 6375
rect 9956 6341 9990 6375
rect 13829 6341 13863 6375
rect 13921 6341 13955 6375
rect 22043 6341 22077 6375
rect 22217 6341 22251 6375
rect 25390 6341 25424 6375
rect 1593 6273 1627 6307
rect 3525 6273 3559 6307
rect 4353 6273 4387 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 9689 6273 9723 6307
rect 11713 6273 11747 6307
rect 11980 6273 12014 6307
rect 13553 6273 13587 6307
rect 13646 6273 13680 6307
rect 14059 6273 14093 6307
rect 14749 6273 14783 6307
rect 14933 6273 14967 6307
rect 15025 6273 15059 6307
rect 15117 6273 15151 6307
rect 15945 6273 15979 6307
rect 16037 6273 16071 6307
rect 16221 6273 16255 6307
rect 16313 6273 16347 6307
rect 17592 6273 17626 6307
rect 19165 6273 19199 6307
rect 19432 6273 19466 6307
rect 23561 6273 23595 6307
rect 5917 6205 5951 6239
rect 7297 6205 7331 6239
rect 17325 6205 17359 6239
rect 23305 6205 23339 6239
rect 25145 6205 25179 6239
rect 4537 6137 4571 6171
rect 3709 6069 3743 6103
rect 8677 6069 8711 6103
rect 11069 6069 11103 6103
rect 13093 6069 13127 6103
rect 14197 6069 14231 6103
rect 18705 6069 18739 6103
rect 22201 6069 22235 6103
rect 2973 5865 3007 5899
rect 3341 5865 3375 5899
rect 4353 5865 4387 5899
rect 5181 5865 5215 5899
rect 8033 5865 8067 5899
rect 10517 5865 10551 5899
rect 11805 5865 11839 5899
rect 15485 5865 15519 5899
rect 18705 5865 18739 5899
rect 18889 5865 18923 5899
rect 21557 5865 21591 5899
rect 22569 5865 22603 5899
rect 25973 5865 26007 5899
rect 12817 5797 12851 5831
rect 17969 5797 18003 5831
rect 1593 5729 1627 5763
rect 3985 5729 4019 5763
rect 6653 5729 6687 5763
rect 9137 5729 9171 5763
rect 12449 5729 12483 5763
rect 20177 5729 20211 5763
rect 24593 5729 24627 5763
rect 1860 5661 1894 5695
rect 4169 5661 4203 5695
rect 4997 5661 5031 5695
rect 9393 5661 9427 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 12633 5661 12667 5695
rect 13369 5661 13403 5695
rect 13461 5661 13495 5695
rect 14841 5661 14875 5695
rect 14989 5661 15023 5695
rect 15117 5661 15151 5695
rect 15306 5661 15340 5695
rect 17417 5661 17451 5695
rect 17785 5661 17819 5695
rect 22017 5661 22051 5695
rect 22385 5661 22419 5695
rect 26985 5661 27019 5695
rect 4813 5593 4847 5627
rect 6920 5593 6954 5627
rect 11437 5593 11471 5627
rect 15209 5593 15243 5627
rect 16589 5593 16623 5627
rect 17601 5593 17635 5627
rect 17693 5593 17727 5627
rect 18521 5593 18555 5627
rect 20444 5593 20478 5627
rect 22201 5593 22235 5627
rect 22293 5593 22327 5627
rect 24860 5593 24894 5627
rect 27230 5593 27264 5627
rect 13645 5525 13679 5559
rect 16681 5525 16715 5559
rect 18731 5525 18765 5559
rect 28365 5525 28399 5559
rect 6009 5321 6043 5355
rect 9321 5321 9355 5355
rect 11161 5321 11195 5355
rect 12541 5321 12575 5355
rect 15577 5321 15611 5355
rect 19533 5321 19567 5355
rect 26617 5321 26651 5355
rect 2964 5253 2998 5287
rect 12173 5253 12207 5287
rect 13544 5253 13578 5287
rect 17233 5253 17267 5287
rect 18420 5253 18454 5287
rect 19993 5253 20027 5287
rect 20209 5253 20243 5287
rect 25482 5253 25516 5287
rect 1961 5185 1995 5219
rect 2697 5185 2731 5219
rect 4629 5185 4663 5219
rect 4896 5185 4930 5219
rect 7941 5185 7975 5219
rect 8208 5185 8242 5219
rect 9781 5185 9815 5219
rect 10048 5185 10082 5219
rect 11989 5185 12023 5219
rect 12265 5185 12299 5219
rect 12357 5185 12391 5219
rect 13277 5185 13311 5219
rect 15117 5185 15151 5219
rect 15393 5185 15427 5219
rect 16129 5185 16163 5219
rect 17049 5185 17083 5219
rect 25237 5185 25271 5219
rect 27445 5185 27479 5219
rect 15301 5117 15335 5151
rect 16865 5117 16899 5151
rect 18153 5117 18187 5151
rect 27169 5117 27203 5151
rect 2145 4981 2179 5015
rect 4077 4981 4111 5015
rect 14657 4981 14691 5015
rect 15393 4981 15427 5015
rect 16221 4981 16255 5015
rect 20177 4981 20211 5015
rect 20361 4981 20395 5015
rect 3157 4777 3191 4811
rect 5917 4777 5951 4811
rect 10793 4777 10827 4811
rect 13737 4777 13771 4811
rect 14841 4777 14875 4811
rect 18245 4777 18279 4811
rect 21925 4777 21959 4811
rect 24041 4777 24075 4811
rect 25973 4777 26007 4811
rect 27813 4777 27847 4811
rect 15025 4709 15059 4743
rect 18429 4709 18463 4743
rect 20085 4709 20119 4743
rect 1777 4641 1811 4675
rect 4537 4641 4571 4675
rect 12357 4641 12391 4675
rect 26433 4641 26467 4675
rect 2033 4573 2067 4607
rect 7205 4573 7239 4607
rect 7472 4573 7506 4607
rect 9413 4573 9447 4607
rect 15577 4573 15611 4607
rect 15844 4573 15878 4607
rect 19441 4573 19475 4607
rect 19589 4573 19623 4607
rect 19906 4573 19940 4607
rect 20545 4573 20579 4607
rect 20812 4573 20846 4607
rect 22661 4573 22695 4607
rect 22928 4573 22962 4607
rect 24593 4573 24627 4607
rect 24849 4573 24883 4607
rect 26689 4573 26723 4607
rect 4782 4505 4816 4539
rect 9680 4505 9714 4539
rect 12624 4505 12658 4539
rect 14657 4505 14691 4539
rect 14857 4505 14891 4539
rect 18061 4505 18095 4539
rect 18261 4505 18295 4539
rect 19717 4505 19751 4539
rect 19809 4505 19843 4539
rect 8585 4437 8619 4471
rect 16957 4437 16991 4471
rect 5181 4233 5215 4267
rect 8125 4233 8159 4267
rect 15945 4233 15979 4267
rect 10517 4165 10551 4199
rect 13737 4165 13771 4199
rect 13937 4165 13971 4199
rect 14810 4165 14844 4199
rect 17110 4165 17144 4199
rect 22109 4165 22143 4199
rect 22293 4165 22327 4199
rect 1685 4097 1719 4131
rect 1952 4097 1986 4131
rect 3801 4097 3835 4131
rect 4068 4097 4102 4131
rect 7012 4097 7046 4131
rect 8852 4097 8886 4131
rect 10701 4097 10735 4131
rect 11897 4097 11931 4131
rect 12164 4097 12198 4131
rect 19165 4097 19199 4131
rect 19432 4097 19466 4131
rect 25504 4097 25538 4131
rect 6745 4029 6779 4063
rect 8585 4029 8619 4063
rect 14565 4029 14599 4063
rect 16865 4029 16899 4063
rect 25237 4029 25271 4063
rect 3065 3961 3099 3995
rect 9965 3961 9999 3995
rect 26617 3961 26651 3995
rect 13277 3893 13311 3927
rect 13921 3893 13955 3927
rect 14105 3893 14139 3927
rect 18245 3893 18279 3927
rect 20545 3893 20579 3927
rect 4169 3689 4203 3723
rect 6837 3689 6871 3723
rect 13277 3689 13311 3723
rect 23765 3689 23799 3723
rect 28365 3689 28399 3723
rect 3341 3621 3375 3655
rect 1961 3553 1995 3587
rect 5457 3553 5491 3587
rect 10885 3553 10919 3587
rect 20545 3553 20579 3587
rect 22385 3553 22419 3587
rect 26985 3553 27019 3587
rect 4077 3485 4111 3519
rect 5724 3485 5758 3519
rect 11152 3485 11186 3519
rect 12725 3485 12759 3519
rect 13001 3485 13035 3519
rect 13093 3485 13127 3519
rect 14749 3485 14783 3519
rect 17417 3485 17451 3519
rect 20812 3485 20846 3519
rect 22641 3485 22675 3519
rect 25145 3485 25179 3519
rect 27241 3485 27275 3519
rect 2206 3417 2240 3451
rect 12909 3417 12943 3451
rect 15016 3417 15050 3451
rect 17684 3417 17718 3451
rect 25412 3417 25446 3451
rect 12265 3349 12299 3383
rect 16129 3349 16163 3383
rect 18797 3349 18831 3383
rect 21925 3349 21959 3383
rect 26525 3349 26559 3383
rect 3617 3145 3651 3179
rect 11161 3145 11195 3179
rect 13829 3145 13863 3179
rect 18245 3145 18279 3179
rect 20913 3145 20947 3179
rect 23489 3145 23523 3179
rect 10048 3077 10082 3111
rect 12716 3077 12750 3111
rect 17132 3077 17166 3111
rect 19778 3077 19812 3111
rect 24216 3077 24250 3111
rect 2237 3009 2271 3043
rect 2513 3009 2547 3043
rect 4353 3009 4387 3043
rect 4620 3009 4654 3043
rect 9781 3009 9815 3043
rect 12449 3009 12483 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 15025 3009 15059 3043
rect 15761 3009 15795 3043
rect 15945 3009 15979 3043
rect 16865 3009 16899 3043
rect 22109 3009 22143 3043
rect 22376 3009 22410 3043
rect 23949 3009 23983 3043
rect 19533 2941 19567 2975
rect 15209 2873 15243 2907
rect 5733 2805 5767 2839
rect 25329 2805 25363 2839
rect 1685 2601 1719 2635
rect 3341 2601 3375 2635
rect 5365 2601 5399 2635
rect 7297 2601 7331 2635
rect 11253 2601 11287 2635
rect 13645 2601 13679 2635
rect 17969 2601 18003 2635
rect 18429 2601 18463 2635
rect 18889 2601 18923 2635
rect 28365 2601 28399 2635
rect 12541 2533 12575 2567
rect 16221 2533 16255 2567
rect 1961 2465 1995 2499
rect 9873 2465 9907 2499
rect 14841 2465 14875 2499
rect 18521 2465 18555 2499
rect 24593 2465 24627 2499
rect 26985 2465 27019 2499
rect 3985 2397 4019 2431
rect 5917 2397 5951 2431
rect 6184 2397 6218 2431
rect 10140 2397 10174 2431
rect 11989 2397 12023 2431
rect 12173 2397 12207 2431
rect 12357 2397 12391 2431
rect 13001 2397 13035 2431
rect 13094 2397 13128 2431
rect 13277 2397 13311 2431
rect 13369 2397 13403 2431
rect 13507 2397 13541 2431
rect 17325 2397 17359 2431
rect 17473 2397 17507 2431
rect 17601 2397 17635 2431
rect 17693 2397 17727 2431
rect 17790 2397 17824 2431
rect 18705 2397 18739 2431
rect 21281 2397 21315 2431
rect 27241 2397 27275 2431
rect 2206 2329 2240 2363
rect 4252 2329 4286 2363
rect 5825 2329 5859 2363
rect 12265 2329 12299 2363
rect 15108 2329 15142 2363
rect 18429 2329 18463 2363
rect 21548 2329 21582 2363
rect 24860 2329 24894 2363
rect 22661 2261 22695 2295
rect 25973 2261 26007 2295
rect 2329 2057 2363 2091
rect 5549 2057 5583 2091
rect 9321 2057 9355 2091
rect 13921 2057 13955 2091
rect 18337 2057 18371 2091
rect 20177 2057 20211 2091
rect 21281 2057 21315 2091
rect 23397 2057 23431 2091
rect 25237 2057 25271 2091
rect 8208 1989 8242 2023
rect 11713 1989 11747 2023
rect 11929 1989 11963 2023
rect 12808 1989 12842 2023
rect 15200 1989 15234 2023
rect 17224 1989 17258 2023
rect 24102 1989 24136 2023
rect 25973 1989 26007 2023
rect 3709 1921 3743 1955
rect 4169 1921 4203 1955
rect 4436 1921 4470 1955
rect 9781 1921 9815 1955
rect 10048 1921 10082 1955
rect 12541 1921 12575 1955
rect 19053 1921 19087 1955
rect 20637 1921 20671 1955
rect 20730 1921 20764 1955
rect 20913 1921 20947 1955
rect 21005 1921 21039 1955
rect 21102 1921 21136 1955
rect 22017 1921 22051 1955
rect 22284 1921 22318 1955
rect 23857 1921 23891 1955
rect 25697 1921 25731 1955
rect 25881 1921 25915 1955
rect 26065 1921 26099 1955
rect 1777 1853 1811 1887
rect 3433 1853 3467 1887
rect 7941 1853 7975 1887
rect 14933 1853 14967 1887
rect 16957 1853 16991 1887
rect 18797 1853 18831 1887
rect 11161 1785 11195 1819
rect 16313 1785 16347 1819
rect 11897 1717 11931 1751
rect 12081 1717 12115 1751
rect 26249 1717 26283 1751
rect 14565 1513 14599 1547
rect 14749 1513 14783 1547
rect 14657 1445 14691 1479
rect 1961 1377 1995 1411
rect 13001 1377 13035 1411
rect 3985 1309 4019 1343
rect 9137 1309 9171 1343
rect 9404 1309 9438 1343
rect 11989 1309 12023 1343
rect 12173 1309 12207 1343
rect 14381 1309 14415 1343
rect 14841 1309 14875 1343
rect 15761 1309 15795 1343
rect 16037 1309 16071 1343
rect 16129 1309 16163 1343
rect 17509 1309 17543 1343
rect 19901 1309 19935 1343
rect 20269 1309 20303 1343
rect 20913 1309 20947 1343
rect 21097 1309 21131 1343
rect 21281 1309 21315 1343
rect 22385 1309 22419 1343
rect 22652 1309 22686 1343
rect 25237 1309 25271 1343
rect 1685 1241 1719 1275
rect 2228 1241 2262 1275
rect 4252 1241 4286 1275
rect 15945 1241 15979 1275
rect 17776 1241 17810 1275
rect 20085 1241 20119 1275
rect 20177 1241 20211 1275
rect 21189 1241 21223 1275
rect 25482 1241 25516 1275
rect 3341 1173 3375 1207
rect 5365 1173 5399 1207
rect 5733 1173 5767 1207
rect 10517 1173 10551 1207
rect 14933 1173 14967 1207
rect 16313 1173 16347 1207
rect 18889 1173 18923 1207
rect 20453 1173 20487 1207
rect 21465 1173 21499 1207
rect 23765 1173 23799 1207
rect 26617 1173 26651 1207
<< metal1 >>
rect 1104 32666 29048 32688
rect 1104 32614 7896 32666
rect 7948 32614 7960 32666
rect 8012 32614 8024 32666
rect 8076 32614 8088 32666
rect 8140 32614 8152 32666
rect 8204 32614 14842 32666
rect 14894 32614 14906 32666
rect 14958 32614 14970 32666
rect 15022 32614 15034 32666
rect 15086 32614 15098 32666
rect 15150 32614 21788 32666
rect 21840 32614 21852 32666
rect 21904 32614 21916 32666
rect 21968 32614 21980 32666
rect 22032 32614 22044 32666
rect 22096 32614 28734 32666
rect 28786 32614 28798 32666
rect 28850 32614 28862 32666
rect 28914 32614 28926 32666
rect 28978 32614 28990 32666
rect 29042 32614 29048 32666
rect 1104 32592 29048 32614
rect 4338 32512 4344 32564
rect 4396 32512 4402 32564
rect 5166 32512 5172 32564
rect 5224 32512 5230 32564
rect 8570 32512 8576 32564
rect 8628 32512 8634 32564
rect 9490 32512 9496 32564
rect 9548 32552 9554 32564
rect 11057 32555 11115 32561
rect 11057 32552 11069 32555
rect 9548 32524 11069 32552
rect 9548 32512 9554 32524
rect 11057 32521 11069 32524
rect 11103 32552 11115 32555
rect 11238 32552 11244 32564
rect 11103 32524 11244 32552
rect 11103 32521 11115 32524
rect 11057 32515 11115 32521
rect 11238 32512 11244 32524
rect 11296 32512 11302 32564
rect 3329 32487 3387 32493
rect 3329 32453 3341 32487
rect 3375 32484 3387 32487
rect 8478 32484 8484 32496
rect 3375 32456 8484 32484
rect 3375 32453 3387 32456
rect 3329 32447 3387 32453
rect 8478 32444 8484 32456
rect 8536 32444 8542 32496
rect 12360 32456 15608 32484
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 1670 32416 1676 32428
rect 1627 32388 1676 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 3973 32419 4031 32425
rect 3973 32385 3985 32419
rect 4019 32416 4031 32419
rect 5166 32416 5172 32428
rect 4019 32388 5172 32416
rect 4019 32385 4031 32388
rect 3973 32379 4031 32385
rect 5166 32376 5172 32388
rect 5224 32376 5230 32428
rect 8294 32376 8300 32428
rect 8352 32416 8358 32428
rect 12360 32425 12388 32456
rect 14292 32428 14320 32456
rect 12345 32419 12403 32425
rect 12345 32416 12357 32419
rect 8352 32388 12357 32416
rect 8352 32376 8358 32388
rect 12345 32385 12357 32388
rect 12391 32385 12403 32419
rect 12345 32379 12403 32385
rect 12526 32376 12532 32428
rect 12584 32376 12590 32428
rect 14274 32376 14280 32428
rect 14332 32376 14338 32428
rect 14458 32376 14464 32428
rect 14516 32376 14522 32428
rect 14936 32425 14964 32456
rect 15580 32425 15608 32456
rect 14921 32419 14979 32425
rect 14921 32385 14933 32419
rect 14967 32385 14979 32419
rect 14921 32379 14979 32385
rect 15105 32419 15163 32425
rect 15105 32385 15117 32419
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 15565 32419 15623 32425
rect 15565 32385 15577 32419
rect 15611 32385 15623 32419
rect 15565 32379 15623 32385
rect 4798 32308 4804 32360
rect 4856 32308 4862 32360
rect 8202 32308 8208 32360
rect 8260 32348 8266 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 8260 32320 9137 32348
rect 8260 32308 8266 32320
rect 9125 32317 9137 32320
rect 9171 32317 9183 32351
rect 9125 32311 9183 32317
rect 9490 32308 9496 32360
rect 9548 32308 9554 32360
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32348 10747 32351
rect 11146 32348 11152 32360
rect 10735 32320 11152 32348
rect 10735 32317 10747 32320
rect 10689 32311 10747 32317
rect 11146 32308 11152 32320
rect 11204 32308 11210 32360
rect 3326 32240 3332 32292
rect 3384 32280 3390 32292
rect 4341 32283 4399 32289
rect 4341 32280 4353 32283
rect 3384 32252 4353 32280
rect 3384 32240 3390 32252
rect 4341 32249 4353 32252
rect 4387 32249 4399 32283
rect 4341 32243 4399 32249
rect 5166 32240 5172 32292
rect 5224 32240 5230 32292
rect 5997 32283 6055 32289
rect 5997 32249 6009 32283
rect 6043 32280 6055 32283
rect 8386 32280 8392 32292
rect 6043 32252 8392 32280
rect 6043 32249 6055 32252
rect 5997 32243 6055 32249
rect 8386 32240 8392 32252
rect 8444 32240 8450 32292
rect 8570 32240 8576 32292
rect 8628 32280 8634 32292
rect 9508 32280 9536 32308
rect 11057 32283 11115 32289
rect 8628 32252 9536 32280
rect 10060 32252 11008 32280
rect 8628 32240 8634 32252
rect 4890 32172 4896 32224
rect 4948 32212 4954 32224
rect 6733 32215 6791 32221
rect 6733 32212 6745 32215
rect 4948 32184 6745 32212
rect 4948 32172 4954 32184
rect 6733 32181 6745 32184
rect 6779 32181 6791 32215
rect 6733 32175 6791 32181
rect 7377 32215 7435 32221
rect 7377 32181 7389 32215
rect 7423 32212 7435 32215
rect 10060 32212 10088 32252
rect 7423 32184 10088 32212
rect 7423 32181 7435 32184
rect 7377 32175 7435 32181
rect 10134 32172 10140 32224
rect 10192 32172 10198 32224
rect 10980 32212 11008 32252
rect 11057 32249 11069 32283
rect 11103 32280 11115 32283
rect 11238 32280 11244 32292
rect 11103 32252 11244 32280
rect 11103 32249 11115 32252
rect 11057 32243 11115 32249
rect 11238 32240 11244 32252
rect 11296 32240 11302 32292
rect 11885 32283 11943 32289
rect 11885 32249 11897 32283
rect 11931 32280 11943 32283
rect 15120 32280 15148 32379
rect 15746 32376 15752 32428
rect 15804 32376 15810 32428
rect 11931 32252 15148 32280
rect 11931 32249 11943 32252
rect 11885 32243 11943 32249
rect 13078 32212 13084 32224
rect 10980 32184 13084 32212
rect 13078 32172 13084 32184
rect 13136 32172 13142 32224
rect 13173 32215 13231 32221
rect 13173 32181 13185 32215
rect 13219 32212 13231 32215
rect 15102 32212 15108 32224
rect 13219 32184 15108 32212
rect 13219 32181 13231 32184
rect 13173 32175 13231 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 1104 32122 28888 32144
rect 1104 32070 4423 32122
rect 4475 32070 4487 32122
rect 4539 32070 4551 32122
rect 4603 32070 4615 32122
rect 4667 32070 4679 32122
rect 4731 32070 11369 32122
rect 11421 32070 11433 32122
rect 11485 32070 11497 32122
rect 11549 32070 11561 32122
rect 11613 32070 11625 32122
rect 11677 32070 18315 32122
rect 18367 32070 18379 32122
rect 18431 32070 18443 32122
rect 18495 32070 18507 32122
rect 18559 32070 18571 32122
rect 18623 32070 25261 32122
rect 25313 32070 25325 32122
rect 25377 32070 25389 32122
rect 25441 32070 25453 32122
rect 25505 32070 25517 32122
rect 25569 32070 28888 32122
rect 1104 32048 28888 32070
rect 2774 31968 2780 32020
rect 2832 32008 2838 32020
rect 4525 32011 4583 32017
rect 4525 32008 4537 32011
rect 2832 31980 4537 32008
rect 2832 31968 2838 31980
rect 4525 31977 4537 31980
rect 4571 31977 4583 32011
rect 5258 32008 5264 32020
rect 4525 31971 4583 31977
rect 4632 31980 5264 32008
rect 4632 31940 4660 31980
rect 5258 31968 5264 31980
rect 5316 31968 5322 32020
rect 6733 32011 6791 32017
rect 6733 31977 6745 32011
rect 6779 32008 6791 32011
rect 7377 32011 7435 32017
rect 6779 31980 6914 32008
rect 6779 31977 6791 31980
rect 6733 31971 6791 31977
rect 4172 31912 4660 31940
rect 3326 31832 3332 31884
rect 3384 31832 3390 31884
rect 1578 31764 1584 31816
rect 1636 31764 1642 31816
rect 3973 31807 4031 31813
rect 3973 31773 3985 31807
rect 4019 31804 4031 31807
rect 4172 31804 4200 31912
rect 5166 31900 5172 31952
rect 5224 31940 5230 31952
rect 5905 31943 5963 31949
rect 5905 31940 5917 31943
rect 5224 31912 5917 31940
rect 5224 31900 5230 31912
rect 5905 31909 5917 31912
rect 5951 31909 5963 31943
rect 6886 31940 6914 31980
rect 7377 31977 7389 32011
rect 7423 32008 7435 32011
rect 12526 32008 12532 32020
rect 7423 31980 12532 32008
rect 7423 31977 7435 31980
rect 7377 31971 7435 31977
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 9309 31943 9367 31949
rect 6886 31912 9168 31940
rect 5905 31903 5963 31909
rect 9030 31872 9036 31884
rect 4264 31844 9036 31872
rect 4264 31813 4292 31844
rect 9030 31832 9036 31844
rect 9088 31832 9094 31884
rect 9140 31872 9168 31912
rect 9309 31909 9321 31943
rect 9355 31940 9367 31943
rect 11882 31940 11888 31952
rect 9355 31912 11888 31940
rect 9355 31909 9367 31912
rect 9309 31903 9367 31909
rect 11882 31900 11888 31912
rect 11940 31900 11946 31952
rect 13265 31943 13323 31949
rect 13265 31909 13277 31943
rect 13311 31940 13323 31943
rect 13311 31912 15792 31940
rect 13311 31909 13323 31912
rect 13265 31903 13323 31909
rect 9490 31872 9496 31884
rect 9140 31844 9496 31872
rect 9490 31832 9496 31844
rect 9548 31832 9554 31884
rect 9861 31875 9919 31881
rect 9861 31841 9873 31875
rect 9907 31872 9919 31875
rect 10962 31872 10968 31884
rect 9907 31844 10968 31872
rect 9907 31841 9919 31844
rect 9861 31835 9919 31841
rect 10962 31832 10968 31844
rect 11020 31832 11026 31884
rect 11057 31875 11115 31881
rect 11057 31841 11069 31875
rect 11103 31872 11115 31875
rect 11103 31844 11652 31872
rect 11103 31841 11115 31844
rect 11057 31835 11115 31841
rect 4430 31813 4436 31816
rect 4019 31776 4200 31804
rect 4249 31807 4307 31813
rect 4019 31773 4031 31776
rect 3973 31767 4031 31773
rect 4249 31773 4261 31807
rect 4295 31773 4307 31807
rect 4249 31767 4307 31773
rect 4393 31807 4436 31813
rect 4393 31773 4405 31807
rect 4393 31767 4436 31773
rect 4430 31764 4436 31767
rect 4488 31764 4494 31816
rect 4798 31764 4804 31816
rect 4856 31804 4862 31816
rect 5537 31807 5595 31813
rect 5537 31804 5549 31807
rect 4856 31776 5549 31804
rect 4856 31764 4862 31776
rect 5537 31773 5549 31776
rect 5583 31773 5595 31807
rect 5537 31767 5595 31773
rect 7558 31764 7564 31816
rect 7616 31804 7622 31816
rect 8202 31804 8208 31816
rect 7616 31776 8208 31804
rect 7616 31764 7622 31776
rect 8202 31764 8208 31776
rect 8260 31764 8266 31816
rect 8570 31764 8576 31816
rect 8628 31764 8634 31816
rect 10229 31807 10287 31813
rect 10229 31773 10241 31807
rect 10275 31773 10287 31807
rect 10229 31767 10287 31773
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31804 10747 31807
rect 11146 31804 11152 31816
rect 10735 31776 11152 31804
rect 10735 31773 10747 31776
rect 10689 31767 10747 31773
rect 4157 31739 4215 31745
rect 4157 31705 4169 31739
rect 4203 31736 4215 31739
rect 4706 31736 4712 31748
rect 4203 31708 4712 31736
rect 4203 31705 4215 31708
rect 4157 31699 4215 31705
rect 4706 31696 4712 31708
rect 4764 31696 4770 31748
rect 5902 31628 5908 31680
rect 5960 31628 5966 31680
rect 8588 31677 8616 31764
rect 10244 31680 10272 31767
rect 11146 31764 11152 31776
rect 11204 31804 11210 31816
rect 11514 31804 11520 31816
rect 11204 31776 11520 31804
rect 11204 31764 11210 31776
rect 11514 31764 11520 31776
rect 11572 31764 11578 31816
rect 11624 31804 11652 31844
rect 11698 31832 11704 31884
rect 11756 31872 11762 31884
rect 11756 31844 15608 31872
rect 11756 31832 11762 31844
rect 11885 31807 11943 31813
rect 11885 31804 11897 31807
rect 11624 31776 11897 31804
rect 11885 31773 11897 31776
rect 11931 31804 11943 31807
rect 11931 31776 12020 31804
rect 11931 31773 11943 31776
rect 11885 31767 11943 31773
rect 8573 31671 8631 31677
rect 8573 31637 8585 31671
rect 8619 31637 8631 31671
rect 8573 31631 8631 31637
rect 10226 31628 10232 31680
rect 10284 31668 10290 31680
rect 11057 31671 11115 31677
rect 11057 31668 11069 31671
rect 10284 31640 11069 31668
rect 10284 31628 10290 31640
rect 11057 31637 11069 31640
rect 11103 31668 11115 31671
rect 11885 31671 11943 31677
rect 11885 31668 11897 31671
rect 11103 31640 11897 31668
rect 11103 31637 11115 31640
rect 11057 31631 11115 31637
rect 11885 31637 11897 31640
rect 11931 31668 11943 31671
rect 11992 31668 12020 31776
rect 12342 31764 12348 31816
rect 12400 31764 12406 31816
rect 13078 31764 13084 31816
rect 13136 31804 13142 31816
rect 13136 31776 14228 31804
rect 13136 31764 13142 31776
rect 14200 31736 14228 31776
rect 14274 31764 14280 31816
rect 14332 31764 14338 31816
rect 14936 31813 14964 31844
rect 14461 31807 14519 31813
rect 14461 31804 14473 31807
rect 14384 31776 14473 31804
rect 14384 31736 14412 31776
rect 14461 31773 14473 31776
rect 14507 31773 14519 31807
rect 14461 31767 14519 31773
rect 14921 31807 14979 31813
rect 14921 31773 14933 31807
rect 14967 31773 14979 31807
rect 14921 31767 14979 31773
rect 15102 31764 15108 31816
rect 15160 31764 15166 31816
rect 15580 31813 15608 31844
rect 15764 31813 15792 31912
rect 15565 31807 15623 31813
rect 15565 31773 15577 31807
rect 15611 31804 15623 31807
rect 15749 31807 15807 31813
rect 15611 31776 15700 31804
rect 15611 31773 15623 31776
rect 15565 31767 15623 31773
rect 14200 31708 14412 31736
rect 15672 31736 15700 31776
rect 15749 31773 15761 31807
rect 15795 31773 15807 31807
rect 16209 31807 16267 31813
rect 16209 31804 16221 31807
rect 15749 31767 15807 31773
rect 15856 31776 16221 31804
rect 15856 31736 15884 31776
rect 16209 31773 16221 31776
rect 16255 31773 16267 31807
rect 16209 31767 16267 31773
rect 16390 31764 16396 31816
rect 16448 31764 16454 31816
rect 15672 31708 15884 31736
rect 11931 31640 12020 31668
rect 11931 31637 11943 31640
rect 11885 31631 11943 31637
rect 12158 31628 12164 31680
rect 12216 31668 12222 31680
rect 12529 31671 12587 31677
rect 12529 31668 12541 31671
rect 12216 31640 12541 31668
rect 12216 31628 12222 31640
rect 12529 31637 12541 31640
rect 12575 31637 12587 31671
rect 12529 31631 12587 31637
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 5074 31424 5080 31476
rect 5132 31464 5138 31476
rect 5169 31467 5227 31473
rect 5169 31464 5181 31467
rect 5132 31436 5181 31464
rect 5132 31424 5138 31436
rect 5169 31433 5181 31436
rect 5215 31464 5227 31467
rect 5902 31464 5908 31476
rect 5215 31436 5908 31464
rect 5215 31433 5227 31436
rect 5169 31427 5227 31433
rect 5902 31424 5908 31436
rect 5960 31464 5966 31476
rect 5997 31467 6055 31473
rect 5997 31464 6009 31467
rect 5960 31436 6009 31464
rect 5960 31424 5966 31436
rect 5997 31433 6009 31436
rect 6043 31464 6055 31467
rect 6914 31464 6920 31476
rect 6043 31436 6920 31464
rect 6043 31433 6055 31436
rect 5997 31427 6055 31433
rect 6914 31424 6920 31436
rect 6972 31464 6978 31476
rect 7469 31467 7527 31473
rect 7469 31464 7481 31467
rect 6972 31436 7481 31464
rect 6972 31424 6978 31436
rect 7469 31433 7481 31436
rect 7515 31433 7527 31467
rect 7469 31427 7527 31433
rect 8297 31467 8355 31473
rect 8297 31433 8309 31467
rect 8343 31433 8355 31467
rect 8297 31427 8355 31433
rect 9125 31467 9183 31473
rect 9125 31433 9137 31467
rect 9171 31464 9183 31467
rect 10226 31464 10232 31476
rect 9171 31436 10232 31464
rect 9171 31433 9183 31436
rect 9125 31427 9183 31433
rect 1486 31288 1492 31340
rect 1544 31328 1550 31340
rect 1765 31331 1823 31337
rect 1765 31328 1777 31331
rect 1544 31300 1777 31328
rect 1544 31288 1550 31300
rect 1765 31297 1777 31300
rect 1811 31297 1823 31331
rect 1765 31291 1823 31297
rect 2038 31288 2044 31340
rect 2096 31288 2102 31340
rect 2590 31288 2596 31340
rect 2648 31288 2654 31340
rect 4798 31288 4804 31340
rect 4856 31328 4862 31340
rect 5629 31331 5687 31337
rect 5629 31328 5641 31331
rect 4856 31300 5641 31328
rect 4856 31288 4862 31300
rect 5629 31297 5641 31300
rect 5675 31328 5687 31331
rect 6546 31328 6552 31340
rect 5675 31300 6552 31328
rect 5675 31297 5687 31300
rect 5629 31291 5687 31297
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 7484 31337 7512 31427
rect 7469 31331 7527 31337
rect 7469 31297 7481 31331
rect 7515 31328 7527 31331
rect 7650 31328 7656 31340
rect 7515 31300 7656 31328
rect 7515 31297 7527 31300
rect 7469 31291 7527 31297
rect 7650 31288 7656 31300
rect 7708 31328 7714 31340
rect 8312 31337 8340 31427
rect 9140 31337 9168 31427
rect 10226 31424 10232 31436
rect 10284 31464 10290 31476
rect 10321 31467 10379 31473
rect 10321 31464 10333 31467
rect 10284 31436 10333 31464
rect 10284 31424 10290 31436
rect 10321 31433 10333 31436
rect 10367 31464 10379 31467
rect 11146 31464 11152 31476
rect 10367 31436 11152 31464
rect 10367 31433 10379 31436
rect 10321 31427 10379 31433
rect 10336 31337 10364 31427
rect 11146 31424 11152 31436
rect 11204 31464 11210 31476
rect 12066 31464 12072 31476
rect 11204 31436 12072 31464
rect 11204 31424 11210 31436
rect 12066 31424 12072 31436
rect 12124 31424 12130 31476
rect 13722 31424 13728 31476
rect 13780 31464 13786 31476
rect 14093 31467 14151 31473
rect 14093 31464 14105 31467
rect 13780 31436 14105 31464
rect 13780 31424 13786 31436
rect 14093 31433 14105 31436
rect 14139 31464 14151 31467
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 14139 31436 14933 31464
rect 14139 31433 14151 31436
rect 14093 31427 14151 31433
rect 14921 31433 14933 31436
rect 14967 31433 14979 31467
rect 14921 31427 14979 31433
rect 11054 31396 11060 31408
rect 10796 31368 11060 31396
rect 10796 31337 10824 31368
rect 11054 31356 11060 31368
rect 11112 31396 11118 31408
rect 12342 31396 12348 31408
rect 11112 31368 12348 31396
rect 11112 31356 11118 31368
rect 12342 31356 12348 31368
rect 12400 31356 12406 31408
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 7708 31300 8309 31328
rect 7708 31288 7714 31300
rect 8297 31297 8309 31300
rect 8343 31328 8355 31331
rect 9125 31331 9183 31337
rect 9125 31328 9137 31331
rect 8343 31300 9137 31328
rect 8343 31297 8355 31300
rect 8297 31291 8355 31297
rect 9125 31297 9137 31300
rect 9171 31297 9183 31331
rect 9125 31291 9183 31297
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 10781 31331 10839 31337
rect 10781 31297 10793 31331
rect 10827 31297 10839 31331
rect 10781 31291 10839 31297
rect 11146 31288 11152 31340
rect 11204 31288 11210 31340
rect 11974 31288 11980 31340
rect 12032 31328 12038 31340
rect 13081 31331 13139 31337
rect 13081 31328 13093 31331
rect 12032 31300 13093 31328
rect 12032 31288 12038 31300
rect 13081 31297 13093 31300
rect 13127 31297 13139 31331
rect 13081 31291 13139 31297
rect 2133 31263 2191 31269
rect 2133 31229 2145 31263
rect 2179 31260 2191 31263
rect 3878 31260 3884 31272
rect 2179 31232 3884 31260
rect 2179 31229 2191 31232
rect 2133 31223 2191 31229
rect 3878 31220 3884 31232
rect 3936 31220 3942 31272
rect 7101 31263 7159 31269
rect 7101 31229 7113 31263
rect 7147 31260 7159 31263
rect 7558 31260 7564 31272
rect 7147 31232 7564 31260
rect 7147 31229 7159 31232
rect 7101 31223 7159 31229
rect 7558 31220 7564 31232
rect 7616 31260 7622 31272
rect 7929 31263 7987 31269
rect 7929 31260 7941 31263
rect 7616 31232 7941 31260
rect 7616 31220 7622 31232
rect 7929 31229 7941 31232
rect 7975 31260 7987 31263
rect 8757 31263 8815 31269
rect 8757 31260 8769 31263
rect 7975 31232 8769 31260
rect 7975 31229 7987 31232
rect 7929 31223 7987 31229
rect 8757 31229 8769 31232
rect 8803 31229 8815 31263
rect 8757 31223 8815 31229
rect 9950 31220 9956 31272
rect 10008 31260 10014 31272
rect 11514 31260 11520 31272
rect 10008 31232 11520 31260
rect 10008 31220 10014 31232
rect 11514 31220 11520 31232
rect 11572 31260 11578 31272
rect 11701 31263 11759 31269
rect 11701 31260 11713 31263
rect 11572 31232 11713 31260
rect 11572 31220 11578 31232
rect 11701 31229 11713 31232
rect 11747 31260 11759 31263
rect 12158 31260 12164 31272
rect 11747 31232 12164 31260
rect 11747 31229 11759 31232
rect 11701 31223 11759 31229
rect 12158 31220 12164 31232
rect 12216 31220 12222 31272
rect 13170 31220 13176 31272
rect 13228 31260 13234 31272
rect 13725 31263 13783 31269
rect 13725 31260 13737 31263
rect 13228 31232 13737 31260
rect 13228 31220 13234 31232
rect 13725 31229 13737 31232
rect 13771 31229 13783 31263
rect 14553 31263 14611 31269
rect 14553 31260 14565 31263
rect 13725 31223 13783 31229
rect 14016 31232 14565 31260
rect 5166 31152 5172 31204
rect 5224 31192 5230 31204
rect 5902 31192 5908 31204
rect 5224 31164 5908 31192
rect 5224 31152 5230 31164
rect 5902 31152 5908 31164
rect 5960 31192 5966 31204
rect 5997 31195 6055 31201
rect 5997 31192 6009 31195
rect 5960 31164 6009 31192
rect 5960 31152 5966 31164
rect 5997 31161 6009 31164
rect 6043 31161 6055 31195
rect 5997 31155 6055 31161
rect 12066 31152 12072 31204
rect 12124 31152 12130 31204
rect 14016 31136 14044 31232
rect 14553 31229 14565 31232
rect 14599 31229 14611 31263
rect 14553 31223 14611 31229
rect 14093 31195 14151 31201
rect 14093 31161 14105 31195
rect 14139 31192 14151 31195
rect 14366 31192 14372 31204
rect 14139 31164 14372 31192
rect 14139 31161 14151 31164
rect 14093 31155 14151 31161
rect 14366 31152 14372 31164
rect 14424 31152 14430 31204
rect 14921 31195 14979 31201
rect 14921 31161 14933 31195
rect 14967 31192 14979 31195
rect 15194 31192 15200 31204
rect 14967 31164 15200 31192
rect 14967 31161 14979 31164
rect 14921 31155 14979 31161
rect 15194 31152 15200 31164
rect 15252 31152 15258 31204
rect 3786 31084 3792 31136
rect 3844 31124 3850 31136
rect 3881 31127 3939 31133
rect 3881 31124 3893 31127
rect 3844 31096 3893 31124
rect 3844 31084 3850 31096
rect 3881 31093 3893 31096
rect 3927 31093 3939 31127
rect 3881 31087 3939 31093
rect 4246 31084 4252 31136
rect 4304 31124 4310 31136
rect 4430 31124 4436 31136
rect 4304 31096 4436 31124
rect 4304 31084 4310 31096
rect 4430 31084 4436 31096
rect 4488 31124 4494 31136
rect 6362 31124 6368 31136
rect 4488 31096 6368 31124
rect 4488 31084 4494 31096
rect 6362 31084 6368 31096
rect 6420 31084 6426 31136
rect 12618 31084 12624 31136
rect 12676 31124 12682 31136
rect 13173 31127 13231 31133
rect 13173 31124 13185 31127
rect 12676 31096 13185 31124
rect 12676 31084 12682 31096
rect 13173 31093 13185 31096
rect 13219 31124 13231 31127
rect 13998 31124 14004 31136
rect 13219 31096 14004 31124
rect 13219 31093 13231 31096
rect 13173 31087 13231 31093
rect 13998 31084 14004 31096
rect 14056 31084 14062 31136
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 2590 30920 2596 30932
rect 1688 30892 2596 30920
rect 1688 30725 1716 30892
rect 2590 30880 2596 30892
rect 2648 30920 2654 30932
rect 6273 30923 6331 30929
rect 6273 30920 6285 30923
rect 2648 30892 6285 30920
rect 2648 30880 2654 30892
rect 6273 30889 6285 30892
rect 6319 30889 6331 30923
rect 6273 30883 6331 30889
rect 7650 30880 7656 30932
rect 7708 30920 7714 30932
rect 8573 30923 8631 30929
rect 8573 30920 8585 30923
rect 7708 30892 8585 30920
rect 7708 30880 7714 30892
rect 8573 30889 8585 30892
rect 8619 30889 8631 30923
rect 8573 30883 8631 30889
rect 8294 30852 8300 30864
rect 3436 30824 8300 30852
rect 3436 30793 3464 30824
rect 8294 30812 8300 30824
rect 8352 30812 8358 30864
rect 8588 30852 8616 30883
rect 12066 30880 12072 30932
rect 12124 30920 12130 30932
rect 12161 30923 12219 30929
rect 12161 30920 12173 30923
rect 12124 30892 12173 30920
rect 12124 30880 12130 30892
rect 12161 30889 12173 30892
rect 12207 30889 12219 30923
rect 12161 30883 12219 30889
rect 9582 30852 9588 30864
rect 8588 30824 9588 30852
rect 3421 30787 3479 30793
rect 3421 30753 3433 30787
rect 3467 30753 3479 30787
rect 3421 30747 3479 30753
rect 4065 30787 4123 30793
rect 4065 30753 4077 30787
rect 4111 30784 4123 30787
rect 5626 30784 5632 30796
rect 4111 30756 5632 30784
rect 4111 30753 4123 30756
rect 4065 30747 4123 30753
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 7558 30744 7564 30796
rect 7616 30784 7622 30796
rect 8588 30793 8616 30824
rect 9582 30812 9588 30824
rect 9640 30852 9646 30864
rect 9677 30855 9735 30861
rect 9677 30852 9689 30855
rect 9640 30824 9689 30852
rect 9640 30812 9646 30824
rect 9677 30821 9689 30824
rect 9723 30852 9735 30855
rect 10505 30855 10563 30861
rect 10505 30852 10517 30855
rect 9723 30824 10517 30852
rect 9723 30821 9735 30824
rect 9677 30815 9735 30821
rect 10505 30821 10517 30824
rect 10551 30852 10563 30855
rect 11333 30855 11391 30861
rect 11333 30852 11345 30855
rect 10551 30824 11345 30852
rect 10551 30821 10563 30824
rect 10505 30815 10563 30821
rect 11333 30821 11345 30824
rect 11379 30821 11391 30855
rect 11333 30815 11391 30821
rect 8205 30787 8263 30793
rect 8205 30784 8217 30787
rect 7616 30756 8217 30784
rect 7616 30744 7622 30756
rect 8205 30753 8217 30756
rect 8251 30753 8263 30787
rect 8205 30747 8263 30753
rect 8573 30787 8631 30793
rect 8573 30753 8585 30787
rect 8619 30753 8631 30787
rect 8573 30747 8631 30753
rect 9309 30787 9367 30793
rect 9309 30753 9321 30787
rect 9355 30784 9367 30787
rect 9950 30784 9956 30796
rect 9355 30756 9956 30784
rect 9355 30753 9367 30756
rect 9309 30747 9367 30753
rect 9950 30744 9956 30756
rect 10008 30744 10014 30796
rect 10137 30787 10195 30793
rect 10137 30753 10149 30787
rect 10183 30784 10195 30787
rect 10965 30787 11023 30793
rect 10965 30784 10977 30787
rect 10183 30756 10977 30784
rect 10183 30753 10195 30756
rect 10137 30747 10195 30753
rect 10965 30753 10977 30756
rect 11011 30784 11023 30787
rect 11054 30784 11060 30796
rect 11011 30756 11060 30784
rect 11011 30753 11023 30756
rect 10965 30747 11023 30753
rect 11054 30744 11060 30756
rect 11112 30784 11118 30796
rect 12176 30793 12204 30883
rect 11793 30787 11851 30793
rect 11793 30784 11805 30787
rect 11112 30756 11805 30784
rect 11112 30744 11118 30756
rect 11793 30753 11805 30756
rect 11839 30753 11851 30787
rect 11793 30747 11851 30753
rect 12161 30787 12219 30793
rect 12161 30753 12173 30787
rect 12207 30784 12219 30787
rect 13725 30787 13783 30793
rect 12207 30756 12434 30784
rect 12207 30753 12219 30756
rect 12161 30747 12219 30753
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 4246 30676 4252 30728
rect 4304 30676 4310 30728
rect 4338 30676 4344 30728
rect 4396 30716 4402 30728
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4396 30688 4997 30716
rect 4396 30676 4402 30688
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 4985 30679 5043 30685
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 7285 30719 7343 30725
rect 7285 30716 7297 30719
rect 6604 30688 7297 30716
rect 6604 30676 6610 30688
rect 7285 30685 7297 30688
rect 7331 30685 7343 30719
rect 7285 30679 7343 30685
rect 7650 30676 7656 30728
rect 7708 30676 7714 30728
rect 4525 30651 4583 30657
rect 4525 30617 4537 30651
rect 4571 30648 4583 30651
rect 5994 30648 6000 30660
rect 4571 30620 6000 30648
rect 4571 30617 4583 30620
rect 4525 30611 4583 30617
rect 5994 30608 6000 30620
rect 6052 30608 6058 30660
rect 4154 30540 4160 30592
rect 4212 30580 4218 30592
rect 4433 30583 4491 30589
rect 4433 30580 4445 30583
rect 4212 30552 4445 30580
rect 4212 30540 4218 30552
rect 4433 30549 4445 30552
rect 4479 30549 4491 30583
rect 4433 30543 4491 30549
rect 9582 30540 9588 30592
rect 9640 30580 9646 30592
rect 9677 30583 9735 30589
rect 9677 30580 9689 30583
rect 9640 30552 9689 30580
rect 9640 30540 9646 30552
rect 9677 30549 9689 30552
rect 9723 30580 9735 30583
rect 10505 30583 10563 30589
rect 10505 30580 10517 30583
rect 9723 30552 10517 30580
rect 9723 30549 9735 30552
rect 9677 30543 9735 30549
rect 10505 30549 10517 30552
rect 10551 30580 10563 30583
rect 11333 30583 11391 30589
rect 11333 30580 11345 30583
rect 10551 30552 11345 30580
rect 10551 30549 10563 30552
rect 10505 30543 10563 30549
rect 11333 30549 11345 30552
rect 11379 30549 11391 30583
rect 12406 30580 12434 30756
rect 13725 30753 13737 30787
rect 13771 30784 13783 30787
rect 14366 30784 14372 30796
rect 13771 30756 14372 30784
rect 13771 30753 13783 30756
rect 13725 30747 13783 30753
rect 14366 30744 14372 30756
rect 14424 30784 14430 30796
rect 15933 30787 15991 30793
rect 15933 30784 15945 30787
rect 14424 30756 15945 30784
rect 14424 30744 14430 30756
rect 15933 30753 15945 30756
rect 15979 30753 15991 30787
rect 15933 30747 15991 30753
rect 12618 30676 12624 30728
rect 12676 30676 12682 30728
rect 13170 30676 13176 30728
rect 13228 30716 13234 30728
rect 13357 30719 13415 30725
rect 13357 30716 13369 30719
rect 13228 30688 13369 30716
rect 13228 30676 13234 30688
rect 13357 30685 13369 30688
rect 13403 30685 13415 30719
rect 13357 30679 13415 30685
rect 13998 30676 14004 30728
rect 14056 30716 14062 30728
rect 14829 30719 14887 30725
rect 14829 30716 14841 30719
rect 14056 30688 14841 30716
rect 14056 30676 14062 30688
rect 14829 30685 14841 30688
rect 14875 30685 14887 30719
rect 14829 30679 14887 30685
rect 15194 30676 15200 30728
rect 15252 30676 15258 30728
rect 13262 30608 13268 30660
rect 13320 30648 13326 30660
rect 15749 30651 15807 30657
rect 15749 30648 15761 30651
rect 13320 30620 15761 30648
rect 13320 30608 13326 30620
rect 15749 30617 15761 30620
rect 15795 30617 15807 30651
rect 15749 30611 15807 30617
rect 12710 30580 12716 30592
rect 12406 30552 12716 30580
rect 11333 30543 11391 30549
rect 12710 30540 12716 30552
rect 12768 30540 12774 30592
rect 12805 30583 12863 30589
rect 12805 30549 12817 30583
rect 12851 30580 12863 30583
rect 13170 30580 13176 30592
rect 12851 30552 13176 30580
rect 12851 30549 12863 30552
rect 12805 30543 12863 30549
rect 13170 30540 13176 30552
rect 13228 30540 13234 30592
rect 13722 30540 13728 30592
rect 13780 30580 13786 30592
rect 15197 30583 15255 30589
rect 15197 30580 15209 30583
rect 13780 30552 15209 30580
rect 13780 30540 13786 30552
rect 15197 30549 15209 30552
rect 15243 30549 15255 30583
rect 15197 30543 15255 30549
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 6914 30336 6920 30388
rect 6972 30376 6978 30388
rect 7745 30379 7803 30385
rect 7745 30376 7757 30379
rect 6972 30348 7757 30376
rect 6972 30336 6978 30348
rect 7745 30345 7757 30348
rect 7791 30376 7803 30379
rect 9125 30379 9183 30385
rect 9125 30376 9137 30379
rect 7791 30348 9137 30376
rect 7791 30345 7803 30348
rect 7745 30339 7803 30345
rect 9125 30345 9137 30348
rect 9171 30376 9183 30379
rect 10321 30379 10379 30385
rect 10321 30376 10333 30379
rect 9171 30348 10333 30376
rect 9171 30345 9183 30348
rect 9125 30339 9183 30345
rect 10321 30345 10333 30348
rect 10367 30376 10379 30379
rect 11149 30379 11207 30385
rect 11149 30376 11161 30379
rect 10367 30348 11161 30376
rect 10367 30345 10379 30348
rect 10321 30339 10379 30345
rect 11149 30345 11161 30348
rect 11195 30345 11207 30379
rect 11149 30339 11207 30345
rect 1854 30268 1860 30320
rect 1912 30308 1918 30320
rect 2041 30311 2099 30317
rect 2041 30308 2053 30311
rect 1912 30280 2053 30308
rect 1912 30268 1918 30280
rect 2041 30277 2053 30280
rect 2087 30277 2099 30311
rect 2041 30271 2099 30277
rect 3970 30268 3976 30320
rect 4028 30308 4034 30320
rect 5169 30311 5227 30317
rect 5169 30308 5181 30311
rect 4028 30280 5181 30308
rect 4028 30268 4034 30280
rect 5169 30277 5181 30280
rect 5215 30277 5227 30311
rect 7466 30308 7472 30320
rect 5169 30271 5227 30277
rect 5368 30280 7472 30308
rect 1949 30243 2007 30249
rect 1949 30209 1961 30243
rect 1995 30209 2007 30243
rect 1949 30203 2007 30209
rect 1964 30172 1992 30203
rect 2130 30200 2136 30252
rect 2188 30200 2194 30252
rect 2222 30200 2228 30252
rect 2280 30200 2286 30252
rect 2406 30200 2412 30252
rect 2464 30200 2470 30252
rect 2866 30200 2872 30252
rect 2924 30200 2930 30252
rect 5368 30249 5396 30280
rect 7466 30268 7472 30280
rect 7524 30268 7530 30320
rect 5353 30243 5411 30249
rect 5353 30209 5365 30243
rect 5399 30209 5411 30243
rect 5353 30203 5411 30209
rect 5442 30200 5448 30252
rect 5500 30200 5506 30252
rect 6178 30240 6184 30252
rect 5552 30212 6184 30240
rect 5552 30172 5580 30212
rect 6178 30200 6184 30212
rect 6236 30200 6242 30252
rect 6546 30200 6552 30252
rect 6604 30240 6610 30252
rect 7377 30243 7435 30249
rect 7377 30240 7389 30243
rect 6604 30212 7389 30240
rect 6604 30200 6610 30212
rect 7377 30209 7389 30212
rect 7423 30209 7435 30243
rect 7377 30203 7435 30209
rect 7558 30200 7564 30252
rect 7616 30240 7622 30252
rect 9140 30249 9168 30339
rect 8757 30243 8815 30249
rect 8757 30240 8769 30243
rect 7616 30212 8769 30240
rect 7616 30200 7622 30212
rect 8757 30209 8769 30212
rect 8803 30209 8815 30243
rect 8757 30203 8815 30209
rect 9125 30243 9183 30249
rect 9125 30209 9137 30243
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 9950 30200 9956 30252
rect 10008 30200 10014 30252
rect 10336 30249 10364 30339
rect 10321 30243 10379 30249
rect 10321 30209 10333 30243
rect 10367 30209 10379 30243
rect 10321 30203 10379 30209
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 11054 30240 11060 30252
rect 10827 30212 11060 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 11054 30200 11060 30212
rect 11112 30200 11118 30252
rect 11164 30249 11192 30339
rect 12710 30336 12716 30388
rect 12768 30376 12774 30388
rect 13541 30379 13599 30385
rect 13541 30376 13553 30379
rect 12768 30348 13553 30376
rect 12768 30336 12774 30348
rect 13541 30345 13553 30348
rect 13587 30376 13599 30379
rect 13722 30376 13728 30388
rect 13587 30348 13728 30376
rect 13587 30345 13599 30348
rect 13541 30339 13599 30345
rect 13722 30336 13728 30348
rect 13780 30376 13786 30388
rect 14369 30379 14427 30385
rect 14369 30376 14381 30379
rect 13780 30348 14381 30376
rect 13780 30336 13786 30348
rect 14369 30345 14381 30348
rect 14415 30376 14427 30379
rect 15197 30379 15255 30385
rect 15197 30376 15209 30379
rect 14415 30348 15209 30376
rect 14415 30345 14427 30348
rect 14369 30339 14427 30345
rect 15197 30345 15209 30348
rect 15243 30376 15255 30379
rect 16025 30379 16083 30385
rect 16025 30376 16037 30379
rect 15243 30348 16037 30376
rect 15243 30345 15255 30348
rect 15197 30339 15255 30345
rect 16025 30345 16037 30348
rect 16071 30345 16083 30379
rect 16025 30339 16083 30345
rect 11149 30243 11207 30249
rect 11149 30209 11161 30243
rect 11195 30209 11207 30243
rect 11149 30203 11207 30209
rect 11698 30200 11704 30252
rect 11756 30200 11762 30252
rect 11882 30200 11888 30252
rect 11940 30200 11946 30252
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14826 30240 14832 30252
rect 14056 30212 14832 30240
rect 14056 30200 14062 30212
rect 14826 30200 14832 30212
rect 14884 30240 14890 30252
rect 15657 30243 15715 30249
rect 15657 30240 15669 30243
rect 14884 30212 15669 30240
rect 14884 30200 14890 30212
rect 15657 30209 15669 30212
rect 15703 30209 15715 30243
rect 15657 30203 15715 30209
rect 1964 30144 5580 30172
rect 5626 30132 5632 30184
rect 5684 30132 5690 30184
rect 5721 30175 5779 30181
rect 5721 30141 5733 30175
rect 5767 30141 5779 30175
rect 5721 30135 5779 30141
rect 12345 30175 12403 30181
rect 12345 30141 12357 30175
rect 12391 30172 12403 30175
rect 13170 30172 13176 30184
rect 12391 30144 13176 30172
rect 12391 30141 12403 30144
rect 12345 30135 12403 30141
rect 1765 30107 1823 30113
rect 1765 30073 1777 30107
rect 1811 30104 1823 30107
rect 4338 30104 4344 30116
rect 1811 30076 4344 30104
rect 1811 30073 1823 30076
rect 1765 30067 1823 30073
rect 4338 30064 4344 30076
rect 4396 30064 4402 30116
rect 5074 30064 5080 30116
rect 5132 30104 5138 30116
rect 5736 30104 5764 30135
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 14366 30172 14372 30184
rect 13464 30144 14372 30172
rect 5132 30076 5764 30104
rect 5132 30064 5138 30076
rect 6914 30064 6920 30116
rect 6972 30104 6978 30116
rect 7650 30104 7656 30116
rect 6972 30076 7656 30104
rect 6972 30064 6978 30076
rect 7650 30064 7656 30076
rect 7708 30104 7714 30116
rect 7745 30107 7803 30113
rect 7745 30104 7757 30107
rect 7708 30076 7757 30104
rect 7708 30064 7714 30076
rect 7745 30073 7757 30076
rect 7791 30073 7803 30107
rect 7745 30067 7803 30073
rect 12713 30107 12771 30113
rect 12713 30073 12725 30107
rect 12759 30104 12771 30107
rect 12894 30104 12900 30116
rect 12759 30076 12900 30104
rect 12759 30073 12771 30076
rect 12713 30067 12771 30073
rect 12894 30064 12900 30076
rect 12952 30104 12958 30116
rect 13464 30104 13492 30144
rect 14366 30132 14372 30144
rect 14424 30132 14430 30184
rect 12952 30076 13492 30104
rect 13541 30107 13599 30113
rect 12952 30064 12958 30076
rect 13541 30073 13553 30107
rect 13587 30104 13599 30107
rect 13814 30104 13820 30116
rect 13587 30076 13820 30104
rect 13587 30073 13599 30076
rect 13541 30067 13599 30073
rect 13814 30064 13820 30076
rect 13872 30064 13878 30116
rect 15194 30064 15200 30116
rect 15252 30104 15258 30116
rect 16025 30107 16083 30113
rect 16025 30104 16037 30107
rect 15252 30076 16037 30104
rect 15252 30064 15258 30076
rect 16025 30073 16037 30076
rect 16071 30073 16083 30107
rect 16025 30067 16083 30073
rect 1578 29996 1584 30048
rect 1636 30036 1642 30048
rect 2498 30036 2504 30048
rect 1636 30008 2504 30036
rect 1636 29996 1642 30008
rect 2498 29996 2504 30008
rect 2556 30036 2562 30048
rect 4157 30039 4215 30045
rect 4157 30036 4169 30039
rect 2556 30008 4169 30036
rect 2556 29996 2562 30008
rect 4157 30005 4169 30008
rect 4203 30005 4215 30039
rect 4157 29999 4215 30005
rect 4246 29996 4252 30048
rect 4304 30036 4310 30048
rect 10410 30036 10416 30048
rect 4304 30008 10416 30036
rect 4304 29996 4310 30008
rect 10410 29996 10416 30008
rect 10468 29996 10474 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 5166 29792 5172 29844
rect 5224 29832 5230 29844
rect 5445 29835 5503 29841
rect 5445 29832 5457 29835
rect 5224 29804 5457 29832
rect 5224 29792 5230 29804
rect 5445 29801 5457 29804
rect 5491 29801 5503 29835
rect 7374 29832 7380 29844
rect 5445 29795 5503 29801
rect 5828 29804 7380 29832
rect 2222 29724 2228 29776
rect 2280 29764 2286 29776
rect 4246 29764 4252 29776
rect 2280 29736 4252 29764
rect 2280 29724 2286 29736
rect 4246 29724 4252 29736
rect 4304 29724 4310 29776
rect 5828 29764 5856 29804
rect 7374 29792 7380 29804
rect 7432 29792 7438 29844
rect 9309 29835 9367 29841
rect 9309 29801 9321 29835
rect 9355 29832 9367 29835
rect 14458 29832 14464 29844
rect 9355 29804 14464 29832
rect 9355 29801 9367 29804
rect 9309 29795 9367 29801
rect 14458 29792 14464 29804
rect 14516 29792 14522 29844
rect 4540 29736 5856 29764
rect 1688 29668 4476 29696
rect 1688 29637 1716 29668
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 1946 29588 1952 29640
rect 2004 29628 2010 29640
rect 2406 29628 2412 29640
rect 2004 29600 2412 29628
rect 2004 29588 2010 29600
rect 2406 29588 2412 29600
rect 2464 29628 2470 29640
rect 3973 29631 4031 29637
rect 3973 29628 3985 29631
rect 2464 29600 3985 29628
rect 2464 29588 2470 29600
rect 3973 29597 3985 29600
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 4246 29588 4252 29640
rect 4304 29588 4310 29640
rect 3878 29520 3884 29572
rect 3936 29560 3942 29572
rect 4448 29560 4476 29668
rect 4540 29637 4568 29736
rect 5902 29724 5908 29776
rect 5960 29764 5966 29776
rect 6549 29767 6607 29773
rect 6549 29764 6561 29767
rect 5960 29736 6561 29764
rect 5960 29724 5966 29736
rect 6549 29733 6561 29736
rect 6595 29764 6607 29767
rect 6914 29764 6920 29776
rect 6595 29736 6920 29764
rect 6595 29733 6607 29736
rect 6549 29727 6607 29733
rect 6914 29724 6920 29736
rect 6972 29724 6978 29776
rect 11054 29724 11060 29776
rect 11112 29764 11118 29776
rect 11885 29767 11943 29773
rect 11885 29764 11897 29767
rect 11112 29736 11897 29764
rect 11112 29724 11118 29736
rect 11885 29733 11897 29736
rect 11931 29733 11943 29767
rect 11885 29727 11943 29733
rect 12894 29724 12900 29776
rect 12952 29724 12958 29776
rect 8435 29699 8493 29705
rect 8435 29696 8447 29699
rect 4632 29668 8447 29696
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29597 4583 29631
rect 4525 29591 4583 29597
rect 4632 29560 4660 29668
rect 8435 29665 8447 29668
rect 8481 29665 8493 29699
rect 8435 29659 8493 29665
rect 9950 29656 9956 29708
rect 10008 29696 10014 29708
rect 10686 29696 10692 29708
rect 10008 29668 10692 29696
rect 10008 29656 10014 29668
rect 10686 29656 10692 29668
rect 10744 29696 10750 29708
rect 10781 29699 10839 29705
rect 10781 29696 10793 29699
rect 10744 29668 10793 29696
rect 10744 29656 10750 29668
rect 10781 29665 10793 29668
rect 10827 29665 10839 29699
rect 10781 29659 10839 29665
rect 14826 29656 14832 29708
rect 14884 29656 14890 29708
rect 16025 29699 16083 29705
rect 16025 29696 16037 29699
rect 15212 29668 16037 29696
rect 15212 29640 15240 29668
rect 16025 29665 16037 29668
rect 16071 29665 16083 29699
rect 16025 29659 16083 29665
rect 4801 29631 4859 29637
rect 4801 29597 4813 29631
rect 4847 29628 4859 29631
rect 5534 29628 5540 29640
rect 4847 29600 5540 29628
rect 4847 29597 4859 29600
rect 4801 29591 4859 29597
rect 5534 29588 5540 29600
rect 5592 29588 5598 29640
rect 6181 29631 6239 29637
rect 6181 29597 6193 29631
rect 6227 29628 6239 29631
rect 6454 29628 6460 29640
rect 6227 29600 6460 29628
rect 6227 29597 6239 29600
rect 6181 29591 6239 29597
rect 6454 29588 6460 29600
rect 6512 29588 6518 29640
rect 7466 29588 7472 29640
rect 7524 29588 7530 29640
rect 7558 29588 7564 29640
rect 7616 29628 7622 29640
rect 7653 29631 7711 29637
rect 7653 29628 7665 29631
rect 7616 29600 7665 29628
rect 7616 29588 7622 29600
rect 7653 29597 7665 29600
rect 7699 29597 7711 29631
rect 7653 29591 7711 29597
rect 8294 29588 8300 29640
rect 8352 29637 8358 29640
rect 8352 29631 8390 29637
rect 8378 29597 8390 29631
rect 8352 29591 8390 29597
rect 10321 29631 10379 29637
rect 10321 29597 10333 29631
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29628 11207 29631
rect 12529 29631 12587 29637
rect 11195 29600 12434 29628
rect 11195 29597 11207 29600
rect 11149 29591 11207 29597
rect 8352 29588 8358 29591
rect 3936 29532 4200 29560
rect 4448 29532 4660 29560
rect 5261 29563 5319 29569
rect 3936 29520 3942 29532
rect 1578 29452 1584 29504
rect 1636 29492 1642 29504
rect 2961 29495 3019 29501
rect 2961 29492 2973 29495
rect 1636 29464 2973 29492
rect 1636 29452 1642 29464
rect 2961 29461 2973 29464
rect 3007 29461 3019 29495
rect 2961 29455 3019 29461
rect 3418 29452 3424 29504
rect 3476 29492 3482 29504
rect 4065 29495 4123 29501
rect 4065 29492 4077 29495
rect 3476 29464 4077 29492
rect 3476 29452 3482 29464
rect 4065 29461 4077 29464
rect 4111 29461 4123 29495
rect 4172 29492 4200 29532
rect 5261 29529 5273 29563
rect 5307 29560 5319 29563
rect 5810 29560 5816 29572
rect 5307 29532 5816 29560
rect 5307 29529 5319 29532
rect 5261 29523 5319 29529
rect 5810 29520 5816 29532
rect 5868 29520 5874 29572
rect 6472 29560 6500 29588
rect 6472 29532 7604 29560
rect 5445 29495 5503 29501
rect 5445 29492 5457 29495
rect 4172 29464 5457 29492
rect 4065 29455 4123 29461
rect 5445 29461 5457 29464
rect 5491 29461 5503 29495
rect 5445 29455 5503 29461
rect 5626 29452 5632 29504
rect 5684 29452 5690 29504
rect 6549 29495 6607 29501
rect 6549 29461 6561 29495
rect 6595 29492 6607 29495
rect 6822 29492 6828 29504
rect 6595 29464 6828 29492
rect 6595 29461 6607 29464
rect 6549 29455 6607 29461
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 7576 29501 7604 29532
rect 10336 29501 10364 29591
rect 7561 29495 7619 29501
rect 7561 29461 7573 29495
rect 7607 29461 7619 29495
rect 7561 29455 7619 29461
rect 10321 29495 10379 29501
rect 10321 29461 10333 29495
rect 10367 29492 10379 29495
rect 11054 29492 11060 29504
rect 10367 29464 11060 29492
rect 10367 29461 10379 29464
rect 10321 29455 10379 29461
rect 11054 29452 11060 29464
rect 11112 29492 11118 29504
rect 11164 29501 11192 29591
rect 11701 29563 11759 29569
rect 11701 29529 11713 29563
rect 11747 29560 11759 29563
rect 11882 29560 11888 29572
rect 11747 29532 11888 29560
rect 11747 29529 11759 29532
rect 11701 29523 11759 29529
rect 11882 29520 11888 29532
rect 11940 29520 11946 29572
rect 11149 29495 11207 29501
rect 11149 29492 11161 29495
rect 11112 29464 11161 29492
rect 11112 29452 11118 29464
rect 11149 29461 11161 29464
rect 11195 29461 11207 29495
rect 12406 29492 12434 29600
rect 12529 29597 12541 29631
rect 12575 29628 12587 29631
rect 13170 29628 13176 29640
rect 12575 29600 13176 29628
rect 12575 29597 12587 29600
rect 12529 29591 12587 29597
rect 13170 29588 13176 29600
rect 13228 29628 13234 29640
rect 13357 29631 13415 29637
rect 13357 29628 13369 29631
rect 13228 29600 13369 29628
rect 13228 29588 13234 29600
rect 13357 29597 13369 29600
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 13814 29628 13820 29640
rect 13771 29600 13820 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 13372 29560 13400 29591
rect 13814 29588 13820 29600
rect 13872 29588 13878 29640
rect 15194 29588 15200 29640
rect 15252 29588 15258 29640
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29597 15715 29631
rect 15657 29591 15715 29597
rect 14182 29560 14188 29572
rect 13372 29532 14188 29560
rect 14182 29520 14188 29532
rect 14240 29560 14246 29572
rect 15672 29560 15700 29591
rect 14240 29532 15700 29560
rect 14240 29520 14246 29532
rect 12710 29492 12716 29504
rect 12406 29464 12716 29492
rect 11149 29455 11207 29461
rect 12710 29452 12716 29464
rect 12768 29492 12774 29504
rect 12897 29495 12955 29501
rect 12897 29492 12909 29495
rect 12768 29464 12909 29492
rect 12768 29452 12774 29464
rect 12897 29461 12909 29464
rect 12943 29492 12955 29495
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 12943 29464 13737 29492
rect 12943 29461 12955 29464
rect 12897 29455 12955 29461
rect 13725 29461 13737 29464
rect 13771 29492 13783 29495
rect 15197 29495 15255 29501
rect 15197 29492 15209 29495
rect 13771 29464 15209 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 15197 29461 15209 29464
rect 15243 29492 15255 29495
rect 16025 29495 16083 29501
rect 16025 29492 16037 29495
rect 15243 29464 16037 29492
rect 15243 29461 15255 29464
rect 15197 29455 15255 29461
rect 16025 29461 16037 29464
rect 16071 29461 16083 29495
rect 16025 29455 16083 29461
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 1762 29248 1768 29300
rect 1820 29288 1826 29300
rect 1820 29260 2774 29288
rect 1820 29248 1826 29260
rect 2406 29220 2412 29232
rect 1872 29192 2412 29220
rect 1872 29161 1900 29192
rect 2406 29180 2412 29192
rect 2464 29180 2470 29232
rect 2746 29220 2774 29260
rect 2866 29248 2872 29300
rect 2924 29288 2930 29300
rect 9953 29291 10011 29297
rect 9953 29288 9965 29291
rect 2924 29260 9965 29288
rect 2924 29248 2930 29260
rect 9953 29257 9965 29260
rect 9999 29257 10011 29291
rect 9953 29251 10011 29257
rect 11054 29248 11060 29300
rect 11112 29248 11118 29300
rect 16390 29288 16396 29300
rect 13832 29260 16396 29288
rect 5261 29223 5319 29229
rect 5261 29220 5273 29223
rect 2746 29192 5273 29220
rect 5261 29189 5273 29192
rect 5307 29189 5319 29223
rect 5261 29183 5319 29189
rect 5626 29180 5632 29232
rect 5684 29220 5690 29232
rect 13832 29220 13860 29260
rect 16390 29248 16396 29260
rect 16448 29248 16454 29300
rect 5684 29192 9812 29220
rect 5684 29180 5690 29192
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29121 1915 29155
rect 1857 29115 1915 29121
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29121 2099 29155
rect 2041 29115 2099 29121
rect 2056 29016 2084 29115
rect 2590 29112 2596 29164
rect 2648 29112 2654 29164
rect 5442 29112 5448 29164
rect 5500 29112 5506 29164
rect 6914 29112 6920 29164
rect 6972 29112 6978 29164
rect 9784 29161 9812 29192
rect 10520 29192 13860 29220
rect 9769 29155 9827 29161
rect 9769 29121 9781 29155
rect 9815 29121 9827 29155
rect 9769 29115 9827 29121
rect 2133 29087 2191 29093
rect 2133 29053 2145 29087
rect 2179 29084 2191 29087
rect 3970 29084 3976 29096
rect 2179 29056 3976 29084
rect 2179 29053 2191 29056
rect 2133 29047 2191 29053
rect 3970 29044 3976 29056
rect 4028 29044 4034 29096
rect 4341 29087 4399 29093
rect 4341 29053 4353 29087
rect 4387 29053 4399 29087
rect 4341 29047 4399 29053
rect 5721 29087 5779 29093
rect 5721 29053 5733 29087
rect 5767 29084 5779 29087
rect 6730 29084 6736 29096
rect 5767 29056 6736 29084
rect 5767 29053 5779 29056
rect 5721 29047 5779 29053
rect 4356 29016 4384 29047
rect 6730 29044 6736 29056
rect 6788 29044 6794 29096
rect 7006 29044 7012 29096
rect 7064 29044 7070 29096
rect 7193 29087 7251 29093
rect 7193 29053 7205 29087
rect 7239 29053 7251 29087
rect 7193 29047 7251 29053
rect 8665 29087 8723 29093
rect 8665 29053 8677 29087
rect 8711 29084 8723 29087
rect 10520 29084 10548 29192
rect 14366 29180 14372 29232
rect 14424 29220 14430 29232
rect 14424 29192 15056 29220
rect 14424 29180 14430 29192
rect 10686 29112 10692 29164
rect 10744 29112 10750 29164
rect 11054 29112 11060 29164
rect 11112 29112 11118 29164
rect 11698 29112 11704 29164
rect 11756 29112 11762 29164
rect 11885 29155 11943 29161
rect 11885 29121 11897 29155
rect 11931 29121 11943 29155
rect 11885 29115 11943 29121
rect 13725 29155 13783 29161
rect 13725 29121 13737 29155
rect 13771 29152 13783 29155
rect 13814 29152 13820 29164
rect 13771 29124 13820 29152
rect 13771 29121 13783 29124
rect 13725 29115 13783 29121
rect 8711 29056 10548 29084
rect 8711 29053 8723 29056
rect 8665 29047 8723 29053
rect 5534 29016 5540 29028
rect 2056 28988 5540 29016
rect 5534 28976 5540 28988
rect 5592 29016 5598 29028
rect 6086 29016 6092 29028
rect 5592 28988 6092 29016
rect 5592 28976 5598 28988
rect 6086 28976 6092 28988
rect 6144 28976 6150 29028
rect 6196 28988 6776 29016
rect 5629 28951 5687 28957
rect 5629 28917 5641 28951
rect 5675 28948 5687 28951
rect 5718 28948 5724 28960
rect 5675 28920 5724 28948
rect 5675 28917 5687 28920
rect 5629 28911 5687 28917
rect 5718 28908 5724 28920
rect 5776 28948 5782 28960
rect 6196 28948 6224 28988
rect 5776 28920 6224 28948
rect 6549 28951 6607 28957
rect 5776 28908 5782 28920
rect 6549 28917 6561 28951
rect 6595 28948 6607 28951
rect 6638 28948 6644 28960
rect 6595 28920 6644 28948
rect 6595 28917 6607 28920
rect 6549 28911 6607 28917
rect 6638 28908 6644 28920
rect 6696 28908 6702 28960
rect 6748 28948 6776 28988
rect 7208 28948 7236 29047
rect 7650 28976 7656 29028
rect 7708 29016 7714 29028
rect 8021 29019 8079 29025
rect 8021 29016 8033 29019
rect 7708 28988 8033 29016
rect 7708 28976 7714 28988
rect 8021 28985 8033 28988
rect 8067 28985 8079 29019
rect 8021 28979 8079 28985
rect 9306 28976 9312 29028
rect 9364 28976 9370 29028
rect 10134 28976 10140 29028
rect 10192 29016 10198 29028
rect 11900 29016 11928 29115
rect 13814 29112 13820 29124
rect 13872 29152 13878 29164
rect 15028 29161 15056 29192
rect 14553 29155 14611 29161
rect 14553 29152 14565 29155
rect 13872 29124 14565 29152
rect 13872 29112 13878 29124
rect 14553 29121 14565 29124
rect 14599 29121 14611 29155
rect 14553 29115 14611 29121
rect 15013 29155 15071 29161
rect 15013 29121 15025 29155
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 12342 29044 12348 29096
rect 12400 29044 12406 29096
rect 12713 29087 12771 29093
rect 12713 29053 12725 29087
rect 12759 29053 12771 29087
rect 12713 29047 12771 29053
rect 13357 29087 13415 29093
rect 13357 29053 13369 29087
rect 13403 29084 13415 29087
rect 14182 29084 14188 29096
rect 13403 29056 14188 29084
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 10192 28988 11928 29016
rect 10192 28976 10198 28988
rect 12728 28960 12756 29047
rect 14182 29044 14188 29056
rect 14240 29044 14246 29096
rect 14568 29016 14596 29115
rect 15194 29016 15200 29028
rect 14568 28988 15200 29016
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 11054 28948 11060 28960
rect 6748 28920 11060 28948
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 12710 28908 12716 28960
rect 12768 28908 12774 28960
rect 13725 28951 13783 28957
rect 13725 28917 13737 28951
rect 13771 28948 13783 28951
rect 13814 28948 13820 28960
rect 13771 28920 13820 28948
rect 13771 28917 13783 28920
rect 13725 28911 13783 28917
rect 13814 28908 13820 28920
rect 13872 28948 13878 28960
rect 14553 28951 14611 28957
rect 14553 28948 14565 28951
rect 13872 28920 14565 28948
rect 13872 28908 13878 28920
rect 14553 28917 14565 28920
rect 14599 28917 14611 28951
rect 14553 28911 14611 28917
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 6825 28747 6883 28753
rect 6825 28713 6837 28747
rect 6871 28744 6883 28747
rect 7558 28744 7564 28756
rect 6871 28716 7564 28744
rect 6871 28713 6883 28716
rect 6825 28707 6883 28713
rect 7558 28704 7564 28716
rect 7616 28704 7622 28756
rect 9309 28747 9367 28753
rect 9309 28713 9321 28747
rect 9355 28744 9367 28747
rect 15746 28744 15752 28756
rect 9355 28716 15752 28744
rect 9355 28713 9367 28716
rect 9309 28707 9367 28713
rect 15746 28704 15752 28716
rect 15804 28704 15810 28756
rect 5166 28636 5172 28688
rect 5224 28676 5230 28688
rect 7282 28676 7288 28688
rect 5224 28648 7288 28676
rect 5224 28636 5230 28648
rect 7282 28636 7288 28648
rect 7340 28636 7346 28688
rect 8386 28636 8392 28688
rect 8444 28676 8450 28688
rect 8444 28648 10640 28676
rect 8444 28636 8450 28648
rect 9122 28608 9128 28620
rect 5920 28580 9128 28608
rect 2038 28500 2044 28552
rect 2096 28500 2102 28552
rect 2308 28543 2366 28549
rect 2308 28509 2320 28543
rect 2354 28540 2366 28543
rect 3418 28540 3424 28552
rect 2354 28512 3424 28540
rect 2354 28509 2366 28512
rect 2308 28503 2366 28509
rect 3418 28500 3424 28512
rect 3476 28500 3482 28552
rect 5920 28549 5948 28580
rect 9122 28568 9128 28580
rect 9180 28568 9186 28620
rect 9490 28568 9496 28620
rect 9548 28608 9554 28620
rect 9548 28580 9996 28608
rect 9548 28568 9554 28580
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 5905 28543 5963 28549
rect 5905 28509 5917 28543
rect 5951 28509 5963 28543
rect 5905 28503 5963 28509
rect 2056 28472 2084 28500
rect 2682 28472 2688 28484
rect 2056 28444 2688 28472
rect 2682 28432 2688 28444
rect 2740 28472 2746 28484
rect 3988 28472 4016 28503
rect 6086 28500 6092 28552
rect 6144 28500 6150 28552
rect 6638 28500 6644 28552
rect 6696 28500 6702 28552
rect 7377 28543 7435 28549
rect 7377 28509 7389 28543
rect 7423 28509 7435 28543
rect 7377 28503 7435 28509
rect 2740 28444 4016 28472
rect 4240 28475 4298 28481
rect 2740 28432 2746 28444
rect 4240 28441 4252 28475
rect 4286 28472 4298 28475
rect 4338 28472 4344 28484
rect 4286 28444 4344 28472
rect 4286 28441 4298 28444
rect 4240 28435 4298 28441
rect 4338 28432 4344 28444
rect 4396 28432 4402 28484
rect 7392 28472 7420 28503
rect 7558 28500 7564 28552
rect 7616 28500 7622 28552
rect 8205 28543 8263 28549
rect 8205 28509 8217 28543
rect 8251 28540 8263 28543
rect 9582 28540 9588 28552
rect 8251 28512 9588 28540
rect 8251 28509 8263 28512
rect 8205 28503 8263 28509
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 9968 28549 9996 28580
rect 10612 28549 10640 28648
rect 14366 28636 14372 28688
rect 14424 28676 14430 28688
rect 14645 28679 14703 28685
rect 14645 28676 14657 28679
rect 14424 28648 14657 28676
rect 14424 28636 14430 28648
rect 14645 28645 14657 28648
rect 14691 28645 14703 28679
rect 14645 28639 14703 28645
rect 11885 28611 11943 28617
rect 11885 28577 11897 28611
rect 11931 28608 11943 28611
rect 12710 28608 12716 28620
rect 11931 28580 12716 28608
rect 11931 28577 11943 28580
rect 11885 28571 11943 28577
rect 12710 28568 12716 28580
rect 12768 28608 12774 28620
rect 13541 28611 13599 28617
rect 13541 28608 13553 28611
rect 12768 28580 13553 28608
rect 12768 28568 12774 28580
rect 9769 28543 9827 28549
rect 9769 28509 9781 28543
rect 9815 28509 9827 28543
rect 9769 28503 9827 28509
rect 9953 28543 10011 28549
rect 9953 28509 9965 28543
rect 9999 28509 10011 28543
rect 9953 28503 10011 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28509 10471 28543
rect 10413 28503 10471 28509
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 11517 28543 11575 28549
rect 11517 28509 11529 28543
rect 11563 28540 11575 28543
rect 12342 28540 12348 28552
rect 11563 28512 12348 28540
rect 11563 28509 11575 28512
rect 11517 28503 11575 28509
rect 7392 28444 7696 28472
rect 3421 28407 3479 28413
rect 3421 28373 3433 28407
rect 3467 28404 3479 28407
rect 3510 28404 3516 28416
rect 3467 28376 3516 28404
rect 3467 28373 3479 28376
rect 3421 28367 3479 28373
rect 3510 28364 3516 28376
rect 3568 28364 3574 28416
rect 5166 28364 5172 28416
rect 5224 28404 5230 28416
rect 5353 28407 5411 28413
rect 5353 28404 5365 28407
rect 5224 28376 5365 28404
rect 5224 28364 5230 28376
rect 5353 28373 5365 28376
rect 5399 28373 5411 28407
rect 5353 28367 5411 28373
rect 5442 28364 5448 28416
rect 5500 28404 5506 28416
rect 5905 28407 5963 28413
rect 5905 28404 5917 28407
rect 5500 28376 5917 28404
rect 5500 28364 5506 28376
rect 5905 28373 5917 28376
rect 5951 28373 5963 28407
rect 5905 28367 5963 28373
rect 7466 28364 7472 28416
rect 7524 28364 7530 28416
rect 7668 28404 7696 28444
rect 7742 28432 7748 28484
rect 7800 28472 7806 28484
rect 9784 28472 9812 28503
rect 10428 28472 10456 28503
rect 12342 28500 12348 28512
rect 12400 28540 12406 28552
rect 13173 28543 13231 28549
rect 12400 28500 12434 28540
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 11698 28472 11704 28484
rect 7800 28444 11704 28472
rect 7800 28432 7806 28444
rect 11698 28432 11704 28444
rect 11756 28432 11762 28484
rect 12406 28472 12434 28500
rect 13188 28472 13216 28503
rect 12406 28444 13216 28472
rect 8021 28407 8079 28413
rect 8021 28404 8033 28407
rect 7668 28376 8033 28404
rect 8021 28373 8033 28376
rect 8067 28404 8079 28407
rect 8570 28404 8576 28416
rect 8067 28376 8576 28404
rect 8067 28373 8079 28376
rect 8021 28367 8079 28373
rect 8570 28364 8576 28376
rect 8628 28364 8634 28416
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 11885 28407 11943 28413
rect 11885 28404 11897 28407
rect 11848 28376 11897 28404
rect 11848 28364 11854 28376
rect 11885 28373 11897 28376
rect 11931 28404 11943 28407
rect 12713 28407 12771 28413
rect 12713 28404 12725 28407
rect 11931 28376 12725 28404
rect 11931 28373 11943 28376
rect 11885 28367 11943 28373
rect 12713 28373 12725 28376
rect 12759 28404 12771 28407
rect 13280 28404 13308 28580
rect 13541 28577 13553 28580
rect 13587 28577 13599 28611
rect 13541 28571 13599 28577
rect 14182 28568 14188 28620
rect 14240 28608 14246 28620
rect 14277 28611 14335 28617
rect 14277 28608 14289 28611
rect 14240 28580 14289 28608
rect 14240 28568 14246 28580
rect 14277 28577 14289 28580
rect 14323 28577 14335 28611
rect 14277 28571 14335 28577
rect 13541 28407 13599 28413
rect 13541 28404 13553 28407
rect 12759 28376 13553 28404
rect 12759 28373 12771 28376
rect 12713 28367 12771 28373
rect 13541 28373 13553 28376
rect 13587 28404 13599 28407
rect 13814 28404 13820 28416
rect 13587 28376 13820 28404
rect 13587 28373 13599 28376
rect 13541 28367 13599 28373
rect 13814 28364 13820 28376
rect 13872 28404 13878 28416
rect 14645 28407 14703 28413
rect 14645 28404 14657 28407
rect 13872 28376 14657 28404
rect 13872 28364 13878 28376
rect 14645 28373 14657 28376
rect 14691 28373 14703 28407
rect 14645 28367 14703 28373
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 4065 28203 4123 28209
rect 4065 28169 4077 28203
rect 4111 28200 4123 28203
rect 4154 28200 4160 28212
rect 4111 28172 4160 28200
rect 4111 28169 4123 28172
rect 4065 28163 4123 28169
rect 4154 28160 4160 28172
rect 4212 28160 4218 28212
rect 4246 28160 4252 28212
rect 4304 28200 4310 28212
rect 4893 28203 4951 28209
rect 4893 28200 4905 28203
rect 4304 28172 4905 28200
rect 4304 28160 4310 28172
rect 4893 28169 4905 28172
rect 4939 28169 4951 28203
rect 4893 28163 4951 28169
rect 8113 28203 8171 28209
rect 8113 28169 8125 28203
rect 8159 28200 8171 28203
rect 8846 28200 8852 28212
rect 8159 28172 8852 28200
rect 8159 28169 8171 28172
rect 8113 28163 8171 28169
rect 8846 28160 8852 28172
rect 8904 28200 8910 28212
rect 8941 28203 8999 28209
rect 8941 28200 8953 28203
rect 8904 28172 8953 28200
rect 8904 28160 8910 28172
rect 8941 28169 8953 28172
rect 8987 28200 8999 28203
rect 10229 28203 10287 28209
rect 10229 28200 10241 28203
rect 8987 28172 10241 28200
rect 8987 28169 8999 28172
rect 8941 28163 8999 28169
rect 10229 28169 10241 28172
rect 10275 28169 10287 28203
rect 10229 28163 10287 28169
rect 3418 28132 3424 28144
rect 2056 28104 3424 28132
rect 1670 28024 1676 28076
rect 1728 28064 1734 28076
rect 1765 28067 1823 28073
rect 1765 28064 1777 28067
rect 1728 28036 1777 28064
rect 1728 28024 1734 28036
rect 1765 28033 1777 28036
rect 1811 28064 1823 28067
rect 1946 28064 1952 28076
rect 1811 28036 1952 28064
rect 1811 28033 1823 28036
rect 1765 28027 1823 28033
rect 1946 28024 1952 28036
rect 2004 28024 2010 28076
rect 2056 28073 2084 28104
rect 3418 28092 3424 28104
rect 3476 28092 3482 28144
rect 5902 28092 5908 28144
rect 5960 28092 5966 28144
rect 6549 28135 6607 28141
rect 6549 28101 6561 28135
rect 6595 28132 6607 28135
rect 6914 28132 6920 28144
rect 6595 28104 6920 28132
rect 6595 28101 6607 28104
rect 6549 28095 6607 28101
rect 6914 28092 6920 28104
rect 6972 28132 6978 28144
rect 6972 28104 10180 28132
rect 6972 28092 6978 28104
rect 2041 28067 2099 28073
rect 2041 28033 2053 28067
rect 2087 28033 2099 28067
rect 2041 28027 2099 28033
rect 2498 28024 2504 28076
rect 2556 28064 2562 28076
rect 2593 28067 2651 28073
rect 2593 28064 2605 28067
rect 2556 28036 2605 28064
rect 2556 28024 2562 28036
rect 2593 28033 2605 28036
rect 2639 28033 2651 28067
rect 2593 28027 2651 28033
rect 3510 28024 3516 28076
rect 3568 28064 3574 28076
rect 4893 28067 4951 28073
rect 4893 28064 4905 28067
rect 3568 28036 4905 28064
rect 3568 28024 3574 28036
rect 4893 28033 4905 28036
rect 4939 28033 4951 28067
rect 4893 28027 4951 28033
rect 2133 27999 2191 28005
rect 2133 27965 2145 27999
rect 2179 27996 2191 27999
rect 4246 27996 4252 28008
rect 2179 27968 4252 27996
rect 2179 27965 2191 27968
rect 2133 27959 2191 27965
rect 4246 27956 4252 27968
rect 4304 27956 4310 28008
rect 4908 27996 4936 28027
rect 4982 28024 4988 28076
rect 5040 28024 5046 28076
rect 5718 28024 5724 28076
rect 5776 28024 5782 28076
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 7466 28024 7472 28076
rect 7524 28064 7530 28076
rect 7745 28067 7803 28073
rect 7745 28064 7757 28067
rect 7524 28036 7757 28064
rect 7524 28024 7530 28036
rect 7745 28033 7757 28036
rect 7791 28064 7803 28067
rect 8573 28067 8631 28073
rect 8573 28064 8585 28067
rect 7791 28036 8585 28064
rect 7791 28033 7803 28036
rect 7745 28027 7803 28033
rect 8573 28033 8585 28036
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 7190 27996 7196 28008
rect 4908 27968 7196 27996
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 8294 27956 8300 28008
rect 8352 27996 8358 28008
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 8352 27968 9873 27996
rect 8352 27956 8358 27968
rect 9861 27965 9873 27968
rect 9907 27965 9919 27999
rect 9861 27959 9919 27965
rect 10042 27956 10048 28008
rect 10100 27996 10106 28008
rect 10152 27996 10180 28104
rect 10244 28073 10272 28163
rect 10229 28067 10287 28073
rect 10229 28033 10241 28067
rect 10275 28033 10287 28067
rect 10229 28027 10287 28033
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 11977 28067 12035 28073
rect 11977 28033 11989 28067
rect 12023 28064 12035 28067
rect 12342 28064 12348 28076
rect 12023 28036 12348 28064
rect 12023 28033 12035 28036
rect 11977 28027 12035 28033
rect 10980 27996 11008 28027
rect 12342 28024 12348 28036
rect 12400 28064 12406 28076
rect 12989 28067 13047 28073
rect 12989 28064 13001 28067
rect 12400 28036 13001 28064
rect 12400 28024 12406 28036
rect 12989 28033 13001 28036
rect 13035 28033 13047 28067
rect 12989 28027 13047 28033
rect 13170 28024 13176 28076
rect 13228 28024 13234 28076
rect 15188 28067 15246 28073
rect 15188 28033 15200 28067
rect 15234 28064 15246 28067
rect 17586 28064 17592 28076
rect 15234 28036 17592 28064
rect 15234 28033 15246 28036
rect 15188 28027 15246 28033
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 10100 27968 11008 27996
rect 10100 27956 10106 27968
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14608 27968 14933 27996
rect 14608 27956 14614 27968
rect 14921 27965 14933 27968
rect 14967 27965 14979 27999
rect 14921 27959 14979 27965
rect 8113 27931 8171 27937
rect 8113 27897 8125 27931
rect 8159 27928 8171 27931
rect 8938 27928 8944 27940
rect 8159 27900 8944 27928
rect 8159 27897 8171 27900
rect 8113 27891 8171 27897
rect 8938 27888 8944 27900
rect 8996 27888 9002 27940
rect 11057 27931 11115 27937
rect 11057 27897 11069 27931
rect 11103 27928 11115 27931
rect 13722 27928 13728 27940
rect 11103 27900 13728 27928
rect 11103 27897 11115 27900
rect 11057 27891 11115 27897
rect 13722 27888 13728 27900
rect 13780 27888 13786 27940
rect 6914 27820 6920 27872
rect 6972 27820 6978 27872
rect 12986 27820 12992 27872
rect 13044 27820 13050 27872
rect 16298 27820 16304 27872
rect 16356 27820 16362 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 2590 27616 2596 27668
rect 2648 27656 2654 27668
rect 2648 27628 2912 27656
rect 2648 27616 2654 27628
rect 2884 27588 2912 27628
rect 4062 27616 4068 27668
rect 4120 27656 4126 27668
rect 6546 27656 6552 27668
rect 4120 27628 6552 27656
rect 4120 27616 4126 27628
rect 6546 27616 6552 27628
rect 6604 27616 6610 27668
rect 8846 27616 8852 27668
rect 8904 27656 8910 27668
rect 10594 27656 10600 27668
rect 8904 27628 10600 27656
rect 8904 27616 8910 27628
rect 10594 27616 10600 27628
rect 10652 27656 10658 27668
rect 11425 27659 11483 27665
rect 11425 27656 11437 27659
rect 10652 27628 11437 27656
rect 10652 27616 10658 27628
rect 11425 27625 11437 27628
rect 11471 27656 11483 27659
rect 11790 27656 11796 27668
rect 11471 27628 11796 27656
rect 11471 27625 11483 27628
rect 11425 27619 11483 27625
rect 5997 27591 6055 27597
rect 5997 27588 6009 27591
rect 2884 27560 6009 27588
rect 5997 27557 6009 27560
rect 6043 27557 6055 27591
rect 5997 27551 6055 27557
rect 6086 27548 6092 27600
rect 6144 27588 6150 27600
rect 6144 27560 7788 27588
rect 6144 27548 6150 27560
rect 7760 27529 7788 27560
rect 9030 27548 9036 27600
rect 9088 27588 9094 27600
rect 9263 27591 9321 27597
rect 9263 27588 9275 27591
rect 9088 27560 9275 27588
rect 9088 27548 9094 27560
rect 9263 27557 9275 27560
rect 9309 27557 9321 27591
rect 9263 27551 9321 27557
rect 7009 27523 7067 27529
rect 7009 27520 7021 27523
rect 3988 27492 7021 27520
rect 1949 27455 2007 27461
rect 1949 27421 1961 27455
rect 1995 27452 2007 27455
rect 2038 27452 2044 27464
rect 1995 27424 2044 27452
rect 1995 27421 2007 27424
rect 1949 27415 2007 27421
rect 2038 27412 2044 27424
rect 2096 27412 2102 27464
rect 2216 27455 2274 27461
rect 2216 27421 2228 27455
rect 2262 27452 2274 27455
rect 3988 27452 4016 27492
rect 7009 27489 7021 27492
rect 7055 27489 7067 27523
rect 7009 27483 7067 27489
rect 7745 27523 7803 27529
rect 7745 27489 7757 27523
rect 7791 27489 7803 27523
rect 7745 27483 7803 27489
rect 8570 27480 8576 27532
rect 8628 27520 8634 27532
rect 11440 27529 11468 27619
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 10229 27523 10287 27529
rect 10229 27520 10241 27523
rect 8628 27492 10241 27520
rect 8628 27480 8634 27492
rect 10229 27489 10241 27492
rect 10275 27520 10287 27523
rect 11057 27523 11115 27529
rect 11057 27520 11069 27523
rect 10275 27492 11069 27520
rect 10275 27489 10287 27492
rect 10229 27483 10287 27489
rect 11057 27489 11069 27492
rect 11103 27489 11115 27523
rect 11057 27483 11115 27489
rect 11425 27523 11483 27529
rect 11425 27489 11437 27523
rect 11471 27489 11483 27523
rect 11425 27483 11483 27489
rect 11974 27480 11980 27532
rect 12032 27480 12038 27532
rect 2262 27424 4016 27452
rect 2262 27421 2274 27424
rect 2216 27415 2274 27421
rect 4062 27412 4068 27464
rect 4120 27412 4126 27464
rect 4172 27424 4844 27452
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 4172 27384 4200 27424
rect 4028 27356 4200 27384
rect 4709 27387 4767 27393
rect 4028 27344 4034 27356
rect 4709 27353 4721 27387
rect 4755 27353 4767 27387
rect 4816 27384 4844 27424
rect 5626 27412 5632 27464
rect 5684 27452 5690 27464
rect 6917 27455 6975 27461
rect 6917 27452 6929 27455
rect 5684 27424 6929 27452
rect 5684 27412 5690 27424
rect 6917 27421 6929 27424
rect 6963 27421 6975 27455
rect 6917 27415 6975 27421
rect 7101 27455 7159 27461
rect 7101 27421 7113 27455
rect 7147 27421 7159 27455
rect 7101 27415 7159 27421
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27421 7527 27455
rect 8205 27455 8263 27461
rect 8205 27452 8217 27455
rect 7469 27415 7527 27421
rect 7760 27424 8217 27452
rect 7116 27384 7144 27415
rect 4816 27356 7144 27384
rect 4709 27347 4767 27353
rect 3329 27319 3387 27325
rect 3329 27285 3341 27319
rect 3375 27316 3387 27319
rect 4154 27316 4160 27328
rect 3375 27288 4160 27316
rect 3375 27285 3387 27288
rect 3329 27279 3387 27285
rect 4154 27276 4160 27288
rect 4212 27276 4218 27328
rect 4249 27319 4307 27325
rect 4249 27285 4261 27319
rect 4295 27316 4307 27319
rect 4724 27316 4752 27347
rect 4295 27288 4752 27316
rect 7484 27316 7512 27415
rect 7760 27396 7788 27424
rect 8205 27421 8217 27424
rect 8251 27421 8263 27455
rect 8205 27415 8263 27421
rect 8386 27412 8392 27464
rect 8444 27412 8450 27464
rect 8478 27412 8484 27464
rect 8536 27452 8542 27464
rect 9160 27455 9218 27461
rect 9160 27452 9172 27455
rect 8536 27424 9172 27452
rect 8536 27412 8542 27424
rect 9160 27421 9172 27424
rect 9206 27421 9218 27455
rect 9160 27415 9218 27421
rect 10594 27412 10600 27464
rect 10652 27412 10658 27464
rect 11882 27412 11888 27464
rect 11940 27412 11946 27464
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 13170 27452 13176 27464
rect 12115 27424 13176 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 7742 27344 7748 27396
rect 7800 27344 7806 27396
rect 9398 27344 9404 27396
rect 9456 27384 9462 27396
rect 12084 27384 12112 27415
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27452 18107 27455
rect 18322 27452 18328 27464
rect 18095 27424 18328 27452
rect 18095 27421 18107 27424
rect 18049 27415 18107 27421
rect 18322 27412 18328 27424
rect 18380 27412 18386 27464
rect 18417 27455 18475 27461
rect 18417 27421 18429 27455
rect 18463 27421 18475 27455
rect 18417 27415 18475 27421
rect 9456 27356 12112 27384
rect 9456 27344 9462 27356
rect 10134 27316 10140 27328
rect 7484 27288 10140 27316
rect 4295 27285 4307 27288
rect 4249 27279 4307 27285
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 14277 27319 14335 27325
rect 14277 27285 14289 27319
rect 14323 27316 14335 27319
rect 14366 27316 14372 27328
rect 14323 27288 14372 27316
rect 14323 27285 14335 27288
rect 14277 27279 14335 27285
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 14458 27276 14464 27328
rect 14516 27316 14522 27328
rect 18432 27325 18460 27415
rect 20714 27412 20720 27464
rect 20772 27412 20778 27464
rect 20254 27344 20260 27396
rect 20312 27384 20318 27396
rect 20962 27387 21020 27393
rect 20962 27384 20974 27387
rect 20312 27356 20974 27384
rect 20312 27344 20318 27356
rect 20962 27353 20974 27356
rect 21008 27353 21020 27387
rect 20962 27347 21020 27353
rect 18417 27319 18475 27325
rect 18417 27316 18429 27319
rect 14516 27288 18429 27316
rect 14516 27276 14522 27288
rect 18417 27285 18429 27288
rect 18463 27285 18475 27319
rect 18417 27279 18475 27285
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22554 27316 22560 27328
rect 22143 27288 22560 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22554 27276 22560 27288
rect 22612 27276 22618 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 1854 27072 1860 27124
rect 1912 27112 1918 27124
rect 1949 27115 2007 27121
rect 1949 27112 1961 27115
rect 1912 27084 1961 27112
rect 1912 27072 1918 27084
rect 1949 27081 1961 27084
rect 1995 27081 2007 27115
rect 1949 27075 2007 27081
rect 2225 27115 2283 27121
rect 2225 27081 2237 27115
rect 2271 27112 2283 27115
rect 4062 27112 4068 27124
rect 2271 27084 4068 27112
rect 2271 27081 2283 27084
rect 2225 27075 2283 27081
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 7466 27112 7472 27124
rect 4212 27084 7472 27112
rect 4212 27072 4218 27084
rect 7466 27072 7472 27084
rect 7524 27072 7530 27124
rect 7558 27072 7564 27124
rect 7616 27112 7622 27124
rect 9398 27112 9404 27124
rect 7616 27084 9404 27112
rect 7616 27072 7622 27084
rect 9398 27072 9404 27084
rect 9456 27072 9462 27124
rect 11698 27072 11704 27124
rect 11756 27072 11762 27124
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 13814 27112 13820 27124
rect 13596 27084 13820 27112
rect 13596 27072 13602 27084
rect 13814 27072 13820 27084
rect 13872 27112 13878 27124
rect 14369 27115 14427 27121
rect 14369 27112 14381 27115
rect 13872 27084 14381 27112
rect 13872 27072 13878 27084
rect 14369 27081 14381 27084
rect 14415 27112 14427 27115
rect 14458 27112 14464 27124
rect 14415 27084 14464 27112
rect 14415 27081 14427 27084
rect 14369 27075 14427 27081
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 5442 27044 5448 27056
rect 5000 27016 5448 27044
rect 2682 26936 2688 26988
rect 2740 26976 2746 26988
rect 5000 26985 5028 27016
rect 5442 27004 5448 27016
rect 5500 27004 5506 27056
rect 7098 27004 7104 27056
rect 7156 27044 7162 27056
rect 7576 27044 7604 27072
rect 7156 27016 7604 27044
rect 7156 27004 7162 27016
rect 2777 26979 2835 26985
rect 2777 26976 2789 26979
rect 2740 26948 2789 26976
rect 2740 26936 2746 26948
rect 2777 26945 2789 26948
rect 2823 26945 2835 26979
rect 2777 26939 2835 26945
rect 3044 26979 3102 26985
rect 3044 26945 3056 26979
rect 3090 26976 3102 26979
rect 4801 26979 4859 26985
rect 4801 26976 4813 26979
rect 3090 26948 4813 26976
rect 3090 26945 3102 26948
rect 3044 26939 3102 26945
rect 4801 26945 4813 26948
rect 4847 26945 4859 26979
rect 4801 26939 4859 26945
rect 4985 26979 5043 26985
rect 4985 26945 4997 26979
rect 5031 26945 5043 26979
rect 4985 26939 5043 26945
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26945 5319 26979
rect 5261 26939 5319 26945
rect 5537 26979 5595 26985
rect 5537 26945 5549 26979
rect 5583 26976 5595 26979
rect 6086 26976 6092 26988
rect 5583 26948 6092 26976
rect 5583 26945 5595 26948
rect 5537 26939 5595 26945
rect 1581 26911 1639 26917
rect 1581 26877 1593 26911
rect 1627 26877 1639 26911
rect 1581 26871 1639 26877
rect 1596 26772 1624 26871
rect 1854 26868 1860 26920
rect 1912 26868 1918 26920
rect 2041 26911 2099 26917
rect 2041 26877 2053 26911
rect 2087 26908 2099 26911
rect 2406 26908 2412 26920
rect 2087 26880 2412 26908
rect 2087 26877 2099 26880
rect 2041 26871 2099 26877
rect 2406 26868 2412 26880
rect 2464 26868 2470 26920
rect 4706 26868 4712 26920
rect 4764 26868 4770 26920
rect 5166 26840 5172 26852
rect 4080 26812 5172 26840
rect 4080 26772 4108 26812
rect 5166 26800 5172 26812
rect 5224 26800 5230 26852
rect 5276 26840 5304 26939
rect 6086 26936 6092 26948
rect 6144 26936 6150 26988
rect 6362 26936 6368 26988
rect 6420 26976 6426 26988
rect 7576 26985 7604 27016
rect 7650 27004 7656 27056
rect 7708 27044 7714 27056
rect 20714 27044 20720 27056
rect 7708 27016 8248 27044
rect 7708 27004 7714 27016
rect 6549 26979 6607 26985
rect 6549 26976 6561 26979
rect 6420 26948 6561 26976
rect 6420 26936 6426 26948
rect 6549 26945 6561 26948
rect 6595 26945 6607 26979
rect 6549 26939 6607 26945
rect 6733 26979 6791 26985
rect 6733 26945 6745 26979
rect 6779 26945 6791 26979
rect 6733 26939 6791 26945
rect 7377 26979 7435 26985
rect 7377 26945 7389 26979
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 7561 26979 7619 26985
rect 7561 26945 7573 26979
rect 7607 26945 7619 26979
rect 7561 26939 7619 26945
rect 6454 26868 6460 26920
rect 6512 26908 6518 26920
rect 6748 26908 6776 26939
rect 6512 26880 6776 26908
rect 7392 26908 7420 26939
rect 7742 26936 7748 26988
rect 7800 26976 7806 26988
rect 8220 26985 8248 27016
rect 19168 27016 20720 27044
rect 19168 26988 19196 27016
rect 20714 27004 20720 27016
rect 20772 27004 20778 27056
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 7800 26948 8033 26976
rect 7800 26936 7806 26948
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 8205 26979 8263 26985
rect 8205 26945 8217 26979
rect 8251 26945 8263 26979
rect 8205 26939 8263 26945
rect 12066 26936 12072 26988
rect 12124 26936 12130 26988
rect 12986 26936 12992 26988
rect 13044 26976 13050 26988
rect 13173 26979 13231 26985
rect 13173 26976 13185 26979
rect 13044 26948 13185 26976
rect 13044 26936 13050 26948
rect 13173 26945 13185 26948
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13722 26936 13728 26988
rect 13780 26976 13786 26988
rect 14001 26979 14059 26985
rect 14001 26976 14013 26979
rect 13780 26948 14013 26976
rect 13780 26936 13786 26948
rect 14001 26945 14013 26948
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14366 26936 14372 26988
rect 14424 26936 14430 26988
rect 18322 26936 18328 26988
rect 18380 26936 18386 26988
rect 19150 26936 19156 26988
rect 19208 26936 19214 26988
rect 19420 26979 19478 26985
rect 19420 26945 19432 26979
rect 19466 26976 19478 26979
rect 20622 26976 20628 26988
rect 19466 26948 20628 26976
rect 19466 26945 19478 26948
rect 19420 26939 19478 26945
rect 20622 26936 20628 26948
rect 20680 26936 20686 26988
rect 22830 26936 22836 26988
rect 22888 26976 22894 26988
rect 23273 26979 23331 26985
rect 23273 26976 23285 26979
rect 22888 26948 23285 26976
rect 22888 26936 22894 26948
rect 23273 26945 23285 26948
rect 23319 26945 23331 26979
rect 23273 26939 23331 26945
rect 8294 26908 8300 26920
rect 7392 26880 8300 26908
rect 6512 26868 6518 26880
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 10042 26868 10048 26920
rect 10100 26908 10106 26920
rect 12161 26911 12219 26917
rect 12161 26908 12173 26911
rect 10100 26880 12173 26908
rect 10100 26868 10106 26880
rect 12161 26877 12173 26880
rect 12207 26877 12219 26911
rect 12161 26871 12219 26877
rect 12345 26911 12403 26917
rect 12345 26877 12357 26911
rect 12391 26908 12403 26911
rect 12710 26908 12716 26920
rect 12391 26880 12716 26908
rect 12391 26877 12403 26880
rect 12345 26871 12403 26877
rect 12710 26868 12716 26880
rect 12768 26908 12774 26920
rect 13541 26911 13599 26917
rect 13541 26908 13553 26911
rect 12768 26880 13553 26908
rect 12768 26868 12774 26880
rect 13541 26877 13553 26880
rect 13587 26877 13599 26911
rect 13541 26871 13599 26877
rect 21818 26868 21824 26920
rect 21876 26908 21882 26920
rect 23017 26911 23075 26917
rect 23017 26908 23029 26911
rect 21876 26880 23029 26908
rect 21876 26868 21882 26880
rect 23017 26877 23029 26880
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 9858 26840 9864 26852
rect 5276 26812 9864 26840
rect 9858 26800 9864 26812
rect 9916 26800 9922 26852
rect 1596 26744 4108 26772
rect 4154 26732 4160 26784
rect 4212 26732 4218 26784
rect 4706 26732 4712 26784
rect 4764 26772 4770 26784
rect 5626 26772 5632 26784
rect 4764 26744 5632 26772
rect 4764 26732 4770 26744
rect 5626 26732 5632 26744
rect 5684 26732 5690 26784
rect 5718 26732 5724 26784
rect 5776 26772 5782 26784
rect 6641 26775 6699 26781
rect 6641 26772 6653 26775
rect 5776 26744 6653 26772
rect 5776 26732 5782 26744
rect 6641 26741 6653 26744
rect 6687 26741 6699 26775
rect 6641 26735 6699 26741
rect 7377 26775 7435 26781
rect 7377 26741 7389 26775
rect 7423 26772 7435 26775
rect 8202 26772 8208 26784
rect 7423 26744 8208 26772
rect 7423 26741 7435 26744
rect 7377 26735 7435 26741
rect 8202 26732 8208 26744
rect 8260 26732 8266 26784
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 20533 26775 20591 26781
rect 20533 26772 20545 26775
rect 20312 26744 20545 26772
rect 20312 26732 20318 26744
rect 20533 26741 20545 26744
rect 20579 26741 20591 26775
rect 20533 26735 20591 26741
rect 24394 26732 24400 26784
rect 24452 26732 24458 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 7377 26571 7435 26577
rect 2464 26540 7328 26568
rect 2464 26528 2470 26540
rect 5350 26460 5356 26512
rect 5408 26460 5414 26512
rect 7098 26500 7104 26512
rect 5460 26472 7104 26500
rect 2038 26392 2044 26444
rect 2096 26432 2102 26444
rect 2682 26432 2688 26444
rect 2096 26404 2688 26432
rect 2096 26392 2102 26404
rect 2682 26392 2688 26404
rect 2740 26432 2746 26444
rect 3973 26435 4031 26441
rect 3973 26432 3985 26435
rect 2740 26404 3985 26432
rect 2740 26392 2746 26404
rect 3973 26401 3985 26404
rect 4019 26401 4031 26435
rect 3973 26395 4031 26401
rect 1578 26324 1584 26376
rect 1636 26324 1642 26376
rect 4246 26373 4252 26376
rect 4240 26327 4252 26373
rect 4246 26324 4252 26327
rect 4304 26324 4310 26376
rect 5460 26364 5488 26472
rect 7098 26460 7104 26472
rect 7156 26460 7162 26512
rect 7300 26500 7328 26540
rect 7377 26537 7389 26571
rect 7423 26568 7435 26571
rect 8294 26568 8300 26580
rect 7423 26540 8300 26568
rect 7423 26537 7435 26540
rect 7377 26531 7435 26537
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8846 26568 8852 26580
rect 8619 26540 8852 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8846 26528 8852 26540
rect 8904 26528 8910 26580
rect 9582 26528 9588 26580
rect 9640 26528 9646 26580
rect 12713 26571 12771 26577
rect 12713 26537 12725 26571
rect 12759 26568 12771 26571
rect 13538 26568 13544 26580
rect 12759 26540 13544 26568
rect 12759 26537 12771 26540
rect 12713 26531 12771 26537
rect 13538 26528 13544 26540
rect 13596 26528 13602 26580
rect 17586 26528 17592 26580
rect 17644 26528 17650 26580
rect 22830 26528 22836 26580
rect 22888 26568 22894 26580
rect 26973 26571 27031 26577
rect 26973 26568 26985 26571
rect 22888 26540 26985 26568
rect 22888 26528 22894 26540
rect 26973 26537 26985 26540
rect 27019 26537 27031 26571
rect 26973 26531 27031 26537
rect 9950 26500 9956 26512
rect 7300 26472 9956 26500
rect 9950 26460 9956 26472
rect 10008 26460 10014 26512
rect 5534 26392 5540 26444
rect 5592 26432 5598 26444
rect 6917 26435 6975 26441
rect 6917 26432 6929 26435
rect 5592 26404 6929 26432
rect 5592 26392 5598 26404
rect 6917 26401 6929 26404
rect 6963 26401 6975 26435
rect 6917 26395 6975 26401
rect 8202 26392 8208 26444
rect 8260 26392 8266 26444
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26401 10195 26435
rect 10137 26395 10195 26401
rect 12345 26435 12403 26441
rect 12345 26401 12357 26435
rect 12391 26432 12403 26435
rect 12986 26432 12992 26444
rect 12391 26404 12992 26432
rect 12391 26401 12403 26404
rect 12345 26395 12403 26401
rect 5813 26367 5871 26373
rect 5813 26364 5825 26367
rect 5460 26336 5825 26364
rect 5813 26333 5825 26336
rect 5859 26333 5871 26367
rect 5813 26327 5871 26333
rect 5994 26324 6000 26376
rect 6052 26324 6058 26376
rect 6549 26367 6607 26373
rect 6549 26333 6561 26367
rect 6595 26364 6607 26367
rect 7561 26367 7619 26373
rect 6595 26336 7512 26364
rect 6595 26333 6607 26336
rect 6549 26327 6607 26333
rect 4798 26256 4804 26308
rect 4856 26296 4862 26308
rect 5905 26299 5963 26305
rect 5905 26296 5917 26299
rect 4856 26268 5917 26296
rect 4856 26256 4862 26268
rect 5905 26265 5917 26268
rect 5951 26265 5963 26299
rect 5905 26259 5963 26265
rect 6730 26256 6736 26308
rect 6788 26256 6794 26308
rect 7484 26296 7512 26336
rect 7561 26333 7573 26367
rect 7607 26364 7619 26367
rect 8478 26364 8484 26376
rect 7607 26336 8484 26364
rect 7607 26333 7619 26336
rect 7561 26327 7619 26333
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 8570 26324 8576 26376
rect 8628 26324 8634 26376
rect 9674 26324 9680 26376
rect 9732 26364 9738 26376
rect 9953 26367 10011 26373
rect 9953 26364 9965 26367
rect 9732 26336 9965 26364
rect 9732 26324 9738 26336
rect 9953 26333 9965 26336
rect 9999 26364 10011 26367
rect 10042 26364 10048 26376
rect 9999 26336 10048 26364
rect 9999 26333 10011 26336
rect 9953 26327 10011 26333
rect 10042 26324 10048 26336
rect 10100 26324 10106 26376
rect 8846 26296 8852 26308
rect 7484 26268 8852 26296
rect 8846 26256 8852 26268
rect 8904 26296 8910 26308
rect 10152 26296 10180 26395
rect 12986 26392 12992 26404
rect 13044 26432 13050 26444
rect 13173 26435 13231 26441
rect 13173 26432 13185 26435
rect 13044 26404 13185 26432
rect 13044 26392 13050 26404
rect 13173 26401 13185 26404
rect 13219 26401 13231 26435
rect 13173 26395 13231 26401
rect 21450 26392 21456 26444
rect 21508 26432 21514 26444
rect 21818 26432 21824 26444
rect 21508 26404 21824 26432
rect 21508 26392 21514 26404
rect 21818 26392 21824 26404
rect 21876 26392 21882 26444
rect 12710 26324 12716 26376
rect 12768 26364 12774 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 12768 26336 13553 26364
rect 12768 26324 12774 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26364 16267 26367
rect 18322 26364 18328 26376
rect 16255 26336 18328 26364
rect 16255 26333 16267 26336
rect 16209 26327 16267 26333
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 25593 26367 25651 26373
rect 25593 26364 25605 26367
rect 25188 26336 25605 26364
rect 25188 26324 25194 26336
rect 25593 26333 25605 26336
rect 25639 26333 25651 26367
rect 25593 26327 25651 26333
rect 10226 26296 10232 26308
rect 8904 26268 10232 26296
rect 8904 26256 8910 26268
rect 10226 26256 10232 26268
rect 10284 26256 10290 26308
rect 16476 26299 16534 26305
rect 12636 26268 12848 26296
rect 2682 26188 2688 26240
rect 2740 26228 2746 26240
rect 2869 26231 2927 26237
rect 2869 26228 2881 26231
rect 2740 26200 2881 26228
rect 2740 26188 2746 26200
rect 2869 26197 2881 26200
rect 2915 26197 2927 26231
rect 2869 26191 2927 26197
rect 5350 26188 5356 26240
rect 5408 26228 5414 26240
rect 9766 26228 9772 26240
rect 5408 26200 9772 26228
rect 5408 26188 5414 26200
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 12066 26228 12072 26240
rect 10100 26200 12072 26228
rect 10100 26188 10106 26200
rect 12066 26188 12072 26200
rect 12124 26188 12130 26240
rect 12158 26188 12164 26240
rect 12216 26228 12222 26240
rect 12636 26228 12664 26268
rect 12216 26200 12664 26228
rect 12820 26228 12848 26268
rect 16476 26265 16488 26299
rect 16522 26296 16534 26299
rect 17402 26296 17408 26308
rect 16522 26268 17408 26296
rect 16522 26265 16534 26268
rect 16476 26259 16534 26265
rect 17402 26256 17408 26268
rect 17460 26256 17466 26308
rect 22088 26299 22146 26305
rect 22088 26265 22100 26299
rect 22134 26296 22146 26299
rect 22554 26296 22560 26308
rect 22134 26268 22560 26296
rect 22134 26265 22146 26268
rect 22088 26259 22146 26265
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 25038 26256 25044 26308
rect 25096 26296 25102 26308
rect 25838 26299 25896 26305
rect 25838 26296 25850 26299
rect 25096 26268 25850 26296
rect 25096 26256 25102 26268
rect 25838 26265 25850 26268
rect 25884 26296 25896 26299
rect 26142 26296 26148 26308
rect 25884 26268 26148 26296
rect 25884 26265 25896 26268
rect 25838 26259 25896 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 17678 26234 17684 26240
rect 13464 26228 13676 26234
rect 17512 26228 17684 26234
rect 12820 26206 17684 26228
rect 12820 26200 13492 26206
rect 13648 26200 17540 26206
rect 12216 26188 12222 26200
rect 17678 26188 17684 26206
rect 17736 26188 17742 26240
rect 18322 26188 18328 26240
rect 18380 26228 18386 26240
rect 19150 26228 19156 26240
rect 18380 26200 19156 26228
rect 18380 26188 18386 26200
rect 19150 26188 19156 26200
rect 19208 26188 19214 26240
rect 23198 26188 23204 26240
rect 23256 26188 23262 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 4415 26027 4473 26033
rect 4415 26024 4427 26027
rect 1964 25996 4427 26024
rect 1964 25956 1992 25996
rect 4415 25993 4427 25996
rect 4461 25993 4473 26027
rect 4415 25987 4473 25993
rect 4893 26027 4951 26033
rect 4893 25993 4905 26027
rect 4939 26024 4951 26027
rect 5350 26024 5356 26036
rect 4939 25996 5356 26024
rect 4939 25993 4951 25996
rect 4893 25987 4951 25993
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 5442 25984 5448 26036
rect 5500 26024 5506 26036
rect 5500 25996 6684 26024
rect 5500 25984 5506 25996
rect 1872 25928 1992 25956
rect 5000 25928 5764 25956
rect 1670 25848 1676 25900
rect 1728 25888 1734 25900
rect 1872 25897 1900 25928
rect 1857 25891 1915 25897
rect 1728 25860 1808 25888
rect 1728 25848 1734 25860
rect 1780 25684 1808 25860
rect 1857 25857 1869 25891
rect 1903 25857 1915 25891
rect 1857 25851 1915 25857
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25888 2007 25891
rect 2665 25891 2723 25897
rect 2665 25888 2677 25891
rect 1995 25860 2677 25888
rect 1995 25857 2007 25860
rect 1949 25851 2007 25857
rect 2665 25857 2677 25860
rect 2711 25857 2723 25891
rect 2665 25851 2723 25857
rect 4062 25848 4068 25900
rect 4120 25888 4126 25900
rect 5000 25888 5028 25928
rect 4120 25860 5028 25888
rect 4120 25848 4126 25860
rect 5626 25848 5632 25900
rect 5684 25848 5690 25900
rect 5736 25897 5764 25928
rect 6546 25916 6552 25968
rect 6604 25916 6610 25968
rect 6656 25956 6684 25996
rect 6822 25984 6828 26036
rect 6880 25984 6886 26036
rect 6917 26027 6975 26033
rect 6917 25993 6929 26027
rect 6963 25993 6975 26027
rect 6917 25987 6975 25993
rect 6932 25956 6960 25987
rect 8938 25984 8944 26036
rect 8996 25984 9002 26036
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 11790 26024 11796 26036
rect 9824 25996 11796 26024
rect 9824 25984 9830 25996
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 13538 25984 13544 26036
rect 13596 25984 13602 26036
rect 26142 25984 26148 26036
rect 26200 26024 26206 26036
rect 26605 26027 26663 26033
rect 26605 26024 26617 26027
rect 26200 25996 26617 26024
rect 26200 25984 26206 25996
rect 26605 25993 26617 25996
rect 26651 25993 26663 26027
rect 26605 25987 26663 25993
rect 6656 25928 6960 25956
rect 7190 25916 7196 25968
rect 7248 25956 7254 25968
rect 9214 25956 9220 25968
rect 7248 25928 9220 25956
rect 7248 25916 7254 25928
rect 9214 25916 9220 25928
rect 9272 25916 9278 25968
rect 10873 25959 10931 25965
rect 10873 25925 10885 25959
rect 10919 25956 10931 25959
rect 12342 25956 12348 25968
rect 10919 25928 12348 25956
rect 10919 25925 10931 25928
rect 10873 25919 10931 25925
rect 12342 25916 12348 25928
rect 12400 25916 12406 25968
rect 13262 25956 13268 25968
rect 12728 25928 13268 25956
rect 12728 25900 12756 25928
rect 13262 25916 13268 25928
rect 13320 25916 13326 25968
rect 16209 25959 16267 25965
rect 16209 25925 16221 25959
rect 16255 25956 16267 25959
rect 16574 25956 16580 25968
rect 16255 25928 16580 25956
rect 16255 25925 16267 25928
rect 16209 25919 16267 25925
rect 16574 25916 16580 25928
rect 16632 25916 16638 25968
rect 18592 25959 18650 25965
rect 18592 25925 18604 25959
rect 18638 25956 18650 25959
rect 19242 25956 19248 25968
rect 18638 25928 19248 25956
rect 18638 25925 18650 25928
rect 18592 25919 18650 25925
rect 19242 25916 19248 25928
rect 19300 25916 19306 25968
rect 25492 25959 25550 25965
rect 25492 25925 25504 25959
rect 25538 25956 25550 25959
rect 25590 25956 25596 25968
rect 25538 25928 25596 25956
rect 25538 25925 25550 25928
rect 25492 25919 25550 25925
rect 25590 25916 25596 25928
rect 25648 25916 25654 25968
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25888 6791 25891
rect 6914 25888 6920 25900
rect 6779 25860 6920 25888
rect 6779 25857 6791 25860
rect 6733 25851 6791 25857
rect 6914 25848 6920 25860
rect 6972 25848 6978 25900
rect 7098 25848 7104 25900
rect 7156 25848 7162 25900
rect 8846 25848 8852 25900
rect 8904 25848 8910 25900
rect 10410 25848 10416 25900
rect 10468 25888 10474 25900
rect 10689 25891 10747 25897
rect 10689 25888 10701 25891
rect 10468 25860 10701 25888
rect 10468 25848 10474 25860
rect 10689 25857 10701 25860
rect 10735 25857 10747 25891
rect 10689 25851 10747 25857
rect 10962 25848 10968 25900
rect 11020 25848 11026 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 12710 25888 12716 25900
rect 12299 25860 12716 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 12710 25848 12716 25860
rect 12768 25848 12774 25900
rect 12986 25848 12992 25900
rect 13044 25888 13050 25900
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 13044 25860 13185 25888
rect 13044 25848 13050 25860
rect 13173 25857 13185 25860
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 16022 25848 16028 25900
rect 16080 25848 16086 25900
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 17218 25888 17224 25900
rect 16347 25860 17224 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 17218 25848 17224 25860
rect 17276 25848 17282 25900
rect 18322 25848 18328 25900
rect 18380 25848 18386 25900
rect 2038 25780 2044 25832
rect 2096 25820 2102 25832
rect 2409 25823 2467 25829
rect 2409 25820 2421 25823
rect 2096 25792 2421 25820
rect 2096 25780 2102 25792
rect 2409 25789 2421 25792
rect 2455 25789 2467 25823
rect 2409 25783 2467 25789
rect 4798 25780 4804 25832
rect 4856 25780 4862 25832
rect 4982 25780 4988 25832
rect 5040 25780 5046 25832
rect 5166 25780 5172 25832
rect 5224 25820 5230 25832
rect 10505 25823 10563 25829
rect 10505 25820 10517 25823
rect 5224 25792 10517 25820
rect 5224 25780 5230 25792
rect 10505 25789 10517 25792
rect 10551 25789 10563 25823
rect 10505 25783 10563 25789
rect 25130 25780 25136 25832
rect 25188 25820 25194 25832
rect 25225 25823 25283 25829
rect 25225 25820 25237 25823
rect 25188 25792 25237 25820
rect 25188 25780 25194 25792
rect 25225 25789 25237 25792
rect 25271 25789 25283 25823
rect 25225 25783 25283 25789
rect 3712 25724 4108 25752
rect 3712 25684 3740 25724
rect 1780 25656 3740 25684
rect 3789 25687 3847 25693
rect 3789 25653 3801 25687
rect 3835 25684 3847 25687
rect 3970 25684 3976 25696
rect 3835 25656 3976 25684
rect 3835 25653 3847 25656
rect 3789 25647 3847 25653
rect 3970 25644 3976 25656
rect 4028 25644 4034 25696
rect 4080 25684 4108 25724
rect 4246 25712 4252 25764
rect 4304 25752 4310 25764
rect 5813 25755 5871 25761
rect 5813 25752 5825 25755
rect 4304 25724 5825 25752
rect 4304 25712 4310 25724
rect 5813 25721 5825 25724
rect 5859 25721 5871 25755
rect 5813 25715 5871 25721
rect 12618 25712 12624 25764
rect 12676 25752 12682 25764
rect 13541 25755 13599 25761
rect 13541 25752 13553 25755
rect 12676 25724 13553 25752
rect 12676 25712 12682 25724
rect 13541 25721 13553 25724
rect 13587 25721 13599 25755
rect 13541 25715 13599 25721
rect 5626 25684 5632 25696
rect 4080 25656 5632 25684
rect 5626 25644 5632 25656
rect 5684 25684 5690 25696
rect 5994 25684 6000 25696
rect 5684 25656 6000 25684
rect 5684 25644 5690 25656
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 12345 25687 12403 25693
rect 12345 25684 12357 25687
rect 12308 25656 12357 25684
rect 12308 25644 12314 25656
rect 12345 25653 12357 25656
rect 12391 25653 12403 25687
rect 12345 25647 12403 25653
rect 15838 25644 15844 25696
rect 15896 25644 15902 25696
rect 19702 25644 19708 25696
rect 19760 25644 19766 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 1946 25440 1952 25492
rect 2004 25480 2010 25492
rect 2004 25452 3372 25480
rect 2004 25440 2010 25452
rect 3344 25412 3372 25452
rect 3418 25440 3424 25492
rect 3476 25480 3482 25492
rect 4065 25483 4123 25489
rect 4065 25480 4077 25483
rect 3476 25452 4077 25480
rect 3476 25440 3482 25452
rect 4065 25449 4077 25452
rect 4111 25449 4123 25483
rect 4065 25443 4123 25449
rect 5810 25440 5816 25492
rect 5868 25480 5874 25492
rect 6089 25483 6147 25489
rect 6089 25480 6101 25483
rect 5868 25452 6101 25480
rect 5868 25440 5874 25452
rect 6089 25449 6101 25452
rect 6135 25449 6147 25483
rect 6089 25443 6147 25449
rect 6273 25483 6331 25489
rect 6273 25449 6285 25483
rect 6319 25480 6331 25483
rect 7098 25480 7104 25492
rect 6319 25452 7104 25480
rect 6319 25449 6331 25452
rect 6273 25443 6331 25449
rect 3344 25384 5856 25412
rect 5828 25356 5856 25384
rect 4617 25347 4675 25353
rect 4617 25313 4629 25347
rect 4663 25344 4675 25347
rect 4982 25344 4988 25356
rect 4663 25316 4988 25344
rect 4663 25313 4675 25316
rect 4617 25307 4675 25313
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 5166 25304 5172 25356
rect 5224 25344 5230 25356
rect 5721 25347 5779 25353
rect 5721 25344 5733 25347
rect 5224 25316 5733 25344
rect 5224 25304 5230 25316
rect 5721 25313 5733 25316
rect 5767 25313 5779 25347
rect 5721 25307 5779 25313
rect 2038 25236 2044 25288
rect 2096 25236 2102 25288
rect 2308 25279 2366 25285
rect 2308 25245 2320 25279
rect 2354 25276 2366 25279
rect 4246 25276 4252 25288
rect 2354 25248 4252 25276
rect 2354 25245 2366 25248
rect 2308 25239 2366 25245
rect 4246 25236 4252 25248
rect 4304 25236 4310 25288
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25276 4399 25279
rect 5350 25276 5356 25288
rect 4387 25248 5356 25276
rect 4387 25245 4399 25248
rect 4341 25239 4399 25245
rect 5350 25236 5356 25248
rect 5408 25236 5414 25288
rect 5736 25276 5764 25307
rect 5810 25304 5816 25356
rect 5868 25304 5874 25356
rect 6104 25344 6132 25443
rect 7098 25440 7104 25452
rect 7156 25440 7162 25492
rect 7374 25440 7380 25492
rect 7432 25480 7438 25492
rect 7561 25483 7619 25489
rect 7561 25480 7573 25483
rect 7432 25452 7573 25480
rect 7432 25440 7438 25452
rect 7561 25449 7573 25452
rect 7607 25449 7619 25483
rect 7561 25443 7619 25449
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 8570 25480 8576 25492
rect 8435 25452 8576 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 8570 25440 8576 25452
rect 8628 25440 8634 25492
rect 11609 25483 11667 25489
rect 11609 25449 11621 25483
rect 11655 25480 11667 25483
rect 11882 25480 11888 25492
rect 11655 25452 11888 25480
rect 11655 25449 11667 25452
rect 11609 25443 11667 25449
rect 11882 25440 11888 25452
rect 11940 25440 11946 25492
rect 17678 25440 17684 25492
rect 17736 25480 17742 25492
rect 25317 25483 25375 25489
rect 25317 25480 25329 25483
rect 17736 25452 25329 25480
rect 17736 25440 17742 25452
rect 25317 25449 25329 25452
rect 25363 25449 25375 25483
rect 25317 25443 25375 25449
rect 7006 25372 7012 25424
rect 7064 25412 7070 25424
rect 7745 25415 7803 25421
rect 7745 25412 7757 25415
rect 7064 25384 7757 25412
rect 7064 25372 7070 25384
rect 7745 25381 7757 25384
rect 7791 25412 7803 25415
rect 8202 25412 8208 25424
rect 7791 25384 8208 25412
rect 7791 25381 7803 25384
rect 7745 25375 7803 25381
rect 8202 25372 8208 25384
rect 8260 25372 8266 25424
rect 8478 25372 8484 25424
rect 8536 25412 8542 25424
rect 9125 25415 9183 25421
rect 9125 25412 9137 25415
rect 8536 25384 9137 25412
rect 8536 25372 8542 25384
rect 9125 25381 9137 25384
rect 9171 25381 9183 25415
rect 9125 25375 9183 25381
rect 10410 25372 10416 25424
rect 10468 25412 10474 25424
rect 10468 25384 13032 25412
rect 10468 25372 10474 25384
rect 7650 25344 7656 25356
rect 6104 25316 7656 25344
rect 7650 25304 7656 25316
rect 7708 25344 7714 25356
rect 8570 25344 8576 25356
rect 7708 25316 8576 25344
rect 7708 25304 7714 25316
rect 8570 25304 8576 25316
rect 8628 25304 8634 25356
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 8680 25316 9689 25344
rect 7190 25276 7196 25288
rect 5736 25248 7196 25276
rect 7190 25236 7196 25248
rect 7248 25276 7254 25288
rect 7248 25248 7420 25276
rect 7248 25236 7254 25248
rect 4522 25168 4528 25220
rect 4580 25168 4586 25220
rect 6086 25168 6092 25220
rect 6144 25168 6150 25220
rect 7392 25217 7420 25248
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8680 25276 8708 25316
rect 9677 25313 9689 25316
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 12250 25304 12256 25356
rect 12308 25304 12314 25356
rect 8352 25248 8708 25276
rect 11793 25279 11851 25285
rect 8352 25236 8358 25248
rect 11793 25245 11805 25279
rect 11839 25245 11851 25279
rect 11793 25239 11851 25245
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25276 12035 25279
rect 12023 25248 12296 25276
rect 12023 25245 12035 25248
rect 11977 25239 12035 25245
rect 7377 25211 7435 25217
rect 7377 25177 7389 25211
rect 7423 25177 7435 25211
rect 7377 25171 7435 25177
rect 7561 25211 7619 25217
rect 7561 25177 7573 25211
rect 7607 25208 7619 25211
rect 7650 25208 7656 25220
rect 7607 25180 7656 25208
rect 7607 25177 7619 25180
rect 7561 25171 7619 25177
rect 7650 25168 7656 25180
rect 7708 25168 7714 25220
rect 8938 25208 8944 25220
rect 8128 25180 8944 25208
rect 3421 25143 3479 25149
rect 3421 25109 3433 25143
rect 3467 25140 3479 25143
rect 8128 25140 8156 25180
rect 8938 25168 8944 25180
rect 8996 25168 9002 25220
rect 9493 25211 9551 25217
rect 9493 25177 9505 25211
rect 9539 25208 9551 25211
rect 9674 25208 9680 25220
rect 9539 25180 9680 25208
rect 9539 25177 9551 25180
rect 9493 25171 9551 25177
rect 9674 25168 9680 25180
rect 9732 25208 9738 25220
rect 11698 25208 11704 25220
rect 9732 25180 11704 25208
rect 9732 25168 9738 25180
rect 11698 25168 11704 25180
rect 11756 25208 11762 25220
rect 11808 25208 11836 25239
rect 11756 25180 11836 25208
rect 11885 25211 11943 25217
rect 11756 25168 11762 25180
rect 11885 25177 11897 25211
rect 11931 25177 11943 25211
rect 11885 25171 11943 25177
rect 3467 25112 8156 25140
rect 3467 25109 3479 25112
rect 3421 25103 3479 25109
rect 8202 25100 8208 25152
rect 8260 25140 8266 25152
rect 9585 25143 9643 25149
rect 9585 25140 9597 25143
rect 8260 25112 9597 25140
rect 8260 25100 8266 25112
rect 9585 25109 9597 25112
rect 9631 25140 9643 25143
rect 10042 25140 10048 25152
rect 9631 25112 10048 25140
rect 9631 25109 9643 25112
rect 9585 25103 9643 25109
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 10962 25100 10968 25152
rect 11020 25140 11026 25152
rect 11900 25140 11928 25171
rect 12066 25168 12072 25220
rect 12124 25217 12130 25220
rect 12124 25211 12153 25217
rect 12141 25177 12153 25211
rect 12268 25208 12296 25248
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 13004 25285 13032 25384
rect 12805 25279 12863 25285
rect 12805 25276 12817 25279
rect 12400 25248 12817 25276
rect 12400 25236 12406 25248
rect 12805 25245 12817 25248
rect 12851 25245 12863 25279
rect 12805 25239 12863 25245
rect 12989 25279 13047 25285
rect 12989 25245 13001 25279
rect 13035 25245 13047 25279
rect 25332 25276 25360 25443
rect 25958 25440 25964 25492
rect 26016 25440 26022 25492
rect 25869 25279 25927 25285
rect 25869 25276 25881 25279
rect 25332 25248 25881 25276
rect 12989 25239 13047 25245
rect 25869 25245 25881 25248
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 26970 25236 26976 25288
rect 27028 25236 27034 25288
rect 12434 25208 12440 25220
rect 12268 25180 12440 25208
rect 12124 25171 12153 25177
rect 12124 25168 12130 25171
rect 12434 25168 12440 25180
rect 12492 25168 12498 25220
rect 13170 25168 13176 25220
rect 13228 25168 13234 25220
rect 25682 25168 25688 25220
rect 25740 25168 25746 25220
rect 27246 25217 27252 25220
rect 27240 25208 27252 25217
rect 27207 25180 27252 25208
rect 27240 25171 27252 25180
rect 27246 25168 27252 25171
rect 27304 25168 27310 25220
rect 11020 25112 11928 25140
rect 11020 25100 11026 25112
rect 27522 25100 27528 25152
rect 27580 25140 27586 25152
rect 28353 25143 28411 25149
rect 28353 25140 28365 25143
rect 27580 25112 28365 25140
rect 27580 25100 27586 25112
rect 28353 25109 28365 25112
rect 28399 25109 28411 25143
rect 28353 25103 28411 25109
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 3786 24896 3792 24948
rect 3844 24936 3850 24948
rect 3844 24908 4108 24936
rect 3844 24896 3850 24908
rect 3142 24828 3148 24880
rect 3200 24828 3206 24880
rect 2000 24803 2058 24809
rect 2000 24769 2012 24803
rect 2046 24800 2058 24803
rect 2682 24800 2688 24812
rect 2046 24772 2688 24800
rect 2046 24769 2058 24772
rect 2000 24763 2058 24769
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 2958 24760 2964 24812
rect 3016 24760 3022 24812
rect 3804 24809 3832 24896
rect 3789 24803 3847 24809
rect 3789 24769 3801 24803
rect 3835 24769 3847 24803
rect 3789 24763 3847 24769
rect 3878 24760 3884 24812
rect 3936 24798 3942 24812
rect 3973 24803 4031 24809
rect 3973 24798 3985 24803
rect 3936 24770 3985 24798
rect 3936 24760 3942 24770
rect 3973 24769 3985 24770
rect 4019 24769 4031 24803
rect 4080 24800 4108 24908
rect 4522 24896 4528 24948
rect 4580 24936 4586 24948
rect 5445 24939 5503 24945
rect 4580 24908 5396 24936
rect 4580 24896 4586 24908
rect 5368 24868 5396 24908
rect 5445 24905 5457 24939
rect 5491 24936 5503 24939
rect 5626 24936 5632 24948
rect 5491 24908 5632 24936
rect 5491 24905 5503 24908
rect 5445 24899 5503 24905
rect 5626 24896 5632 24908
rect 5684 24936 5690 24948
rect 6086 24936 6092 24948
rect 5684 24908 6092 24936
rect 5684 24896 5690 24908
rect 6086 24896 6092 24908
rect 6144 24896 6150 24948
rect 7650 24936 7656 24948
rect 7484 24908 7656 24936
rect 7484 24868 7512 24908
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 10226 24896 10232 24948
rect 10284 24896 10290 24948
rect 11054 24896 11060 24948
rect 11112 24936 11118 24948
rect 11885 24939 11943 24945
rect 11885 24936 11897 24939
rect 11112 24908 11897 24936
rect 11112 24896 11118 24908
rect 11885 24905 11897 24908
rect 11931 24905 11943 24939
rect 11885 24899 11943 24905
rect 4540 24840 4752 24868
rect 5368 24840 7512 24868
rect 4433 24803 4491 24809
rect 4433 24800 4445 24803
rect 4080 24772 4445 24800
rect 3973 24763 4031 24769
rect 4433 24769 4445 24772
rect 4479 24800 4491 24803
rect 4540 24800 4568 24840
rect 4479 24772 4568 24800
rect 4479 24769 4491 24772
rect 4433 24763 4491 24769
rect 4614 24760 4620 24812
rect 4672 24760 4678 24812
rect 4724 24800 4752 24840
rect 7558 24828 7564 24880
rect 7616 24868 7622 24880
rect 12158 24868 12164 24880
rect 7616 24840 12164 24868
rect 7616 24828 7622 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 12434 24828 12440 24880
rect 12492 24868 12498 24880
rect 12492 24840 13124 24868
rect 12492 24828 12498 24840
rect 5353 24803 5411 24809
rect 4724 24772 5304 24800
rect 1854 24692 1860 24744
rect 1912 24732 1918 24744
rect 2087 24735 2145 24741
rect 2087 24732 2099 24735
rect 1912 24704 2099 24732
rect 1912 24692 1918 24704
rect 2087 24701 2099 24704
rect 2133 24701 2145 24735
rect 2087 24695 2145 24701
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24732 3295 24735
rect 4982 24732 4988 24744
rect 3283 24704 4988 24732
rect 3283 24701 3295 24704
rect 3237 24695 3295 24701
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 2685 24667 2743 24673
rect 2685 24633 2697 24667
rect 2731 24664 2743 24667
rect 4062 24664 4068 24676
rect 2731 24636 4068 24664
rect 2731 24633 2743 24636
rect 2685 24627 2743 24633
rect 4062 24624 4068 24636
rect 4120 24624 4126 24676
rect 4614 24624 4620 24676
rect 4672 24664 4678 24676
rect 4890 24664 4896 24676
rect 4672 24636 4896 24664
rect 4672 24624 4678 24636
rect 4890 24624 4896 24636
rect 4948 24624 4954 24676
rect 5276 24664 5304 24772
rect 5353 24769 5365 24803
rect 5399 24800 5411 24803
rect 5442 24800 5448 24812
rect 5399 24772 5448 24800
rect 5399 24769 5411 24772
rect 5353 24763 5411 24769
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 5537 24803 5595 24809
rect 5537 24769 5549 24803
rect 5583 24800 5595 24803
rect 5810 24800 5816 24812
rect 5583 24772 5816 24800
rect 5583 24769 5595 24772
rect 5537 24763 5595 24769
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 10229 24803 10287 24809
rect 10229 24800 10241 24803
rect 10192 24772 10241 24800
rect 10192 24760 10198 24772
rect 10229 24769 10241 24772
rect 10275 24769 10287 24803
rect 10962 24800 10968 24812
rect 10229 24763 10287 24769
rect 10428 24772 10968 24800
rect 7742 24732 7748 24744
rect 6104 24704 7748 24732
rect 6104 24664 6132 24704
rect 7742 24692 7748 24704
rect 7800 24692 7806 24744
rect 10045 24735 10103 24741
rect 10045 24701 10057 24735
rect 10091 24732 10103 24735
rect 10428 24732 10456 24772
rect 10962 24760 10968 24772
rect 11020 24760 11026 24812
rect 11054 24760 11060 24812
rect 11112 24800 11118 24812
rect 11790 24800 11796 24812
rect 11112 24772 11796 24800
rect 11112 24760 11118 24772
rect 11790 24760 11796 24772
rect 11848 24800 11854 24812
rect 11885 24803 11943 24809
rect 11885 24800 11897 24803
rect 11848 24772 11897 24800
rect 11848 24760 11854 24772
rect 11885 24769 11897 24772
rect 11931 24769 11943 24803
rect 12250 24800 12256 24812
rect 12211 24772 12256 24800
rect 11885 24763 11943 24769
rect 12250 24760 12256 24772
rect 12308 24800 12314 24812
rect 13096 24809 13124 24840
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12308 24772 12909 24800
rect 12308 24760 12314 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 14553 24803 14611 24809
rect 14553 24769 14565 24803
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 10091 24704 10456 24732
rect 10091 24701 10103 24704
rect 10045 24695 10103 24701
rect 5276 24636 6132 24664
rect 6178 24624 6184 24676
rect 6236 24664 6242 24676
rect 10060 24664 10088 24695
rect 10502 24692 10508 24744
rect 10560 24732 10566 24744
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 10560 24704 10609 24732
rect 10560 24692 10566 24704
rect 10597 24701 10609 24704
rect 10643 24701 10655 24735
rect 10980 24732 11008 24760
rect 11701 24735 11759 24741
rect 11701 24732 11713 24735
rect 10980 24704 11713 24732
rect 10597 24695 10655 24701
rect 11701 24701 11713 24704
rect 11747 24732 11759 24735
rect 11974 24732 11980 24744
rect 11747 24704 11980 24732
rect 11747 24701 11759 24704
rect 11701 24695 11759 24701
rect 11974 24692 11980 24704
rect 12032 24732 12038 24744
rect 13188 24732 13216 24763
rect 12032 24704 13216 24732
rect 14568 24732 14596 24763
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 16482 24760 16488 24812
rect 16540 24800 16546 24812
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 16540 24772 16865 24800
rect 16540 24760 16546 24772
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 17034 24760 17040 24812
rect 17092 24760 17098 24812
rect 17218 24760 17224 24812
rect 17276 24760 17282 24812
rect 15562 24732 15568 24744
rect 14568 24704 15568 24732
rect 12032 24692 12038 24704
rect 15562 24692 15568 24704
rect 15620 24732 15626 24744
rect 16022 24732 16028 24744
rect 15620 24704 16028 24732
rect 15620 24692 15626 24704
rect 16022 24692 16028 24704
rect 16080 24692 16086 24744
rect 10226 24664 10232 24676
rect 6236 24636 10232 24664
rect 6236 24624 6242 24636
rect 10226 24624 10232 24636
rect 10284 24624 10290 24676
rect 14369 24667 14427 24673
rect 14369 24664 14381 24667
rect 12406 24636 14381 24664
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 12406 24596 12434 24636
rect 14369 24633 14381 24636
rect 14415 24633 14427 24667
rect 14369 24627 14427 24633
rect 9732 24568 12434 24596
rect 9732 24556 9738 24568
rect 12710 24556 12716 24608
rect 12768 24556 12774 24608
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 2130 24352 2136 24404
rect 2188 24392 2194 24404
rect 2915 24395 2973 24401
rect 2915 24392 2927 24395
rect 2188 24364 2927 24392
rect 2188 24352 2194 24364
rect 2915 24361 2927 24364
rect 2961 24361 2973 24395
rect 2915 24355 2973 24361
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 9306 24392 9312 24404
rect 3936 24364 9312 24392
rect 3936 24352 3942 24364
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 10226 24352 10232 24404
rect 10284 24352 10290 24404
rect 16574 24352 16580 24404
rect 16632 24352 16638 24404
rect 4154 24324 4160 24336
rect 2424 24296 4160 24324
rect 1486 24148 1492 24200
rect 1544 24188 1550 24200
rect 1544 24160 1716 24188
rect 1544 24148 1550 24160
rect 842 24080 848 24132
rect 900 24120 906 24132
rect 1581 24123 1639 24129
rect 1581 24120 1593 24123
rect 900 24092 1593 24120
rect 900 24080 906 24092
rect 1581 24089 1593 24092
rect 1627 24089 1639 24123
rect 1688 24120 1716 24160
rect 1762 24148 1768 24200
rect 1820 24148 1826 24200
rect 2021 24191 2079 24197
rect 2021 24157 2033 24191
rect 2067 24188 2079 24191
rect 2222 24188 2228 24200
rect 2067 24160 2228 24188
rect 2067 24157 2079 24160
rect 2021 24151 2079 24157
rect 2222 24148 2228 24160
rect 2280 24148 2286 24200
rect 2314 24148 2320 24200
rect 2372 24148 2378 24200
rect 2424 24120 2452 24296
rect 4154 24284 4160 24296
rect 4212 24284 4218 24336
rect 4338 24284 4344 24336
rect 4396 24324 4402 24336
rect 5169 24327 5227 24333
rect 5169 24324 5181 24327
rect 4396 24296 5181 24324
rect 4396 24284 4402 24296
rect 5169 24293 5181 24296
rect 5215 24293 5227 24327
rect 10686 24324 10692 24336
rect 5169 24287 5227 24293
rect 8772 24296 10692 24324
rect 3142 24216 3148 24268
rect 3200 24256 3206 24268
rect 8772 24256 8800 24296
rect 10686 24284 10692 24296
rect 10744 24324 10750 24336
rect 10744 24296 12940 24324
rect 10744 24284 10750 24296
rect 3200 24228 8800 24256
rect 11609 24259 11667 24265
rect 3200 24216 3206 24228
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 11698 24256 11704 24268
rect 11655 24228 11704 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 11698 24216 11704 24228
rect 11756 24216 11762 24268
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 12032 24228 12848 24256
rect 12032 24216 12038 24228
rect 2682 24148 2688 24200
rect 2740 24188 2746 24200
rect 2812 24191 2870 24197
rect 2812 24188 2824 24191
rect 2740 24160 2824 24188
rect 2740 24148 2746 24160
rect 2812 24157 2824 24160
rect 2858 24157 2870 24191
rect 2812 24151 2870 24157
rect 4522 24148 4528 24200
rect 4580 24148 4586 24200
rect 4890 24148 4896 24200
rect 4948 24148 4954 24200
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24188 5319 24191
rect 5718 24188 5724 24200
rect 5307 24160 5724 24188
rect 5307 24157 5319 24160
rect 5261 24151 5319 24157
rect 1688 24092 2452 24120
rect 1581 24083 1639 24089
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 2038 24052 2044 24064
rect 1912 24024 2044 24052
rect 1912 24012 1918 24024
rect 2038 24012 2044 24024
rect 2096 24052 2102 24064
rect 2240 24061 2268 24092
rect 4062 24080 4068 24132
rect 4120 24120 4126 24132
rect 5276 24120 5304 24151
rect 5718 24148 5724 24160
rect 5776 24148 5782 24200
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 8294 24188 8300 24200
rect 6595 24160 8300 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 8294 24148 8300 24160
rect 8352 24148 8358 24200
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 10137 24191 10195 24197
rect 10137 24188 10149 24191
rect 10008 24160 10149 24188
rect 10008 24148 10014 24160
rect 10137 24157 10149 24160
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 10502 24148 10508 24200
rect 10560 24188 10566 24200
rect 11241 24191 11299 24197
rect 11241 24188 11253 24191
rect 10560 24160 11253 24188
rect 10560 24148 10566 24160
rect 11241 24157 11253 24160
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24188 11575 24191
rect 12066 24188 12072 24200
rect 11563 24160 12072 24188
rect 11563 24157 11575 24160
rect 11517 24151 11575 24157
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12820 24197 12848 24228
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12308 24160 12541 24188
rect 12308 24148 12314 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24157 12863 24191
rect 12805 24151 12863 24157
rect 6270 24120 6276 24132
rect 4120 24092 5304 24120
rect 5368 24092 6276 24120
rect 4120 24080 4126 24092
rect 2133 24055 2191 24061
rect 2133 24052 2145 24055
rect 2096 24024 2145 24052
rect 2096 24012 2102 24024
rect 2133 24021 2145 24024
rect 2179 24021 2191 24055
rect 2133 24015 2191 24021
rect 2225 24055 2283 24061
rect 2225 24021 2237 24055
rect 2271 24021 2283 24055
rect 2225 24015 2283 24021
rect 2314 24012 2320 24064
rect 2372 24052 2378 24064
rect 4522 24052 4528 24064
rect 2372 24024 4528 24052
rect 2372 24012 2378 24024
rect 4522 24012 4528 24024
rect 4580 24052 4586 24064
rect 5368 24052 5396 24092
rect 6270 24080 6276 24092
rect 6328 24080 6334 24132
rect 6365 24123 6423 24129
rect 6365 24089 6377 24123
rect 6411 24120 6423 24123
rect 6638 24120 6644 24132
rect 6411 24092 6644 24120
rect 6411 24089 6423 24092
rect 6365 24083 6423 24089
rect 6638 24080 6644 24092
rect 6696 24080 6702 24132
rect 10962 24080 10968 24132
rect 11020 24120 11026 24132
rect 12345 24123 12403 24129
rect 12345 24120 12357 24123
rect 11020 24092 12357 24120
rect 11020 24080 11026 24092
rect 12345 24089 12357 24092
rect 12391 24120 12403 24123
rect 12618 24120 12624 24132
rect 12391 24092 12624 24120
rect 12391 24089 12403 24092
rect 12345 24083 12403 24089
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 12713 24123 12771 24129
rect 12713 24089 12725 24123
rect 12759 24120 12771 24123
rect 12912 24120 12940 24296
rect 20714 24216 20720 24268
rect 20772 24256 20778 24268
rect 20993 24259 21051 24265
rect 20993 24256 21005 24259
rect 20772 24228 21005 24256
rect 20772 24216 20778 24228
rect 20993 24225 21005 24228
rect 21039 24225 21051 24259
rect 20993 24219 21051 24225
rect 13262 24148 13268 24200
rect 13320 24188 13326 24200
rect 16482 24188 16488 24200
rect 13320 24160 16488 24188
rect 13320 24148 13326 24160
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24188 16727 24191
rect 17034 24188 17040 24200
rect 16715 24160 17040 24188
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 16114 24120 16120 24132
rect 12759 24092 16120 24120
rect 12759 24089 12771 24092
rect 12713 24083 12771 24089
rect 16114 24080 16120 24092
rect 16172 24120 16178 24132
rect 16684 24120 16712 24151
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 24578 24148 24584 24200
rect 24636 24188 24642 24200
rect 25130 24188 25136 24200
rect 24636 24160 25136 24188
rect 24636 24148 24642 24160
rect 25130 24148 25136 24160
rect 25188 24188 25194 24200
rect 26970 24188 26976 24200
rect 25188 24160 26976 24188
rect 25188 24148 25194 24160
rect 26970 24148 26976 24160
rect 27028 24148 27034 24200
rect 16172 24092 16712 24120
rect 16172 24080 16178 24092
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 21238 24123 21296 24129
rect 21238 24120 21250 24123
rect 19208 24092 21250 24120
rect 19208 24080 19214 24092
rect 21238 24089 21250 24092
rect 21284 24120 21296 24123
rect 23198 24120 23204 24132
rect 21284 24092 23204 24120
rect 21284 24089 21296 24092
rect 21238 24083 21296 24089
rect 23198 24080 23204 24092
rect 23256 24080 23262 24132
rect 27240 24123 27298 24129
rect 27240 24089 27252 24123
rect 27286 24120 27298 24123
rect 27338 24120 27344 24132
rect 27286 24092 27344 24120
rect 27286 24089 27298 24092
rect 27240 24083 27298 24089
rect 27338 24080 27344 24092
rect 27396 24080 27402 24132
rect 4580 24024 5396 24052
rect 4580 24012 4586 24024
rect 5718 24012 5724 24064
rect 5776 24052 5782 24064
rect 6733 24055 6791 24061
rect 6733 24052 6745 24055
rect 5776 24024 6745 24052
rect 5776 24012 5782 24024
rect 6733 24021 6745 24024
rect 6779 24021 6791 24055
rect 6733 24015 6791 24021
rect 21542 24012 21548 24064
rect 21600 24052 21606 24064
rect 22373 24055 22431 24061
rect 22373 24052 22385 24055
rect 21600 24024 22385 24052
rect 21600 24012 21606 24024
rect 22373 24021 22385 24024
rect 22419 24021 22431 24055
rect 22373 24015 22431 24021
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 28353 24055 28411 24061
rect 28353 24052 28365 24055
rect 24176 24024 28365 24052
rect 24176 24012 24182 24024
rect 28353 24021 28365 24024
rect 28399 24021 28411 24055
rect 28353 24015 28411 24021
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 4065 23851 4123 23857
rect 4065 23817 4077 23851
rect 4111 23848 4123 23851
rect 4982 23848 4988 23860
rect 4111 23820 4988 23848
rect 4111 23817 4123 23820
rect 4065 23811 4123 23817
rect 4982 23808 4988 23820
rect 5040 23808 5046 23860
rect 5442 23808 5448 23860
rect 5500 23808 5506 23860
rect 6362 23808 6368 23860
rect 6420 23848 6426 23860
rect 6749 23851 6807 23857
rect 6749 23848 6761 23851
rect 6420 23820 6761 23848
rect 6420 23808 6426 23820
rect 6749 23817 6761 23820
rect 6795 23817 6807 23851
rect 6749 23811 6807 23817
rect 7006 23808 7012 23860
rect 7064 23848 7070 23860
rect 7834 23848 7840 23860
rect 7064 23820 7840 23848
rect 7064 23808 7070 23820
rect 7834 23808 7840 23820
rect 7892 23808 7898 23860
rect 8294 23808 8300 23860
rect 8352 23848 8358 23860
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 8352 23820 9873 23848
rect 8352 23808 8358 23820
rect 9861 23817 9873 23820
rect 9907 23817 9919 23851
rect 9861 23811 9919 23817
rect 2590 23740 2596 23792
rect 2648 23740 2654 23792
rect 4706 23740 4712 23792
rect 4764 23780 4770 23792
rect 4801 23783 4859 23789
rect 4801 23780 4813 23783
rect 4764 23752 4813 23780
rect 4764 23740 4770 23752
rect 4801 23749 4813 23752
rect 4847 23749 4859 23783
rect 5460 23780 5488 23808
rect 4801 23743 4859 23749
rect 5368 23752 5488 23780
rect 3602 23672 3608 23724
rect 3660 23712 3666 23724
rect 4982 23712 4988 23724
rect 3660 23684 4988 23712
rect 3660 23672 3666 23684
rect 4982 23672 4988 23684
rect 5040 23712 5046 23724
rect 5077 23715 5135 23721
rect 5077 23712 5089 23715
rect 5040 23684 5089 23712
rect 5040 23672 5046 23684
rect 5077 23681 5089 23684
rect 5123 23681 5135 23715
rect 5077 23675 5135 23681
rect 5169 23715 5227 23721
rect 5169 23681 5181 23715
rect 5215 23681 5227 23715
rect 5169 23675 5227 23681
rect 5184 23644 5212 23675
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5368 23712 5396 23752
rect 5810 23740 5816 23792
rect 5868 23780 5874 23792
rect 6549 23783 6607 23789
rect 6549 23780 6561 23783
rect 5868 23752 6561 23780
rect 5868 23740 5874 23752
rect 6549 23749 6561 23752
rect 6595 23780 6607 23783
rect 7098 23780 7104 23792
rect 6595 23752 7104 23780
rect 6595 23749 6607 23752
rect 6549 23743 6607 23749
rect 7098 23740 7104 23752
rect 7156 23740 7162 23792
rect 7469 23783 7527 23789
rect 7469 23749 7481 23783
rect 7515 23780 7527 23783
rect 10594 23780 10600 23792
rect 7515 23752 10600 23780
rect 7515 23749 7527 23752
rect 7469 23743 7527 23749
rect 10594 23740 10600 23752
rect 10652 23740 10658 23792
rect 14734 23780 14740 23792
rect 12406 23752 14740 23780
rect 5316 23684 5396 23712
rect 5316 23672 5322 23684
rect 5442 23672 5448 23724
rect 5500 23672 5506 23724
rect 7190 23672 7196 23724
rect 7248 23712 7254 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7248 23684 7665 23712
rect 7248 23672 7254 23684
rect 7653 23681 7665 23684
rect 7699 23712 7711 23715
rect 9766 23712 9772 23724
rect 7699 23684 9772 23712
rect 7699 23681 7711 23684
rect 7653 23675 7711 23681
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 9858 23672 9864 23724
rect 9916 23672 9922 23724
rect 11146 23672 11152 23724
rect 11204 23712 11210 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11204 23684 11897 23712
rect 11204 23672 11210 23684
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 5810 23644 5816 23656
rect 5184 23616 5816 23644
rect 5810 23604 5816 23616
rect 5868 23604 5874 23656
rect 6454 23604 6460 23656
rect 6512 23644 6518 23656
rect 9677 23647 9735 23653
rect 6512 23616 9628 23644
rect 6512 23604 6518 23616
rect 8386 23576 8392 23588
rect 2746 23548 8392 23576
rect 1765 23511 1823 23517
rect 1765 23477 1777 23511
rect 1811 23508 1823 23511
rect 2746 23508 2774 23548
rect 8386 23536 8392 23548
rect 8444 23536 8450 23588
rect 9600 23576 9628 23616
rect 9677 23613 9689 23647
rect 9723 23644 9735 23647
rect 10134 23644 10140 23656
rect 9723 23616 10140 23644
rect 9723 23613 9735 23616
rect 9677 23607 9735 23613
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 10229 23647 10287 23653
rect 10229 23613 10241 23647
rect 10275 23644 10287 23647
rect 10502 23644 10508 23656
rect 10275 23616 10508 23644
rect 10275 23613 10287 23616
rect 10229 23607 10287 23613
rect 10244 23576 10272 23607
rect 10502 23604 10508 23616
rect 10560 23644 10566 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 10560 23616 12173 23644
rect 10560 23604 10566 23616
rect 12161 23613 12173 23616
rect 12207 23644 12219 23647
rect 12250 23644 12256 23656
rect 12207 23616 12256 23644
rect 12207 23613 12219 23616
rect 12161 23607 12219 23613
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 12406 23576 12434 23752
rect 14734 23740 14740 23752
rect 14792 23740 14798 23792
rect 24394 23780 24400 23792
rect 22066 23752 24400 23780
rect 14550 23672 14556 23724
rect 14608 23672 14614 23724
rect 14820 23715 14878 23721
rect 14820 23681 14832 23715
rect 14866 23712 14878 23715
rect 16298 23712 16304 23724
rect 14866 23684 16304 23712
rect 14866 23681 14878 23684
rect 14820 23675 14878 23681
rect 16298 23672 16304 23684
rect 16356 23672 16362 23724
rect 21174 23604 21180 23656
rect 21232 23644 21238 23656
rect 22066 23644 22094 23752
rect 24394 23740 24400 23752
rect 24452 23780 24458 23792
rect 25010 23783 25068 23789
rect 25010 23780 25022 23783
rect 24452 23752 25022 23780
rect 24452 23740 24458 23752
rect 25010 23749 25022 23752
rect 25056 23749 25068 23783
rect 25010 23743 25068 23749
rect 21232 23616 22094 23644
rect 21232 23604 21238 23616
rect 24578 23604 24584 23656
rect 24636 23644 24642 23656
rect 24765 23647 24823 23653
rect 24765 23644 24777 23647
rect 24636 23616 24777 23644
rect 24636 23604 24642 23616
rect 24765 23613 24777 23616
rect 24811 23613 24823 23647
rect 24765 23607 24823 23613
rect 9600 23548 10272 23576
rect 11992 23548 12434 23576
rect 1811 23480 2774 23508
rect 1811 23477 1823 23480
rect 1765 23471 1823 23477
rect 4154 23468 4160 23520
rect 4212 23508 4218 23520
rect 6454 23508 6460 23520
rect 4212 23480 6460 23508
rect 4212 23468 4218 23480
rect 6454 23468 6460 23480
rect 6512 23468 6518 23520
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 6733 23511 6791 23517
rect 6733 23508 6745 23511
rect 6696 23480 6745 23508
rect 6696 23468 6702 23480
rect 6733 23477 6745 23480
rect 6779 23477 6791 23511
rect 6733 23471 6791 23477
rect 6914 23468 6920 23520
rect 6972 23468 6978 23520
rect 7834 23468 7840 23520
rect 7892 23508 7898 23520
rect 11992 23508 12020 23548
rect 7892 23480 12020 23508
rect 7892 23468 7898 23480
rect 12066 23468 12072 23520
rect 12124 23508 12130 23520
rect 15562 23508 15568 23520
rect 12124 23480 15568 23508
rect 12124 23468 12130 23480
rect 15562 23468 15568 23480
rect 15620 23468 15626 23520
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16022 23508 16028 23520
rect 15979 23480 16028 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 26050 23468 26056 23520
rect 26108 23508 26114 23520
rect 26145 23511 26203 23517
rect 26145 23508 26157 23511
rect 26108 23480 26157 23508
rect 26108 23468 26114 23480
rect 26145 23477 26157 23480
rect 26191 23477 26203 23511
rect 26145 23471 26203 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 1578 23264 1584 23316
rect 1636 23304 1642 23316
rect 11698 23304 11704 23316
rect 1636 23276 11704 23304
rect 1636 23264 1642 23276
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 11793 23307 11851 23313
rect 11793 23273 11805 23307
rect 11839 23304 11851 23307
rect 11974 23304 11980 23316
rect 11839 23276 11980 23304
rect 11839 23273 11851 23276
rect 11793 23267 11851 23273
rect 11974 23264 11980 23276
rect 12032 23304 12038 23316
rect 12342 23304 12348 23316
rect 12032 23276 12348 23304
rect 12032 23264 12038 23276
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 12526 23264 12532 23316
rect 12584 23264 12590 23316
rect 5350 23196 5356 23248
rect 5408 23236 5414 23248
rect 9030 23236 9036 23248
rect 5408 23208 9036 23236
rect 5408 23196 5414 23208
rect 9030 23196 9036 23208
rect 9088 23196 9094 23248
rect 9950 23196 9956 23248
rect 10008 23236 10014 23248
rect 10137 23239 10195 23245
rect 10137 23236 10149 23239
rect 10008 23208 10149 23236
rect 10008 23196 10014 23208
rect 10137 23205 10149 23208
rect 10183 23205 10195 23239
rect 10137 23199 10195 23205
rect 5534 23168 5540 23180
rect 4908 23140 5540 23168
rect 4908 23109 4936 23140
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 5626 23128 5632 23180
rect 5684 23128 5690 23180
rect 5721 23171 5779 23177
rect 5721 23137 5733 23171
rect 5767 23168 5779 23171
rect 6178 23168 6184 23180
rect 5767 23140 6184 23168
rect 5767 23137 5779 23140
rect 5721 23131 5779 23137
rect 6178 23128 6184 23140
rect 6236 23168 6242 23180
rect 6638 23168 6644 23180
rect 6236 23140 6644 23168
rect 6236 23128 6242 23140
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 9766 23128 9772 23180
rect 9824 23168 9830 23180
rect 10410 23168 10416 23180
rect 9824 23140 10416 23168
rect 9824 23128 9830 23140
rect 10410 23128 10416 23140
rect 10468 23128 10474 23180
rect 24578 23128 24584 23180
rect 24636 23168 24642 23180
rect 25869 23171 25927 23177
rect 25869 23168 25881 23171
rect 24636 23140 25881 23168
rect 24636 23128 24642 23140
rect 25869 23137 25881 23140
rect 25915 23137 25927 23171
rect 25869 23131 25927 23137
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23069 5135 23103
rect 5077 23063 5135 23069
rect 4154 22992 4160 23044
rect 4212 23032 4218 23044
rect 4341 23035 4399 23041
rect 4341 23032 4353 23035
rect 4212 23004 4353 23032
rect 4212 22992 4218 23004
rect 4341 23001 4353 23004
rect 4387 23001 4399 23035
rect 5092 23032 5120 23063
rect 5258 23060 5264 23112
rect 5316 23060 5322 23112
rect 9950 23060 9956 23112
rect 10008 23060 10014 23112
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 10870 23100 10876 23112
rect 10652 23072 10876 23100
rect 10652 23060 10658 23072
rect 10870 23060 10876 23072
rect 10928 23100 10934 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 10928 23072 11529 23100
rect 10928 23060 10934 23072
rect 11517 23069 11529 23072
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 12342 23060 12348 23112
rect 12400 23060 12406 23112
rect 13262 23060 13268 23112
rect 13320 23060 13326 23112
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23100 17279 23103
rect 18230 23100 18236 23112
rect 17267 23072 18236 23100
rect 17267 23069 17279 23072
rect 17221 23063 17279 23069
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21269 23103 21327 23109
rect 21269 23100 21281 23103
rect 20772 23072 21281 23100
rect 20772 23060 20778 23072
rect 21269 23069 21281 23072
rect 21315 23069 21327 23103
rect 21269 23063 21327 23069
rect 6178 23032 6184 23044
rect 5092 23004 6184 23032
rect 4341 22995 4399 23001
rect 6178 22992 6184 23004
rect 6236 22992 6242 23044
rect 12894 22992 12900 23044
rect 12952 23032 12958 23044
rect 14550 23032 14556 23044
rect 12952 23004 14556 23032
rect 12952 22992 12958 23004
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 17488 23035 17546 23041
rect 17488 23001 17500 23035
rect 17534 23032 17546 23035
rect 17954 23032 17960 23044
rect 17534 23004 17960 23032
rect 17534 23001 17546 23004
rect 17488 22995 17546 23001
rect 17954 22992 17960 23004
rect 18012 22992 18018 23044
rect 26136 23035 26194 23041
rect 26136 23001 26148 23035
rect 26182 23001 26194 23035
rect 26136 22995 26194 23001
rect 6638 22924 6644 22976
rect 6696 22964 6702 22976
rect 9674 22964 9680 22976
rect 6696 22936 9680 22964
rect 6696 22924 6702 22936
rect 9674 22924 9680 22936
rect 9732 22924 9738 22976
rect 12802 22924 12808 22976
rect 12860 22924 12866 22976
rect 13354 22924 13360 22976
rect 13412 22924 13418 22976
rect 18138 22924 18144 22976
rect 18196 22964 18202 22976
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 18196 22936 18613 22964
rect 18196 22924 18202 22936
rect 18601 22933 18613 22936
rect 18647 22933 18659 22967
rect 18601 22927 18659 22933
rect 21453 22967 21511 22973
rect 21453 22933 21465 22967
rect 21499 22964 21511 22967
rect 21634 22964 21640 22976
rect 21499 22936 21640 22964
rect 21499 22933 21511 22936
rect 21453 22927 21511 22933
rect 21634 22924 21640 22936
rect 21692 22924 21698 22976
rect 26050 22924 26056 22976
rect 26108 22964 26114 22976
rect 26160 22964 26188 22995
rect 26108 22936 26188 22964
rect 26108 22924 26114 22936
rect 27246 22924 27252 22976
rect 27304 22924 27310 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 4890 22720 4896 22772
rect 4948 22760 4954 22772
rect 10502 22760 10508 22772
rect 4948 22732 10508 22760
rect 4948 22720 4954 22732
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 11698 22720 11704 22772
rect 11756 22720 11762 22772
rect 12069 22763 12127 22769
rect 12069 22729 12081 22763
rect 12115 22760 12127 22763
rect 13354 22760 13360 22772
rect 12115 22732 13360 22760
rect 12115 22729 12127 22732
rect 12069 22723 12127 22729
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 16022 22760 16028 22772
rect 13832 22732 16028 22760
rect 6917 22695 6975 22701
rect 6917 22661 6929 22695
rect 6963 22692 6975 22695
rect 7561 22695 7619 22701
rect 7561 22692 7573 22695
rect 6963 22664 7573 22692
rect 6963 22661 6975 22664
rect 6917 22655 6975 22661
rect 7561 22661 7573 22664
rect 7607 22661 7619 22695
rect 7561 22655 7619 22661
rect 9944 22695 10002 22701
rect 9944 22661 9956 22695
rect 9990 22692 10002 22695
rect 13722 22692 13728 22704
rect 9990 22664 13728 22692
rect 9990 22661 10002 22664
rect 9944 22655 10002 22661
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 4890 22584 4896 22636
rect 4948 22624 4954 22636
rect 6733 22627 6791 22633
rect 6733 22624 6745 22627
rect 4948 22596 6745 22624
rect 4948 22584 4954 22596
rect 6733 22593 6745 22596
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 2498 22516 2504 22568
rect 2556 22556 2562 22568
rect 6638 22556 6644 22568
rect 2556 22528 6644 22556
rect 2556 22516 2562 22528
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 1394 22380 1400 22432
rect 1452 22420 1458 22432
rect 6549 22423 6607 22429
rect 6549 22420 6561 22423
rect 1452 22392 6561 22420
rect 1452 22380 1458 22392
rect 6549 22389 6561 22392
rect 6595 22389 6607 22423
rect 6748 22420 6776 22587
rect 7006 22584 7012 22636
rect 7064 22584 7070 22636
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 7248 22596 7481 22624
rect 7248 22584 7254 22596
rect 7469 22593 7481 22596
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7668 22556 7696 22587
rect 9398 22584 9404 22636
rect 9456 22624 9462 22636
rect 9677 22627 9735 22633
rect 9677 22624 9689 22627
rect 9456 22596 9689 22624
rect 9456 22584 9462 22596
rect 9677 22593 9689 22596
rect 9723 22624 9735 22627
rect 9723 22596 10732 22624
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 7432 22528 7696 22556
rect 10704 22556 10732 22596
rect 11698 22584 11704 22636
rect 11756 22624 11762 22636
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 11756 22596 11897 22624
rect 11756 22584 11762 22596
rect 11885 22593 11897 22596
rect 11931 22624 11943 22627
rect 12066 22624 12072 22636
rect 11931 22596 12072 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 12158 22584 12164 22636
rect 12216 22584 12222 22636
rect 12894 22584 12900 22636
rect 12952 22584 12958 22636
rect 13164 22627 13222 22633
rect 13164 22593 13176 22627
rect 13210 22624 13222 22627
rect 13832 22624 13860 22732
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18782 22760 18788 22772
rect 18012 22732 18788 22760
rect 18012 22720 18018 22732
rect 18782 22720 18788 22732
rect 18840 22760 18846 22772
rect 21361 22763 21419 22769
rect 21361 22760 21373 22763
rect 18840 22732 21373 22760
rect 18840 22720 18846 22732
rect 21361 22729 21373 22732
rect 21407 22729 21419 22763
rect 21361 22723 21419 22729
rect 20714 22692 20720 22704
rect 19996 22664 20720 22692
rect 19996 22633 20024 22664
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 22020 22664 23888 22692
rect 13210 22596 13860 22624
rect 19981 22627 20039 22633
rect 13210 22593 13222 22596
rect 13164 22587 13222 22593
rect 19981 22593 19993 22627
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 20070 22584 20076 22636
rect 20128 22624 20134 22636
rect 20237 22627 20295 22633
rect 20237 22624 20249 22627
rect 20128 22596 20249 22624
rect 20128 22584 20134 22596
rect 20237 22593 20249 22596
rect 20283 22593 20295 22627
rect 20237 22587 20295 22593
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 22020 22633 22048 22664
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21692 22596 22017 22624
rect 21692 22584 21698 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22272 22627 22330 22633
rect 22272 22593 22284 22627
rect 22318 22624 22330 22627
rect 23382 22624 23388 22636
rect 22318 22596 23388 22624
rect 22318 22593 22330 22596
rect 22272 22587 22330 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 23860 22633 23888 22664
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 24118 22701 24124 22704
rect 24112 22692 24124 22701
rect 23992 22664 24124 22692
rect 23992 22652 23998 22664
rect 24112 22655 24124 22664
rect 24118 22652 24124 22655
rect 24176 22652 24182 22704
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22624 23903 22627
rect 24578 22624 24584 22636
rect 23891 22596 24584 22624
rect 23891 22593 23903 22596
rect 23845 22587 23903 22593
rect 24578 22584 24584 22596
rect 24636 22584 24642 22636
rect 10704 22528 12434 22556
rect 7432 22516 7438 22528
rect 11057 22491 11115 22497
rect 11057 22457 11069 22491
rect 11103 22488 11115 22491
rect 12406 22488 12434 22528
rect 12912 22488 12940 22584
rect 11103 22460 11836 22488
rect 12406 22460 12940 22488
rect 11103 22457 11115 22460
rect 11057 22451 11115 22457
rect 11698 22420 11704 22432
rect 6748 22392 11704 22420
rect 6549 22383 6607 22389
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 11808 22420 11836 22460
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 13964 22460 14320 22488
rect 13964 22448 13970 22460
rect 14090 22420 14096 22432
rect 11808 22392 14096 22420
rect 14090 22380 14096 22392
rect 14148 22380 14154 22432
rect 14292 22429 14320 22460
rect 14277 22423 14335 22429
rect 14277 22389 14289 22423
rect 14323 22420 14335 22423
rect 15746 22420 15752 22432
rect 14323 22392 15752 22420
rect 14323 22389 14335 22392
rect 14277 22383 14335 22389
rect 15746 22380 15752 22392
rect 15804 22380 15810 22432
rect 20622 22380 20628 22432
rect 20680 22420 20686 22432
rect 23385 22423 23443 22429
rect 23385 22420 23397 22423
rect 20680 22392 23397 22420
rect 20680 22380 20686 22392
rect 23385 22389 23397 22392
rect 23431 22389 23443 22423
rect 23385 22383 23443 22389
rect 25130 22380 25136 22432
rect 25188 22420 25194 22432
rect 25225 22423 25283 22429
rect 25225 22420 25237 22423
rect 25188 22392 25237 22420
rect 25188 22380 25194 22392
rect 25225 22389 25237 22392
rect 25271 22389 25283 22423
rect 25225 22383 25283 22389
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 7006 22176 7012 22228
rect 7064 22216 7070 22228
rect 7561 22219 7619 22225
rect 7561 22216 7573 22219
rect 7064 22188 7573 22216
rect 7064 22176 7070 22188
rect 7561 22185 7573 22188
rect 7607 22185 7619 22219
rect 7561 22179 7619 22185
rect 10870 22176 10876 22228
rect 10928 22216 10934 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10928 22188 10977 22216
rect 10928 22176 10934 22188
rect 10965 22185 10977 22188
rect 11011 22216 11023 22219
rect 11238 22216 11244 22228
rect 11011 22188 11244 22216
rect 11011 22185 11023 22188
rect 10965 22179 11023 22185
rect 11238 22176 11244 22188
rect 11296 22176 11302 22228
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 10042 22148 10048 22160
rect 9824 22120 10048 22148
rect 9824 22108 9830 22120
rect 10042 22108 10048 22120
rect 10100 22108 10106 22160
rect 10410 22108 10416 22160
rect 10468 22148 10474 22160
rect 10597 22151 10655 22157
rect 10597 22148 10609 22151
rect 10468 22120 10609 22148
rect 10468 22108 10474 22120
rect 10597 22117 10609 22120
rect 10643 22117 10655 22151
rect 10597 22111 10655 22117
rect 1946 22040 1952 22092
rect 2004 22040 2010 22092
rect 5074 22040 5080 22092
rect 5132 22080 5138 22092
rect 6089 22083 6147 22089
rect 6089 22080 6101 22083
rect 5132 22052 6101 22080
rect 5132 22040 5138 22052
rect 6089 22049 6101 22052
rect 6135 22049 6147 22083
rect 6089 22043 6147 22049
rect 7282 22040 7288 22092
rect 7340 22040 7346 22092
rect 7374 22040 7380 22092
rect 7432 22080 7438 22092
rect 8570 22080 8576 22092
rect 7432 22052 8576 22080
rect 7432 22040 7438 22052
rect 8570 22040 8576 22052
rect 8628 22080 8634 22092
rect 9950 22080 9956 22092
rect 8628 22052 9956 22080
rect 8628 22040 8634 22052
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12802 22080 12808 22092
rect 12115 22052 12808 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 24578 22040 24584 22092
rect 24636 22040 24642 22092
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 1673 21975 1731 21981
rect 1688 21944 1716 21975
rect 1854 21972 1860 22024
rect 1912 21972 1918 22024
rect 2130 21972 2136 22024
rect 2188 21972 2194 22024
rect 2314 21972 2320 22024
rect 2372 21972 2378 22024
rect 4062 22012 4068 22024
rect 2700 21984 4068 22012
rect 2700 21944 2728 21984
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 5169 22015 5227 22021
rect 5169 21981 5181 22015
rect 5215 22012 5227 22015
rect 5718 22012 5724 22024
rect 5215 21984 5724 22012
rect 5215 21981 5227 21984
rect 5169 21975 5227 21981
rect 5718 21972 5724 21984
rect 5776 21972 5782 22024
rect 6362 21972 6368 22024
rect 6420 21972 6426 22024
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6730 21972 6736 22024
rect 6788 21972 6794 22024
rect 7300 22012 7328 22040
rect 7300 21984 7420 22012
rect 1688 21916 2728 21944
rect 3878 21904 3884 21956
rect 3936 21944 3942 21956
rect 4985 21947 5043 21953
rect 4985 21944 4997 21947
rect 3936 21916 4997 21944
rect 3936 21904 3942 21916
rect 4985 21913 4997 21916
rect 5031 21913 5043 21947
rect 4985 21907 5043 21913
rect 5537 21947 5595 21953
rect 5537 21913 5549 21947
rect 5583 21944 5595 21947
rect 6914 21944 6920 21956
rect 5583 21916 6920 21944
rect 5583 21913 5595 21916
rect 5537 21907 5595 21913
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 7193 21947 7251 21953
rect 7193 21913 7205 21947
rect 7239 21944 7251 21947
rect 7282 21944 7288 21956
rect 7239 21916 7288 21944
rect 7239 21913 7251 21916
rect 7193 21907 7251 21913
rect 7282 21904 7288 21916
rect 7340 21904 7346 21956
rect 7392 21953 7420 21984
rect 7377 21947 7435 21953
rect 7377 21913 7389 21947
rect 7423 21944 7435 21947
rect 7466 21944 7472 21956
rect 7423 21916 7472 21944
rect 7423 21913 7435 21916
rect 7377 21907 7435 21913
rect 7466 21904 7472 21916
rect 7524 21904 7530 21956
rect 9968 21944 9996 22040
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 10965 21947 11023 21953
rect 10965 21944 10977 21947
rect 7852 21916 9260 21944
rect 9968 21916 10977 21944
rect 7852 21888 7880 21916
rect 5258 21836 5264 21888
rect 5316 21836 5322 21888
rect 5350 21836 5356 21888
rect 5408 21836 5414 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7834 21876 7840 21888
rect 7064 21848 7840 21876
rect 7064 21836 7070 21848
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9122 21876 9128 21888
rect 8904 21848 9128 21876
rect 8904 21836 8910 21848
rect 9122 21836 9128 21848
rect 9180 21836 9186 21888
rect 9232 21876 9260 21916
rect 10965 21913 10977 21916
rect 11011 21913 11023 21947
rect 10965 21907 11023 21913
rect 11072 21916 11284 21944
rect 11072 21876 11100 21916
rect 9232 21848 11100 21876
rect 11146 21836 11152 21888
rect 11204 21836 11210 21888
rect 11256 21876 11284 21916
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 12360 21944 12388 21975
rect 15654 21972 15660 22024
rect 15712 21972 15718 22024
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 18230 22012 18236 22024
rect 16439 21984 18236 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 12124 21916 12388 21944
rect 12124 21904 12130 21916
rect 12434 21876 12440 21888
rect 11256 21848 12440 21876
rect 12434 21836 12440 21848
rect 12492 21876 12498 21888
rect 14182 21876 14188 21888
rect 12492 21848 14188 21876
rect 12492 21836 12498 21848
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 15841 21879 15899 21885
rect 15841 21845 15853 21879
rect 15887 21876 15899 21879
rect 16408 21876 16436 21975
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 21545 22015 21603 22021
rect 21545 21981 21557 22015
rect 21591 22012 21603 22015
rect 21634 22012 21640 22024
rect 21591 21984 21640 22012
rect 21591 21981 21603 21984
rect 21545 21975 21603 21981
rect 21634 21972 21640 21984
rect 21692 21972 21698 22024
rect 25958 21972 25964 22024
rect 26016 22012 26022 22024
rect 26973 22015 27031 22021
rect 26973 22012 26985 22015
rect 26016 21984 26985 22012
rect 26016 21972 26022 21984
rect 26973 21981 26985 21984
rect 27019 21981 27031 22015
rect 26973 21975 27031 21981
rect 16660 21947 16718 21953
rect 16660 21913 16672 21947
rect 16706 21944 16718 21947
rect 18138 21944 18144 21956
rect 16706 21916 18144 21944
rect 16706 21913 16718 21916
rect 16660 21907 16718 21913
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 21790 21947 21848 21953
rect 21790 21944 21802 21947
rect 21560 21916 21802 21944
rect 21560 21888 21588 21916
rect 21790 21913 21802 21916
rect 21836 21913 21848 21947
rect 21790 21907 21848 21913
rect 24486 21904 24492 21956
rect 24544 21944 24550 21956
rect 24826 21947 24884 21953
rect 24826 21944 24838 21947
rect 24544 21916 24838 21944
rect 24544 21904 24550 21916
rect 24826 21913 24838 21916
rect 24872 21944 24884 21947
rect 25130 21944 25136 21956
rect 24872 21916 25136 21944
rect 24872 21913 24884 21916
rect 24826 21907 24884 21913
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 26878 21904 26884 21956
rect 26936 21944 26942 21956
rect 27218 21947 27276 21953
rect 27218 21944 27230 21947
rect 26936 21916 27230 21944
rect 26936 21904 26942 21916
rect 27218 21913 27230 21916
rect 27264 21944 27276 21947
rect 27522 21944 27528 21956
rect 27264 21916 27528 21944
rect 27264 21913 27276 21916
rect 27218 21907 27276 21913
rect 27522 21904 27528 21916
rect 27580 21904 27586 21956
rect 15887 21848 16436 21876
rect 15887 21845 15899 21848
rect 15841 21839 15899 21845
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 20162 21876 20168 21888
rect 17828 21848 20168 21876
rect 17828 21836 17834 21848
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 21542 21836 21548 21888
rect 21600 21836 21606 21888
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22925 21879 22983 21885
rect 22925 21876 22937 21879
rect 22336 21848 22937 21876
rect 22336 21836 22342 21848
rect 22925 21845 22937 21848
rect 22971 21845 22983 21879
rect 22925 21839 22983 21845
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 25961 21879 26019 21885
rect 25961 21876 25973 21879
rect 23348 21848 25973 21876
rect 23348 21836 23354 21848
rect 25961 21845 25973 21848
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26142 21836 26148 21888
rect 26200 21876 26206 21888
rect 28353 21879 28411 21885
rect 28353 21876 28365 21879
rect 26200 21848 28365 21876
rect 26200 21836 26206 21848
rect 28353 21845 28365 21848
rect 28399 21845 28411 21879
rect 28353 21839 28411 21845
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 2314 21632 2320 21684
rect 2372 21672 2378 21684
rect 4065 21675 4123 21681
rect 4065 21672 4077 21675
rect 2372 21644 4077 21672
rect 2372 21632 2378 21644
rect 4065 21641 4077 21644
rect 4111 21641 4123 21675
rect 4065 21635 4123 21641
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 7193 21675 7251 21681
rect 7193 21672 7205 21675
rect 6604 21644 7205 21672
rect 6604 21632 6610 21644
rect 7193 21641 7205 21644
rect 7239 21641 7251 21675
rect 7193 21635 7251 21641
rect 9033 21675 9091 21681
rect 9033 21641 9045 21675
rect 9079 21672 9091 21675
rect 13630 21672 13636 21684
rect 9079 21644 13636 21672
rect 9079 21641 9091 21644
rect 9033 21635 9091 21641
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 17770 21672 17776 21684
rect 13924 21644 17776 21672
rect 2130 21564 2136 21616
rect 2188 21604 2194 21616
rect 7920 21607 7978 21613
rect 2188 21576 7236 21604
rect 2188 21564 2194 21576
rect 7208 21548 7236 21576
rect 7920 21573 7932 21607
rect 7966 21604 7978 21607
rect 12428 21607 12486 21613
rect 7966 21576 11836 21604
rect 7966 21573 7978 21576
rect 7920 21567 7978 21573
rect 3142 21496 3148 21548
rect 3200 21496 3206 21548
rect 3973 21539 4031 21545
rect 3973 21505 3985 21539
rect 4019 21536 4031 21539
rect 4338 21536 4344 21548
rect 4019 21508 4344 21536
rect 4019 21505 4031 21508
rect 3973 21499 4031 21505
rect 4338 21496 4344 21508
rect 4396 21496 4402 21548
rect 5810 21496 5816 21548
rect 5868 21536 5874 21548
rect 6638 21536 6644 21548
rect 5868 21508 6644 21536
rect 5868 21496 5874 21508
rect 6638 21496 6644 21508
rect 6696 21536 6702 21548
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6696 21508 6837 21536
rect 6696 21496 6702 21508
rect 6825 21505 6837 21508
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 7098 21536 7104 21548
rect 7055 21508 7104 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21536 7711 21539
rect 7699 21508 9168 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 3329 21403 3387 21409
rect 3329 21369 3341 21403
rect 3375 21400 3387 21403
rect 5258 21400 5264 21412
rect 3375 21372 5264 21400
rect 3375 21369 3387 21372
rect 3329 21363 3387 21369
rect 5258 21360 5264 21372
rect 5316 21360 5322 21412
rect 9140 21400 9168 21508
rect 9232 21480 9260 21576
rect 9760 21539 9818 21545
rect 9760 21505 9772 21539
rect 9806 21536 9818 21539
rect 11698 21536 11704 21548
rect 9806 21508 11704 21536
rect 9806 21505 9818 21508
rect 9760 21499 9818 21505
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 9214 21428 9220 21480
rect 9272 21428 9278 21480
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 9493 21471 9551 21477
rect 9493 21468 9505 21471
rect 9456 21440 9505 21468
rect 9456 21428 9462 21440
rect 9493 21437 9505 21440
rect 9539 21437 9551 21471
rect 9493 21431 9551 21437
rect 9416 21400 9444 21428
rect 9140 21372 9444 21400
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 9490 21332 9496 21344
rect 7156 21304 9496 21332
rect 7156 21292 7162 21304
rect 9490 21292 9496 21304
rect 9548 21292 9554 21344
rect 10594 21292 10600 21344
rect 10652 21332 10658 21344
rect 10873 21335 10931 21341
rect 10873 21332 10885 21335
rect 10652 21304 10885 21332
rect 10652 21292 10658 21304
rect 10873 21301 10885 21304
rect 10919 21301 10931 21335
rect 11808 21332 11836 21576
rect 12428 21573 12440 21607
rect 12474 21604 12486 21607
rect 13924 21604 13952 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 18500 21607 18558 21613
rect 12474 21576 13952 21604
rect 14016 21576 16252 21604
rect 12474 21573 12486 21576
rect 12428 21567 12486 21573
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12250 21536 12256 21548
rect 12207 21508 12256 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 14016 21545 14044 21576
rect 16224 21548 16252 21576
rect 18500 21573 18512 21607
rect 18546 21604 18558 21607
rect 18690 21604 18696 21616
rect 18546 21576 18696 21604
rect 18546 21573 18558 21576
rect 18500 21567 18558 21573
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 20530 21604 20536 21616
rect 18800 21576 20536 21604
rect 14001 21539 14059 21545
rect 14001 21505 14013 21539
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 15562 21496 15568 21548
rect 15620 21496 15626 21548
rect 15930 21496 15936 21548
rect 15988 21496 15994 21548
rect 16206 21496 16212 21548
rect 16264 21496 16270 21548
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18800 21536 18828 21576
rect 20530 21564 20536 21576
rect 20588 21604 20594 21616
rect 21450 21604 21456 21616
rect 20588 21576 21456 21604
rect 20588 21564 20594 21576
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 23106 21564 23112 21616
rect 23164 21604 23170 21616
rect 25958 21604 25964 21616
rect 23164 21576 23612 21604
rect 23164 21564 23170 21576
rect 20346 21545 20352 21548
rect 20340 21536 20352 21545
rect 18340 21508 18828 21536
rect 20307 21508 20352 21536
rect 15838 21428 15844 21480
rect 15896 21428 15902 21480
rect 18340 21468 18368 21508
rect 20340 21499 20352 21508
rect 20404 21536 20410 21548
rect 23290 21536 23296 21548
rect 20404 21508 23296 21536
rect 20346 21496 20352 21499
rect 20404 21496 20410 21508
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 23474 21545 23480 21548
rect 23468 21536 23480 21545
rect 23435 21508 23480 21536
rect 23468 21499 23480 21508
rect 23474 21496 23480 21499
rect 23532 21496 23538 21548
rect 23584 21536 23612 21576
rect 25240 21576 25964 21604
rect 25240 21545 25268 21576
rect 25958 21564 25964 21576
rect 26016 21564 26022 21616
rect 25225 21539 25283 21545
rect 23584 21508 25176 21536
rect 15948 21440 18368 21468
rect 15286 21360 15292 21412
rect 15344 21400 15350 21412
rect 15654 21400 15660 21412
rect 15344 21372 15660 21400
rect 15344 21360 15350 21372
rect 15654 21360 15660 21372
rect 15712 21400 15718 21412
rect 15948 21400 15976 21440
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 19392 21440 20085 21468
rect 19392 21428 19398 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 23198 21428 23204 21480
rect 23256 21428 23262 21480
rect 25148 21468 25176 21508
rect 25225 21505 25237 21539
rect 25271 21505 25283 21539
rect 25481 21539 25539 21545
rect 25481 21536 25493 21539
rect 25225 21499 25283 21505
rect 25332 21508 25493 21536
rect 25332 21468 25360 21508
rect 25481 21505 25493 21508
rect 25527 21505 25539 21539
rect 25481 21499 25539 21505
rect 25148 21440 25360 21468
rect 15712 21372 15976 21400
rect 15712 21360 15718 21372
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 11808 21304 13553 21332
rect 10873 21295 10931 21301
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 13541 21295 13599 21301
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 19300 21304 19625 21332
rect 19300 21292 19306 21304
rect 19613 21301 19625 21304
rect 19659 21301 19671 21335
rect 19613 21295 19671 21301
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20070 21332 20076 21344
rect 19852 21304 20076 21332
rect 19852 21292 19858 21304
rect 20070 21292 20076 21304
rect 20128 21332 20134 21344
rect 21453 21335 21511 21341
rect 21453 21332 21465 21335
rect 20128 21304 21465 21332
rect 20128 21292 20134 21304
rect 21453 21301 21465 21304
rect 21499 21301 21511 21335
rect 21453 21295 21511 21301
rect 22738 21292 22744 21344
rect 22796 21332 22802 21344
rect 24581 21335 24639 21341
rect 24581 21332 24593 21335
rect 22796 21304 24593 21332
rect 22796 21292 22802 21304
rect 24581 21301 24593 21304
rect 24627 21301 24639 21335
rect 24581 21295 24639 21301
rect 24854 21292 24860 21344
rect 24912 21332 24918 21344
rect 25590 21332 25596 21344
rect 24912 21304 25596 21332
rect 24912 21292 24918 21304
rect 25590 21292 25596 21304
rect 25648 21332 25654 21344
rect 26605 21335 26663 21341
rect 26605 21332 26617 21335
rect 25648 21304 26617 21332
rect 25648 21292 25654 21304
rect 26605 21301 26617 21304
rect 26651 21301 26663 21335
rect 26605 21295 26663 21301
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 6457 21131 6515 21137
rect 6457 21097 6469 21131
rect 6503 21128 6515 21131
rect 6914 21128 6920 21140
rect 6503 21100 6920 21128
rect 6503 21097 6515 21100
rect 6457 21091 6515 21097
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 7190 21088 7196 21140
rect 7248 21128 7254 21140
rect 10226 21128 10232 21140
rect 7248 21100 10232 21128
rect 7248 21088 7254 21100
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 12342 21128 12348 21140
rect 11112 21100 12348 21128
rect 11112 21088 11118 21100
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 16482 21128 16488 21140
rect 12728 21100 16488 21128
rect 12728 21069 12756 21100
rect 7101 21063 7159 21069
rect 7101 21029 7113 21063
rect 7147 21029 7159 21063
rect 7101 21023 7159 21029
rect 12713 21063 12771 21069
rect 12713 21029 12725 21063
rect 12759 21029 12771 21063
rect 12713 21023 12771 21029
rect 7116 20992 7144 21023
rect 5184 20964 7144 20992
rect 7392 20964 11468 20992
rect 4890 20884 4896 20936
rect 4948 20884 4954 20936
rect 5184 20933 5212 20964
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20893 5227 20927
rect 5169 20887 5227 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 7282 20924 7288 20936
rect 5399 20896 5488 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 1486 20748 1492 20800
rect 1544 20788 1550 20800
rect 5077 20791 5135 20797
rect 5077 20788 5089 20791
rect 1544 20760 5089 20788
rect 1544 20748 1550 20760
rect 5077 20757 5089 20760
rect 5123 20757 5135 20791
rect 5077 20751 5135 20757
rect 5350 20748 5356 20800
rect 5408 20788 5414 20800
rect 5460 20788 5488 20896
rect 7024 20896 7288 20924
rect 6270 20816 6276 20868
rect 6328 20816 6334 20868
rect 6489 20859 6547 20865
rect 6489 20825 6501 20859
rect 6535 20856 6547 20859
rect 7024 20856 7052 20896
rect 7282 20884 7288 20896
rect 7340 20924 7346 20936
rect 7392 20933 7420 20964
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 7340 20896 7389 20924
rect 7340 20884 7346 20896
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 9306 20924 9312 20936
rect 8619 20896 9312 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 9306 20884 9312 20896
rect 9364 20924 9370 20936
rect 9364 20896 10088 20924
rect 9364 20884 9370 20896
rect 6535 20828 7052 20856
rect 7101 20859 7159 20865
rect 6535 20825 6547 20828
rect 6489 20819 6547 20825
rect 7101 20825 7113 20859
rect 7147 20825 7159 20859
rect 7101 20819 7159 20825
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 5408 20760 6653 20788
rect 5408 20748 5414 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 6914 20748 6920 20800
rect 6972 20788 6978 20800
rect 7116 20788 7144 20819
rect 7190 20816 7196 20868
rect 7248 20856 7254 20868
rect 8205 20859 8263 20865
rect 8205 20856 8217 20859
rect 7248 20828 8217 20856
rect 7248 20816 7254 20828
rect 8205 20825 8217 20828
rect 8251 20825 8263 20859
rect 8205 20819 8263 20825
rect 9582 20816 9588 20868
rect 9640 20816 9646 20868
rect 9766 20816 9772 20868
rect 9824 20816 9830 20868
rect 6972 20760 7144 20788
rect 6972 20748 6978 20760
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 7466 20788 7472 20800
rect 7340 20760 7472 20788
rect 7340 20748 7346 20760
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 9950 20748 9956 20800
rect 10008 20748 10014 20800
rect 10060 20788 10088 20896
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11333 20927 11391 20933
rect 11333 20924 11345 20927
rect 11204 20896 11345 20924
rect 11204 20884 11210 20896
rect 11333 20893 11345 20896
rect 11379 20893 11391 20927
rect 11440 20924 11468 20964
rect 12986 20924 12992 20936
rect 11440 20896 12992 20924
rect 11333 20887 11391 20893
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 11606 20865 11612 20868
rect 11600 20856 11612 20865
rect 11567 20828 11612 20856
rect 11600 20819 11612 20828
rect 11606 20816 11612 20819
rect 11664 20816 11670 20868
rect 11698 20816 11704 20868
rect 11756 20856 11762 20868
rect 13096 20856 13124 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 22738 21128 22744 21140
rect 22066 21100 22744 21128
rect 14182 20952 14188 21004
rect 14240 20992 14246 21004
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 14240 20964 14289 20992
rect 14240 20952 14246 20964
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20924 14519 20927
rect 15473 20927 15531 20933
rect 14507 20896 15148 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 11756 20828 13124 20856
rect 11756 20816 11762 20828
rect 11790 20788 11796 20800
rect 10060 20760 11796 20788
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 13872 20760 14657 20788
rect 13872 20748 13878 20760
rect 14645 20757 14657 20760
rect 14691 20757 14703 20791
rect 15120 20788 15148 20896
rect 15473 20893 15485 20927
rect 15519 20924 15531 20927
rect 16758 20924 16764 20936
rect 15519 20896 16764 20924
rect 15519 20893 15531 20896
rect 15473 20887 15531 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 20625 20927 20683 20933
rect 20625 20924 20637 20927
rect 19392 20896 20637 20924
rect 19392 20884 19398 20896
rect 20625 20893 20637 20896
rect 20671 20924 20683 20927
rect 20714 20924 20720 20936
rect 20671 20896 20720 20924
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 20892 20927 20950 20933
rect 20892 20893 20904 20927
rect 20938 20924 20950 20927
rect 22066 20924 22094 21100
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 20938 20896 22094 20924
rect 22465 20927 22523 20933
rect 20938 20893 20950 20896
rect 20892 20887 20950 20893
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 23198 20924 23204 20936
rect 22511 20896 23204 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 25958 20884 25964 20936
rect 26016 20924 26022 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 26016 20896 26065 20924
rect 26016 20884 26022 20896
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 15562 20816 15568 20868
rect 15620 20856 15626 20868
rect 15718 20859 15776 20865
rect 15718 20856 15730 20859
rect 15620 20828 15730 20856
rect 15620 20816 15626 20828
rect 15718 20825 15730 20828
rect 15764 20825 15776 20859
rect 15718 20819 15776 20825
rect 22370 20816 22376 20868
rect 22428 20856 22434 20868
rect 22710 20859 22768 20865
rect 22710 20856 22722 20859
rect 22428 20828 22722 20856
rect 22428 20816 22434 20828
rect 22710 20825 22722 20828
rect 22756 20825 22768 20859
rect 22710 20819 22768 20825
rect 25130 20816 25136 20868
rect 25188 20856 25194 20868
rect 26298 20859 26356 20865
rect 26298 20856 26310 20859
rect 25188 20828 26310 20856
rect 25188 20816 25194 20828
rect 26298 20825 26310 20828
rect 26344 20825 26356 20859
rect 26298 20819 26356 20825
rect 16206 20788 16212 20800
rect 15120 20760 16212 20788
rect 14645 20751 14703 20757
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 16853 20791 16911 20797
rect 16853 20757 16865 20791
rect 16899 20788 16911 20791
rect 18046 20788 18052 20800
rect 16899 20760 18052 20788
rect 16899 20757 16911 20760
rect 16853 20751 16911 20757
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 21634 20748 21640 20800
rect 21692 20788 21698 20800
rect 22005 20791 22063 20797
rect 22005 20788 22017 20791
rect 21692 20760 22017 20788
rect 21692 20748 21698 20760
rect 22005 20757 22017 20760
rect 22051 20757 22063 20791
rect 22005 20751 22063 20757
rect 23842 20748 23848 20800
rect 23900 20748 23906 20800
rect 26510 20748 26516 20800
rect 26568 20788 26574 20800
rect 27433 20791 27491 20797
rect 27433 20788 27445 20791
rect 26568 20760 27445 20788
rect 26568 20748 26574 20760
rect 27433 20757 27445 20760
rect 27479 20757 27491 20791
rect 27433 20751 27491 20757
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 5166 20584 5172 20596
rect 4304 20556 5172 20584
rect 4304 20544 4310 20556
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 5353 20587 5411 20593
rect 5353 20553 5365 20587
rect 5399 20584 5411 20587
rect 5442 20584 5448 20596
rect 5399 20556 5448 20584
rect 5399 20553 5411 20556
rect 5353 20547 5411 20553
rect 5442 20544 5448 20556
rect 5500 20544 5506 20596
rect 5721 20587 5779 20593
rect 5721 20553 5733 20587
rect 5767 20584 5779 20587
rect 6270 20584 6276 20596
rect 5767 20556 6276 20584
rect 5767 20553 5779 20556
rect 5721 20547 5779 20553
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6880 20556 7021 20584
rect 6880 20544 6886 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 7377 20587 7435 20593
rect 7377 20553 7389 20587
rect 7423 20584 7435 20587
rect 10318 20584 10324 20596
rect 7423 20556 10324 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 10502 20544 10508 20596
rect 10560 20544 10566 20596
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20584 11759 20587
rect 12158 20584 12164 20596
rect 11747 20556 12164 20584
rect 11747 20553 11759 20556
rect 11701 20547 11759 20553
rect 12158 20544 12164 20556
rect 12216 20544 12222 20596
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 3234 20476 3240 20528
rect 3292 20516 3298 20528
rect 8110 20516 8116 20528
rect 3292 20488 5580 20516
rect 3292 20476 3298 20488
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20448 4215 20451
rect 4982 20448 4988 20460
rect 4203 20420 4988 20448
rect 4203 20417 4215 20420
rect 4157 20411 4215 20417
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 5552 20457 5580 20488
rect 7392 20488 8116 20516
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 4246 20340 4252 20392
rect 4304 20340 4310 20392
rect 4798 20340 4804 20392
rect 4856 20380 4862 20392
rect 5442 20380 5448 20392
rect 4856 20352 5448 20380
rect 4856 20340 4862 20352
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 5828 20380 5856 20411
rect 5902 20408 5908 20460
rect 5960 20448 5966 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 5960 20420 7205 20448
rect 5960 20408 5966 20420
rect 7193 20417 7205 20420
rect 7239 20448 7251 20451
rect 7392 20448 7420 20488
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 8389 20519 8447 20525
rect 8389 20485 8401 20519
rect 8435 20516 8447 20519
rect 9674 20516 9680 20528
rect 8435 20488 9680 20516
rect 8435 20485 8447 20488
rect 8389 20479 8447 20485
rect 9674 20476 9680 20488
rect 9732 20516 9738 20528
rect 10410 20516 10416 20528
rect 9732 20488 10416 20516
rect 9732 20476 9738 20488
rect 10410 20476 10416 20488
rect 10468 20476 10474 20528
rect 11057 20519 11115 20525
rect 11057 20485 11069 20519
rect 11103 20516 11115 20519
rect 12710 20516 12716 20528
rect 11103 20488 12716 20516
rect 11103 20485 11115 20488
rect 11057 20479 11115 20485
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 14338 20519 14396 20525
rect 14338 20516 14350 20519
rect 13964 20488 14350 20516
rect 13964 20476 13970 20488
rect 14338 20485 14350 20488
rect 14384 20485 14396 20519
rect 19334 20516 19340 20528
rect 14338 20479 14396 20485
rect 18156 20488 19340 20516
rect 7239 20420 7420 20448
rect 7239 20417 7251 20420
rect 7193 20411 7251 20417
rect 7466 20408 7472 20460
rect 7524 20408 7530 20460
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9306 20448 9312 20460
rect 9263 20420 9312 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 6270 20380 6276 20392
rect 5828 20352 6276 20380
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 8220 20380 8248 20411
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 9490 20408 9496 20460
rect 9548 20408 9554 20460
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 14182 20448 14188 20460
rect 10827 20420 14188 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15620 20420 15945 20448
rect 15620 20408 15626 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 7156 20352 9444 20380
rect 7156 20340 7162 20352
rect 4525 20315 4583 20321
rect 4525 20281 4537 20315
rect 4571 20312 4583 20315
rect 6730 20312 6736 20324
rect 4571 20284 6736 20312
rect 4571 20281 4583 20284
rect 4525 20275 4583 20281
rect 6730 20272 6736 20284
rect 6788 20272 6794 20324
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 9033 20315 9091 20321
rect 9033 20312 9045 20315
rect 7800 20284 9045 20312
rect 7800 20272 7806 20284
rect 9033 20281 9045 20284
rect 9079 20281 9091 20315
rect 9033 20275 9091 20281
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 4798 20244 4804 20256
rect 4387 20216 4804 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 8570 20204 8576 20256
rect 8628 20204 8634 20256
rect 9416 20253 9444 20352
rect 9508 20312 9536 20408
rect 10502 20340 10508 20392
rect 10560 20380 10566 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10560 20352 10701 20380
rect 10560 20340 10566 20352
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11149 20383 11207 20389
rect 11149 20380 11161 20383
rect 11112 20352 11161 20380
rect 11112 20340 11118 20352
rect 11149 20349 11161 20352
rect 11195 20349 11207 20383
rect 11149 20343 11207 20349
rect 11606 20340 11612 20392
rect 11664 20380 11670 20392
rect 11885 20383 11943 20389
rect 11885 20380 11897 20383
rect 11664 20352 11897 20380
rect 11664 20340 11670 20352
rect 11885 20349 11897 20352
rect 11931 20349 11943 20383
rect 11885 20343 11943 20349
rect 11974 20340 11980 20392
rect 12032 20340 12038 20392
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20349 12127 20383
rect 12069 20343 12127 20349
rect 9508 20284 10548 20312
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 9582 20244 9588 20256
rect 9447 20216 9588 20244
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 9582 20204 9588 20216
rect 9640 20244 9646 20256
rect 10410 20244 10416 20256
rect 9640 20216 10416 20244
rect 9640 20204 9646 20216
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10520 20244 10548 20284
rect 10870 20272 10876 20324
rect 10928 20312 10934 20324
rect 12084 20312 12112 20343
rect 12158 20340 12164 20392
rect 12216 20340 12222 20392
rect 12250 20340 12256 20392
rect 12308 20380 12314 20392
rect 14093 20383 14151 20389
rect 14093 20380 14105 20383
rect 12308 20352 14105 20380
rect 12308 20340 12314 20352
rect 14093 20349 14105 20352
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 15654 20340 15660 20392
rect 15712 20380 15718 20392
rect 16224 20380 16252 20411
rect 15712 20352 16252 20380
rect 15712 20340 15718 20352
rect 16758 20340 16764 20392
rect 16816 20380 16822 20392
rect 18156 20389 18184 20488
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 21634 20516 21640 20528
rect 19812 20488 21640 20516
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 18397 20451 18455 20457
rect 18397 20448 18409 20451
rect 18288 20420 18409 20448
rect 18288 20408 18294 20420
rect 18397 20417 18409 20420
rect 18443 20448 18455 20451
rect 19812 20448 19840 20488
rect 21634 20476 21640 20488
rect 21692 20476 21698 20528
rect 23198 20516 23204 20528
rect 22020 20488 23204 20516
rect 18443 20420 19840 20448
rect 18443 20417 18455 20420
rect 18397 20411 18455 20417
rect 19886 20408 19892 20460
rect 19944 20448 19950 20460
rect 22020 20457 22048 20488
rect 23198 20476 23204 20488
rect 23256 20516 23262 20528
rect 25958 20516 25964 20528
rect 23256 20488 25964 20516
rect 23256 20476 23262 20488
rect 22278 20457 22284 20460
rect 20237 20451 20295 20457
rect 20237 20448 20249 20451
rect 19944 20420 20249 20448
rect 19944 20408 19950 20420
rect 20237 20417 20249 20420
rect 20283 20417 20295 20451
rect 20237 20411 20295 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22272 20448 22284 20457
rect 22239 20420 22284 20448
rect 22005 20411 22063 20417
rect 22272 20411 22284 20420
rect 22278 20408 22284 20411
rect 22336 20408 22342 20460
rect 23860 20457 23888 20488
rect 25958 20476 25964 20488
rect 26016 20476 26022 20528
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 24112 20451 24170 20457
rect 24112 20417 24124 20451
rect 24158 20448 24170 20451
rect 24394 20448 24400 20460
rect 24158 20420 24400 20448
rect 24158 20417 24170 20420
rect 24112 20411 24170 20417
rect 24394 20408 24400 20420
rect 24452 20408 24458 20460
rect 18141 20383 18199 20389
rect 18141 20380 18153 20383
rect 16816 20352 18153 20380
rect 16816 20340 16822 20352
rect 18141 20349 18153 20352
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 19978 20340 19984 20392
rect 20036 20340 20042 20392
rect 10928 20284 12112 20312
rect 10928 20272 10934 20284
rect 15930 20272 15936 20324
rect 15988 20272 15994 20324
rect 23658 20312 23664 20324
rect 22940 20284 23664 20312
rect 11974 20244 11980 20256
rect 10520 20216 11980 20244
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 16448 20216 19533 20244
rect 16448 20204 16454 20216
rect 19521 20213 19533 20216
rect 19567 20213 19579 20247
rect 19521 20207 19579 20213
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 22940 20244 22968 20284
rect 23658 20272 23664 20284
rect 23716 20272 23722 20324
rect 21407 20216 22968 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 23382 20204 23388 20256
rect 23440 20204 23446 20256
rect 25130 20204 25136 20256
rect 25188 20244 25194 20256
rect 25225 20247 25283 20253
rect 25225 20244 25237 20247
rect 25188 20216 25237 20244
rect 25188 20204 25194 20216
rect 25225 20213 25237 20216
rect 25271 20213 25283 20247
rect 25225 20207 25283 20213
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5626 20040 5632 20052
rect 5040 20012 5632 20040
rect 5040 20000 5046 20012
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 5718 20000 5724 20052
rect 5776 20000 5782 20052
rect 6086 20000 6092 20052
rect 6144 20040 6150 20052
rect 6733 20043 6791 20049
rect 6733 20040 6745 20043
rect 6144 20012 6745 20040
rect 6144 20000 6150 20012
rect 6733 20009 6745 20012
rect 6779 20009 6791 20043
rect 6733 20003 6791 20009
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7190 20040 7196 20052
rect 6963 20012 7196 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 8297 20043 8355 20049
rect 8297 20009 8309 20043
rect 8343 20040 8355 20043
rect 8846 20040 8852 20052
rect 8343 20012 8852 20040
rect 8343 20009 8355 20012
rect 8297 20003 8355 20009
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 9858 20040 9864 20052
rect 9732 20012 9864 20040
rect 9732 20000 9738 20012
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 10226 20000 10232 20052
rect 10284 20000 10290 20052
rect 10410 20000 10416 20052
rect 10468 20040 10474 20052
rect 10778 20040 10784 20052
rect 10468 20012 10784 20040
rect 10468 20000 10474 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17402 20040 17408 20052
rect 17184 20012 17408 20040
rect 17184 20000 17190 20012
rect 17402 20000 17408 20012
rect 17460 20040 17466 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 17460 20012 18153 20040
rect 17460 20000 17466 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 18141 20003 18199 20009
rect 22833 20043 22891 20049
rect 22833 20009 22845 20043
rect 22879 20040 22891 20043
rect 23198 20040 23204 20052
rect 22879 20012 23204 20040
rect 22879 20009 22891 20012
rect 22833 20003 22891 20009
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 26605 20043 26663 20049
rect 26605 20040 26617 20043
rect 23532 20012 26617 20040
rect 23532 20000 23538 20012
rect 26605 20009 26617 20012
rect 26651 20009 26663 20043
rect 26605 20003 26663 20009
rect 2222 19932 2228 19984
rect 2280 19972 2286 19984
rect 7650 19972 7656 19984
rect 2280 19944 7656 19972
rect 2280 19932 2286 19944
rect 7650 19932 7656 19944
rect 7708 19932 7714 19984
rect 12434 19972 12440 19984
rect 9600 19944 12440 19972
rect 4172 19876 5028 19904
rect 4172 19845 4200 19876
rect 5000 19845 5028 19876
rect 5166 19864 5172 19916
rect 5224 19904 5230 19916
rect 5224 19876 5488 19904
rect 5224 19864 5230 19876
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19805 4215 19839
rect 4157 19799 4215 19805
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4387 19808 4905 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4893 19805 4905 19808
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19836 5043 19839
rect 5350 19836 5356 19848
rect 5031 19808 5356 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 4908 19768 4936 19799
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 5460 19836 5488 19876
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 5592 19876 5733 19904
rect 5592 19864 5598 19876
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 5460 19808 5580 19836
rect 5552 19768 5580 19808
rect 5626 19796 5632 19848
rect 5684 19796 5690 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 6472 19808 8033 19836
rect 6472 19768 6500 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 9600 19836 9628 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10870 19904 10876 19916
rect 9916 19876 10876 19904
rect 9916 19864 9922 19876
rect 10870 19864 10876 19876
rect 10928 19904 10934 19916
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 10928 19876 11069 19904
rect 10928 19864 10934 19876
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 16758 19864 16764 19916
rect 16816 19864 16822 19916
rect 19978 19864 19984 19916
rect 20036 19904 20042 19916
rect 20036 19876 20944 19904
rect 20036 19864 20042 19876
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9600 19808 9689 19836
rect 8021 19799 8079 19805
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 10045 19839 10103 19845
rect 9677 19799 9735 19805
rect 9784 19808 9996 19836
rect 4908 19740 5304 19768
rect 5552 19740 6500 19768
rect 3326 19660 3332 19712
rect 3384 19700 3390 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 3384 19672 4261 19700
rect 3384 19660 3390 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4249 19663 4307 19669
rect 5166 19660 5172 19712
rect 5224 19660 5230 19712
rect 5276 19700 5304 19740
rect 6546 19728 6552 19780
rect 6604 19728 6610 19780
rect 7098 19768 7104 19780
rect 6656 19740 7104 19768
rect 5626 19700 5632 19712
rect 5276 19672 5632 19700
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 5997 19703 6055 19709
rect 5997 19669 6009 19703
rect 6043 19700 6055 19703
rect 6656 19700 6684 19740
rect 7098 19728 7104 19740
rect 7156 19728 7162 19780
rect 6043 19672 6684 19700
rect 6043 19669 6055 19672
rect 5997 19663 6055 19669
rect 6730 19660 6736 19712
rect 6788 19709 6794 19712
rect 6788 19703 6807 19709
rect 6795 19669 6807 19703
rect 6788 19663 6807 19669
rect 6788 19660 6794 19663
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7834 19700 7840 19712
rect 7248 19672 7840 19700
rect 7248 19660 7254 19672
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 8036 19700 8064 19799
rect 8110 19728 8116 19780
rect 8168 19768 8174 19780
rect 9784 19768 9812 19808
rect 8168 19740 9812 19768
rect 8168 19728 8174 19740
rect 9858 19728 9864 19780
rect 9916 19728 9922 19780
rect 9968 19777 9996 19808
rect 10045 19805 10057 19839
rect 10091 19836 10103 19839
rect 10962 19836 10968 19848
rect 10091 19808 10968 19836
rect 10091 19805 10103 19808
rect 10045 19799 10103 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11238 19796 11244 19848
rect 11296 19796 11302 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 20809 19839 20867 19845
rect 20809 19836 20821 19839
rect 20772 19808 20821 19836
rect 20772 19796 20778 19808
rect 20809 19805 20821 19808
rect 20855 19805 20867 19839
rect 20916 19836 20944 19876
rect 22646 19836 22652 19848
rect 20916 19808 22652 19836
rect 20809 19799 20867 19805
rect 22646 19796 22652 19808
rect 22704 19796 22710 19848
rect 25225 19839 25283 19845
rect 25225 19805 25237 19839
rect 25271 19836 25283 19839
rect 25958 19836 25964 19848
rect 25271 19808 25964 19836
rect 25271 19805 25283 19808
rect 25225 19799 25283 19805
rect 25958 19796 25964 19808
rect 26016 19836 26022 19848
rect 26970 19836 26976 19848
rect 26016 19808 26976 19836
rect 26016 19796 26022 19808
rect 26970 19796 26976 19808
rect 27028 19796 27034 19848
rect 9953 19771 10011 19777
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 10134 19768 10140 19780
rect 9999 19740 10140 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 10134 19728 10140 19740
rect 10192 19728 10198 19780
rect 11422 19728 11428 19780
rect 11480 19728 11486 19780
rect 11514 19728 11520 19780
rect 11572 19768 11578 19780
rect 12342 19768 12348 19780
rect 11572 19740 12348 19768
rect 11572 19728 11578 19740
rect 12342 19728 12348 19740
rect 12400 19768 12406 19780
rect 15562 19768 15568 19780
rect 12400 19740 15568 19768
rect 12400 19728 12406 19740
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 16390 19728 16396 19780
rect 16448 19768 16454 19780
rect 17006 19771 17064 19777
rect 17006 19768 17018 19771
rect 16448 19740 17018 19768
rect 16448 19728 16454 19740
rect 17006 19737 17018 19740
rect 17052 19737 17064 19771
rect 17006 19731 17064 19737
rect 19058 19728 19064 19780
rect 19116 19768 19122 19780
rect 21054 19771 21112 19777
rect 21054 19768 21066 19771
rect 19116 19740 21066 19768
rect 19116 19728 19122 19740
rect 21054 19737 21066 19740
rect 21100 19768 21112 19771
rect 23382 19768 23388 19780
rect 21100 19740 23388 19768
rect 21100 19737 21112 19740
rect 21054 19731 21112 19737
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 25492 19771 25550 19777
rect 25492 19737 25504 19771
rect 25538 19768 25550 19771
rect 25774 19768 25780 19780
rect 25538 19740 25780 19768
rect 25538 19737 25550 19740
rect 25492 19731 25550 19737
rect 25774 19728 25780 19740
rect 25832 19728 25838 19780
rect 10410 19700 10416 19712
rect 8036 19672 10416 19700
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 11330 19660 11336 19712
rect 11388 19660 11394 19712
rect 11609 19703 11667 19709
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 13262 19700 13268 19712
rect 11655 19672 13268 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 13262 19660 13268 19672
rect 13320 19700 13326 19712
rect 15654 19700 15660 19712
rect 13320 19672 15660 19700
rect 13320 19660 13326 19672
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 22186 19660 22192 19712
rect 22244 19660 22250 19712
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 25222 19700 25228 19712
rect 22704 19672 25228 19700
rect 22704 19660 22710 19672
rect 25222 19660 25228 19672
rect 25280 19660 25286 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 3237 19499 3295 19505
rect 3237 19465 3249 19499
rect 3283 19496 3295 19499
rect 3694 19496 3700 19508
rect 3283 19468 3700 19496
rect 3283 19465 3295 19468
rect 3237 19459 3295 19465
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 4632 19468 7604 19496
rect 3970 19388 3976 19440
rect 4028 19428 4034 19440
rect 4632 19428 4660 19468
rect 4028 19400 4660 19428
rect 7193 19431 7251 19437
rect 4028 19388 4034 19400
rect 7193 19397 7205 19431
rect 7239 19428 7251 19431
rect 7374 19428 7380 19440
rect 7239 19400 7380 19428
rect 7239 19397 7251 19400
rect 7193 19391 7251 19397
rect 7374 19388 7380 19400
rect 7432 19388 7438 19440
rect 7576 19428 7604 19468
rect 7650 19456 7656 19508
rect 7708 19496 7714 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7708 19468 8125 19496
rect 7708 19456 7714 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 9861 19499 9919 19505
rect 9861 19465 9873 19499
rect 9907 19496 9919 19499
rect 10042 19496 10048 19508
rect 9907 19468 10048 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10502 19456 10508 19508
rect 10560 19456 10566 19508
rect 10778 19456 10784 19508
rect 10836 19496 10842 19508
rect 13998 19496 14004 19508
rect 10836 19468 11192 19496
rect 10836 19456 10842 19468
rect 9585 19431 9643 19437
rect 9585 19428 9597 19431
rect 7576 19400 9597 19428
rect 9585 19397 9597 19400
rect 9631 19428 9643 19431
rect 10134 19428 10140 19440
rect 9631 19400 10140 19428
rect 9631 19397 9643 19400
rect 9585 19391 9643 19397
rect 10134 19388 10140 19400
rect 10192 19388 10198 19440
rect 11054 19428 11060 19440
rect 10796 19400 11060 19428
rect 3326 19320 3332 19372
rect 3384 19320 3390 19372
rect 3513 19363 3571 19369
rect 3513 19334 3525 19363
rect 3436 19329 3525 19334
rect 3559 19329 3571 19363
rect 3436 19323 3571 19329
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 5166 19360 5172 19372
rect 4387 19332 5172 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 3436 19306 3556 19323
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 7392 19360 7420 19388
rect 7650 19360 7656 19372
rect 6932 19332 7144 19360
rect 7392 19332 7656 19360
rect 3436 19236 3464 19306
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 3418 19184 3424 19236
rect 3476 19224 3482 19236
rect 4632 19224 4660 19255
rect 5074 19252 5080 19304
rect 5132 19292 5138 19304
rect 6638 19292 6644 19304
rect 5132 19264 6644 19292
rect 5132 19252 5138 19264
rect 6638 19252 6644 19264
rect 6696 19292 6702 19304
rect 6932 19292 6960 19332
rect 6696 19264 6960 19292
rect 6696 19252 6702 19264
rect 7006 19252 7012 19304
rect 7064 19252 7070 19304
rect 7116 19292 7144 19332
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8481 19363 8539 19369
rect 8481 19360 8493 19363
rect 8220 19332 8493 19360
rect 8220 19292 8248 19332
rect 8481 19329 8493 19332
rect 8527 19360 8539 19363
rect 8662 19360 8668 19372
rect 8527 19332 8668 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8662 19320 8668 19332
rect 8720 19360 8726 19372
rect 9306 19360 9312 19372
rect 8720 19332 9312 19360
rect 8720 19320 8726 19332
rect 9306 19320 9312 19332
rect 9364 19360 9370 19372
rect 9364 19332 10180 19360
rect 9364 19320 9370 19332
rect 7116 19264 8248 19292
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19261 8355 19295
rect 8297 19255 8355 19261
rect 3476 19196 4660 19224
rect 3476 19184 3482 19196
rect 6362 19184 6368 19236
rect 6420 19224 6426 19236
rect 8110 19224 8116 19236
rect 6420 19196 8116 19224
rect 6420 19184 6426 19196
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 8312 19224 8340 19255
rect 8386 19252 8392 19304
rect 8444 19252 8450 19304
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19292 8631 19295
rect 9766 19292 9772 19304
rect 8619 19264 9772 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 9766 19252 9772 19264
rect 9824 19252 9830 19304
rect 10152 19292 10180 19332
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 10796 19369 10824 19400
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10744 19332 10793 19360
rect 10744 19320 10750 19332
rect 10781 19329 10793 19332
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 10870 19320 10876 19372
rect 10928 19320 10934 19372
rect 11164 19369 11192 19468
rect 12820 19468 14004 19496
rect 11238 19388 11244 19440
rect 11296 19428 11302 19440
rect 12250 19428 12256 19440
rect 11296 19400 12256 19428
rect 11296 19388 11302 19400
rect 12250 19388 12256 19400
rect 12308 19428 12314 19440
rect 12308 19400 12756 19428
rect 12308 19388 12314 19400
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11149 19363 11207 19369
rect 11011 19332 11100 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 11072 19292 11100 19332
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12345 19363 12403 19369
rect 12345 19360 12357 19363
rect 11940 19332 12357 19360
rect 11940 19320 11946 19332
rect 12345 19329 12357 19332
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 10152 19264 11100 19292
rect 12728 19292 12756 19400
rect 12820 19369 12848 19468
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 15105 19499 15163 19505
rect 15105 19465 15117 19499
rect 15151 19465 15163 19499
rect 15105 19459 15163 19465
rect 12912 19400 13768 19428
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 12912 19292 12940 19400
rect 12986 19320 12992 19372
rect 13044 19320 13050 19372
rect 13630 19320 13636 19372
rect 13688 19320 13694 19372
rect 13740 19369 13768 19400
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13981 19363 14039 19369
rect 13981 19360 13993 19363
rect 13725 19323 13783 19329
rect 13832 19332 13993 19360
rect 12728 19264 12940 19292
rect 13648 19292 13676 19320
rect 13832 19292 13860 19332
rect 13981 19329 13993 19332
rect 14027 19329 14039 19363
rect 15120 19360 15148 19459
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 15765 19499 15823 19505
rect 15765 19496 15777 19499
rect 15712 19468 15777 19496
rect 15712 19456 15718 19468
rect 15765 19465 15777 19468
rect 15811 19465 15823 19499
rect 15765 19459 15823 19465
rect 15933 19499 15991 19505
rect 15933 19465 15945 19499
rect 15979 19496 15991 19499
rect 16206 19496 16212 19508
rect 15979 19468 16212 19496
rect 15979 19465 15991 19468
rect 15933 19459 15991 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17589 19499 17647 19505
rect 17589 19496 17601 19499
rect 16816 19468 17601 19496
rect 16816 19456 16822 19468
rect 17589 19465 17601 19468
rect 17635 19465 17647 19499
rect 17589 19459 17647 19465
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 20273 19499 20331 19505
rect 20273 19496 20285 19499
rect 19392 19468 20285 19496
rect 19392 19456 19398 19468
rect 20273 19465 20285 19468
rect 20319 19465 20331 19499
rect 20273 19459 20331 19465
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 23348 19468 23765 19496
rect 23348 19456 23354 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 15562 19388 15568 19440
rect 15620 19388 15626 19440
rect 17218 19388 17224 19440
rect 17276 19388 17282 19440
rect 17421 19431 17479 19437
rect 17421 19428 17433 19431
rect 17328 19400 17433 19428
rect 16942 19360 16948 19372
rect 15120 19332 16948 19360
rect 13981 19323 14039 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17328 19360 17356 19400
rect 17421 19397 17433 19400
rect 17467 19397 17479 19431
rect 17421 19391 17479 19397
rect 20073 19431 20131 19437
rect 20073 19397 20085 19431
rect 20119 19428 20131 19431
rect 22462 19428 22468 19440
rect 20119 19400 22468 19428
rect 20119 19397 20131 19400
rect 20073 19391 20131 19397
rect 20088 19360 20116 19391
rect 22462 19388 22468 19400
rect 22520 19388 22526 19440
rect 22640 19431 22698 19437
rect 22640 19397 22652 19431
rect 22686 19428 22698 19431
rect 23382 19428 23388 19440
rect 22686 19400 23388 19428
rect 22686 19397 22698 19400
rect 22640 19391 22698 19397
rect 23382 19388 23388 19400
rect 23440 19388 23446 19440
rect 17092 19332 17356 19360
rect 17420 19332 20116 19360
rect 22373 19363 22431 19369
rect 17092 19320 17098 19332
rect 13648 19264 13860 19292
rect 9950 19224 9956 19236
rect 8312 19196 9956 19224
rect 9950 19184 9956 19196
rect 10008 19184 10014 19236
rect 11072 19224 11100 19264
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17420 19292 17448 19332
rect 22373 19329 22385 19363
rect 22419 19360 22431 19363
rect 23198 19360 23204 19372
rect 22419 19332 23204 19360
rect 22419 19329 22431 19332
rect 22373 19323 22431 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 24946 19320 24952 19372
rect 25004 19360 25010 19372
rect 25481 19363 25539 19369
rect 25481 19360 25493 19363
rect 25004 19332 25493 19360
rect 25004 19320 25010 19332
rect 25481 19329 25493 19332
rect 25527 19329 25539 19363
rect 25481 19323 25539 19329
rect 17276 19264 17448 19292
rect 17276 19252 17282 19264
rect 25222 19252 25228 19304
rect 25280 19252 25286 19304
rect 11882 19224 11888 19236
rect 11072 19196 11888 19224
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12805 19227 12863 19233
rect 12805 19193 12817 19227
rect 12851 19224 12863 19227
rect 12986 19224 12992 19236
rect 12851 19196 12992 19224
rect 12851 19193 12863 19196
rect 12805 19187 12863 19193
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 19242 19224 19248 19236
rect 17420 19196 19248 19224
rect 3050 19116 3056 19168
rect 3108 19116 3114 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 8478 19156 8484 19168
rect 5316 19128 8484 19156
rect 5316 19116 5322 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 11514 19156 11520 19168
rect 9824 19128 11520 19156
rect 9824 19116 9830 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19156 15807 19159
rect 16114 19156 16120 19168
rect 15795 19128 16120 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 17420 19165 17448 19196
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 17405 19159 17463 19165
rect 17405 19125 17417 19159
rect 17451 19125 17463 19159
rect 17405 19119 17463 19125
rect 20254 19116 20260 19168
rect 20312 19116 20318 19168
rect 20438 19116 20444 19168
rect 20496 19116 20502 19168
rect 25240 19156 25268 19252
rect 25958 19156 25964 19168
rect 25240 19128 25964 19156
rect 25958 19116 25964 19128
rect 26016 19116 26022 19168
rect 26326 19116 26332 19168
rect 26384 19156 26390 19168
rect 26605 19159 26663 19165
rect 26605 19156 26617 19159
rect 26384 19128 26617 19156
rect 26384 19116 26390 19128
rect 26605 19125 26617 19128
rect 26651 19125 26663 19159
rect 26605 19119 26663 19125
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 4157 18955 4215 18961
rect 4157 18921 4169 18955
rect 4203 18921 4215 18955
rect 4157 18915 4215 18921
rect 4172 18884 4200 18915
rect 4338 18912 4344 18964
rect 4396 18912 4402 18964
rect 6454 18912 6460 18964
rect 6512 18912 6518 18964
rect 7009 18955 7067 18961
rect 7009 18921 7021 18955
rect 7055 18952 7067 18955
rect 7098 18952 7104 18964
rect 7055 18924 7104 18952
rect 7055 18921 7067 18924
rect 7009 18915 7067 18921
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8536 18924 8585 18952
rect 8536 18912 8542 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 10410 18912 10416 18964
rect 10468 18952 10474 18964
rect 13998 18952 14004 18964
rect 10468 18924 14004 18952
rect 10468 18912 10474 18924
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 16022 18912 16028 18964
rect 16080 18952 16086 18964
rect 17313 18955 17371 18961
rect 17313 18952 17325 18955
rect 16080 18924 17325 18952
rect 16080 18912 16086 18924
rect 17313 18921 17325 18924
rect 17359 18921 17371 18955
rect 17313 18915 17371 18921
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 20438 18952 20444 18964
rect 20027 18924 20444 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 4798 18884 4804 18896
rect 4172 18856 4804 18884
rect 4798 18844 4804 18856
rect 4856 18844 4862 18896
rect 9125 18887 9183 18893
rect 9125 18884 9137 18887
rect 5736 18856 9137 18884
rect 3050 18776 3056 18828
rect 3108 18816 3114 18828
rect 4338 18816 4344 18828
rect 3108 18788 4344 18816
rect 3108 18776 3114 18788
rect 4338 18776 4344 18788
rect 4396 18816 4402 18828
rect 4890 18816 4896 18828
rect 4396 18788 4896 18816
rect 4396 18776 4402 18788
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 5534 18776 5540 18828
rect 5592 18776 5598 18828
rect 5552 18748 5580 18776
rect 5736 18757 5764 18856
rect 9125 18853 9137 18856
rect 9171 18853 9183 18887
rect 10962 18884 10968 18896
rect 9125 18847 9183 18853
rect 9600 18856 10968 18884
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 5960 18788 7236 18816
rect 5960 18776 5966 18788
rect 3988 18720 5580 18748
rect 5721 18751 5779 18757
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3988 18689 4016 18720
rect 5721 18717 5733 18751
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 5997 18751 6055 18757
rect 5997 18748 6009 18751
rect 5868 18720 6009 18748
rect 5868 18708 5874 18720
rect 5997 18717 6009 18720
rect 6043 18748 6055 18751
rect 6582 18751 6640 18757
rect 6582 18748 6594 18751
rect 6043 18720 6594 18748
rect 6043 18717 6055 18720
rect 5997 18711 6055 18717
rect 6582 18717 6594 18720
rect 6628 18717 6640 18751
rect 6582 18711 6640 18717
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 7208 18748 7236 18788
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7340 18788 8064 18816
rect 7340 18776 7346 18788
rect 8036 18757 8064 18788
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 9600 18816 9628 18856
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 14369 18887 14427 18893
rect 14369 18853 14381 18887
rect 14415 18884 14427 18887
rect 14642 18884 14648 18896
rect 14415 18856 14648 18884
rect 14415 18853 14427 18856
rect 14369 18847 14427 18853
rect 14642 18844 14648 18856
rect 14700 18844 14706 18896
rect 17954 18884 17960 18896
rect 16040 18856 17960 18884
rect 16040 18825 16068 18856
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 18049 18887 18107 18893
rect 18049 18853 18061 18887
rect 18095 18884 18107 18887
rect 20806 18884 20812 18896
rect 18095 18856 20812 18884
rect 18095 18853 18107 18856
rect 18049 18847 18107 18853
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 22741 18887 22799 18893
rect 22741 18853 22753 18887
rect 22787 18884 22799 18887
rect 23566 18884 23572 18896
rect 22787 18856 23572 18884
rect 22787 18853 22799 18856
rect 22741 18847 22799 18853
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 8352 18788 9628 18816
rect 8352 18776 8358 18788
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 7208 18720 7941 18748
rect 7929 18717 7941 18720
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 8022 18751 8080 18757
rect 8022 18717 8034 18751
rect 8068 18717 8080 18751
rect 8022 18711 8080 18717
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8394 18751 8452 18757
rect 8394 18748 8406 18751
rect 8168 18720 8406 18748
rect 8168 18708 8174 18720
rect 8394 18717 8406 18720
rect 8440 18748 8452 18751
rect 9306 18748 9312 18760
rect 8440 18720 9312 18748
rect 8440 18717 8452 18720
rect 8394 18711 8452 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9600 18757 9628 18788
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 16025 18819 16083 18825
rect 10275 18788 11468 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 10091 18720 11008 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 3973 18683 4031 18689
rect 3973 18680 3985 18683
rect 3568 18652 3985 18680
rect 3568 18640 3574 18652
rect 3973 18649 3985 18652
rect 4019 18649 4031 18683
rect 3973 18643 4031 18649
rect 5537 18683 5595 18689
rect 5537 18649 5549 18683
rect 5583 18680 5595 18683
rect 7466 18680 7472 18692
rect 5583 18652 7472 18680
rect 5583 18649 5595 18652
rect 5537 18643 5595 18649
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 7742 18640 7748 18692
rect 7800 18680 7806 18692
rect 8205 18683 8263 18689
rect 8205 18680 8217 18683
rect 7800 18652 8217 18680
rect 7800 18640 7806 18652
rect 8205 18649 8217 18652
rect 8251 18649 8263 18683
rect 8205 18643 8263 18649
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18680 8355 18683
rect 8478 18680 8484 18692
rect 8343 18652 8484 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 8478 18640 8484 18652
rect 8536 18680 8542 18692
rect 8846 18680 8852 18692
rect 8536 18652 8852 18680
rect 8536 18640 8542 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 10060 18680 10088 18711
rect 9416 18652 10088 18680
rect 4183 18615 4241 18621
rect 4183 18581 4195 18615
rect 4229 18612 4241 18615
rect 4982 18612 4988 18624
rect 4229 18584 4988 18612
rect 4229 18581 4241 18584
rect 4183 18575 4241 18581
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 5902 18572 5908 18624
rect 5960 18572 5966 18624
rect 6638 18572 6644 18624
rect 6696 18572 6702 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 9416 18612 9444 18652
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 10781 18683 10839 18689
rect 10781 18680 10793 18683
rect 10468 18652 10793 18680
rect 10468 18640 10474 18652
rect 10781 18649 10793 18652
rect 10827 18649 10839 18683
rect 10781 18643 10839 18649
rect 7616 18584 9444 18612
rect 7616 18572 7622 18584
rect 9490 18572 9496 18624
rect 9548 18572 9554 18624
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10597 18615 10655 18621
rect 10597 18612 10609 18615
rect 10192 18584 10609 18612
rect 10192 18572 10198 18584
rect 10597 18581 10609 18584
rect 10643 18581 10655 18615
rect 10597 18575 10655 18581
rect 10689 18615 10747 18621
rect 10689 18581 10701 18615
rect 10735 18612 10747 18615
rect 10870 18612 10876 18624
rect 10735 18584 10876 18612
rect 10735 18581 10747 18584
rect 10689 18575 10747 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 10980 18612 11008 18720
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11296 18720 11345 18748
rect 11296 18708 11302 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11440 18748 11468 18788
rect 12452 18788 15424 18816
rect 12452 18748 12480 18788
rect 15396 18760 15424 18788
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16172 18788 16436 18816
rect 16172 18776 16178 18788
rect 12802 18748 12808 18760
rect 11440 18720 12480 18748
rect 12544 18720 12808 18748
rect 11333 18711 11391 18717
rect 11600 18683 11658 18689
rect 11600 18649 11612 18683
rect 11646 18680 11658 18683
rect 12544 18680 12572 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 14274 18748 14280 18760
rect 12912 18720 14280 18748
rect 12912 18692 12940 18720
rect 14274 18708 14280 18720
rect 14332 18748 14338 18760
rect 14829 18751 14887 18757
rect 14829 18748 14841 18751
rect 14332 18720 14841 18748
rect 14332 18708 14338 18720
rect 14829 18717 14841 18720
rect 14875 18717 14887 18751
rect 14829 18711 14887 18717
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 16209 18751 16267 18757
rect 16209 18748 16221 18751
rect 15436 18720 16221 18748
rect 15436 18708 15442 18720
rect 16209 18717 16221 18720
rect 16255 18717 16267 18751
rect 16209 18711 16267 18717
rect 16408 18748 16436 18788
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16669 18819 16727 18825
rect 16669 18816 16681 18819
rect 16632 18788 16681 18816
rect 16632 18776 16638 18788
rect 16669 18785 16681 18788
rect 16715 18785 16727 18819
rect 18693 18819 18751 18825
rect 16669 18779 16727 18785
rect 17236 18788 18460 18816
rect 17236 18748 17264 18788
rect 18432 18757 18460 18788
rect 18693 18785 18705 18819
rect 18739 18816 18751 18819
rect 18782 18816 18788 18828
rect 18739 18788 18788 18816
rect 18739 18785 18751 18788
rect 18693 18779 18751 18785
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 20165 18819 20223 18825
rect 20165 18785 20177 18819
rect 20211 18816 20223 18819
rect 23385 18819 23443 18825
rect 20211 18788 21036 18816
rect 20211 18785 20223 18788
rect 20165 18779 20223 18785
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 16408 18720 17264 18748
rect 17354 18720 18245 18748
rect 12894 18680 12900 18692
rect 11646 18652 12572 18680
rect 12636 18652 12900 18680
rect 11646 18649 11658 18652
rect 11600 18643 11658 18649
rect 12636 18612 12664 18652
rect 12894 18640 12900 18652
rect 12952 18640 12958 18692
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 14056 18652 14381 18680
rect 14056 18640 14062 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 15105 18683 15163 18689
rect 15105 18649 15117 18683
rect 15151 18680 15163 18683
rect 16114 18680 16120 18692
rect 15151 18652 16120 18680
rect 15151 18649 15163 18652
rect 15105 18643 15163 18649
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 16298 18640 16304 18692
rect 16356 18640 16362 18692
rect 16408 18689 16436 18720
rect 17354 18717 17417 18720
rect 17354 18714 17371 18717
rect 16574 18689 16580 18692
rect 16393 18683 16451 18689
rect 16393 18649 16405 18683
rect 16439 18649 16451 18683
rect 16393 18643 16451 18649
rect 16531 18683 16580 18689
rect 16531 18649 16543 18683
rect 16577 18649 16580 18683
rect 16531 18643 16580 18649
rect 16574 18640 16580 18643
rect 16632 18640 16638 18692
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 17129 18683 17187 18689
rect 17129 18680 17141 18683
rect 16724 18652 17141 18680
rect 16724 18640 16730 18652
rect 17129 18649 17141 18652
rect 17175 18680 17187 18683
rect 17218 18680 17224 18692
rect 17175 18652 17224 18680
rect 17175 18649 17187 18652
rect 17129 18643 17187 18649
rect 17218 18640 17224 18652
rect 17276 18640 17282 18692
rect 17344 18683 17371 18714
rect 17405 18692 17417 18717
rect 18233 18717 18245 18720
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18874 18748 18880 18760
rect 18463 18720 18880 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 20070 18708 20076 18760
rect 20128 18708 20134 18760
rect 20254 18708 20260 18760
rect 20312 18708 20318 18760
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18717 20499 18751
rect 20441 18711 20499 18717
rect 17405 18683 17408 18692
rect 17344 18652 17408 18683
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 17586 18640 17592 18692
rect 17644 18680 17650 18692
rect 18325 18683 18383 18689
rect 18325 18680 18337 18683
rect 17644 18652 18337 18680
rect 17644 18640 17650 18652
rect 18325 18649 18337 18652
rect 18371 18649 18383 18683
rect 18325 18643 18383 18649
rect 18535 18683 18593 18689
rect 18535 18649 18547 18683
rect 18581 18680 18593 18683
rect 20456 18680 20484 18711
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20772 18720 20913 18748
rect 20772 18708 20778 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 21008 18748 21036 18788
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 25038 18816 25044 18828
rect 23431 18788 25044 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25958 18776 25964 18828
rect 26016 18816 26022 18828
rect 26237 18819 26295 18825
rect 26237 18816 26249 18819
rect 26016 18788 26249 18816
rect 26016 18776 26022 18788
rect 26237 18785 26249 18788
rect 26283 18785 26295 18819
rect 26237 18779 26295 18785
rect 21450 18748 21456 18760
rect 21008 18720 21456 18748
rect 20901 18711 20959 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18748 23075 18751
rect 23474 18748 23480 18760
rect 23063 18720 23480 18748
rect 23063 18717 23075 18720
rect 23017 18711 23075 18717
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 18581 18652 20484 18680
rect 21168 18683 21226 18689
rect 18581 18649 18593 18652
rect 18535 18643 18593 18649
rect 21168 18649 21180 18683
rect 21214 18680 21226 18683
rect 21266 18680 21272 18692
rect 21214 18652 21272 18680
rect 21214 18649 21226 18652
rect 21168 18643 21226 18649
rect 10980 18584 12664 18612
rect 12713 18615 12771 18621
rect 12713 18581 12725 18615
rect 12759 18612 12771 18615
rect 13906 18612 13912 18624
rect 12759 18584 13912 18612
rect 12759 18581 12771 18584
rect 12713 18575 12771 18581
rect 13906 18572 13912 18584
rect 13964 18572 13970 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14921 18615 14979 18621
rect 14921 18612 14933 18615
rect 14792 18584 14933 18612
rect 14792 18572 14798 18584
rect 14921 18581 14933 18584
rect 14967 18581 14979 18615
rect 14921 18575 14979 18581
rect 17494 18572 17500 18624
rect 17552 18572 17558 18624
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18550 18612 18578 18643
rect 21266 18640 21272 18652
rect 21324 18640 21330 18692
rect 23109 18683 23167 18689
rect 22066 18652 22876 18680
rect 18288 18584 18578 18612
rect 19705 18615 19763 18621
rect 18288 18572 18294 18584
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 19978 18612 19984 18624
rect 19751 18584 19984 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 22066 18612 22094 18652
rect 20772 18584 22094 18612
rect 20772 18572 20778 18584
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22244 18584 22293 18612
rect 22244 18572 22250 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22848 18612 22876 18652
rect 23109 18649 23121 18683
rect 23155 18649 23167 18683
rect 23109 18643 23167 18649
rect 23247 18683 23305 18689
rect 23247 18649 23259 18683
rect 23293 18680 23305 18683
rect 24762 18680 24768 18692
rect 23293 18652 24768 18680
rect 23293 18649 23305 18652
rect 23247 18643 23305 18649
rect 23124 18612 23152 18643
rect 24762 18640 24768 18652
rect 24820 18640 24826 18692
rect 26326 18640 26332 18692
rect 26384 18680 26390 18692
rect 26482 18683 26540 18689
rect 26482 18680 26494 18683
rect 26384 18652 26494 18680
rect 26384 18640 26390 18652
rect 26482 18649 26494 18652
rect 26528 18649 26540 18683
rect 26482 18643 26540 18649
rect 22848 18584 23152 18612
rect 22281 18575 22339 18581
rect 27154 18572 27160 18624
rect 27212 18612 27218 18624
rect 27617 18615 27675 18621
rect 27617 18612 27629 18615
rect 27212 18584 27629 18612
rect 27212 18572 27218 18584
rect 27617 18581 27629 18584
rect 27663 18581 27675 18615
rect 27617 18575 27675 18581
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 2958 18368 2964 18420
rect 3016 18368 3022 18420
rect 5261 18411 5319 18417
rect 5261 18377 5273 18411
rect 5307 18408 5319 18411
rect 5994 18408 6000 18420
rect 5307 18380 6000 18408
rect 5307 18377 5319 18380
rect 5261 18371 5319 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 7285 18411 7343 18417
rect 7285 18408 7297 18411
rect 6236 18380 7297 18408
rect 6236 18368 6242 18380
rect 7285 18377 7297 18380
rect 7331 18377 7343 18411
rect 7285 18371 7343 18377
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 9916 18380 10977 18408
rect 9916 18368 9922 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 12618 18408 12624 18420
rect 10965 18371 11023 18377
rect 12406 18380 12624 18408
rect 2976 18340 3004 18368
rect 6733 18343 6791 18349
rect 6733 18340 6745 18343
rect 2976 18312 6745 18340
rect 6733 18309 6745 18312
rect 6779 18340 6791 18343
rect 8846 18340 8852 18352
rect 6779 18312 8852 18340
rect 6779 18309 6791 18312
rect 6733 18303 6791 18309
rect 8846 18300 8852 18312
rect 8904 18300 8910 18352
rect 8938 18300 8944 18352
rect 8996 18340 9002 18352
rect 9950 18340 9956 18352
rect 8996 18312 9956 18340
rect 8996 18300 9002 18312
rect 9950 18300 9956 18312
rect 10008 18300 10014 18352
rect 12406 18340 12434 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 13136 18380 13553 18408
rect 13136 18368 13142 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15528 18380 17540 18408
rect 15528 18368 15534 18380
rect 10336 18312 12434 18340
rect 13449 18343 13507 18349
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3326 18272 3332 18284
rect 3191 18244 3332 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 2976 18204 3004 18235
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 4246 18232 4252 18284
rect 4304 18232 4310 18284
rect 4798 18232 4804 18284
rect 4856 18232 4862 18284
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 3418 18204 3424 18216
rect 2976 18176 3424 18204
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 3050 18028 3056 18080
rect 3108 18028 3114 18080
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6656 18068 6684 18235
rect 7190 18232 7196 18284
rect 7248 18272 7254 18284
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 7248 18244 7573 18272
rect 7248 18232 7254 18244
rect 7561 18241 7573 18244
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 8662 18272 8668 18284
rect 7699 18244 8668 18272
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 10336 18281 10364 18312
rect 13449 18309 13461 18343
rect 13495 18340 13507 18343
rect 13814 18340 13820 18352
rect 13495 18312 13820 18340
rect 13495 18309 13507 18312
rect 13449 18303 13507 18309
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 14706 18343 14764 18349
rect 14706 18340 14718 18343
rect 14148 18312 14718 18340
rect 14148 18300 14154 18312
rect 14706 18309 14718 18312
rect 14752 18309 14764 18343
rect 14706 18303 14764 18309
rect 16022 18300 16028 18352
rect 16080 18340 16086 18352
rect 17221 18343 17279 18349
rect 17221 18340 17233 18343
rect 16080 18312 17233 18340
rect 16080 18300 16086 18312
rect 17221 18309 17233 18312
rect 17267 18309 17279 18343
rect 17221 18303 17279 18309
rect 10321 18275 10379 18281
rect 10321 18272 10333 18275
rect 9364 18244 10333 18272
rect 9364 18232 9370 18244
rect 10321 18241 10333 18244
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 10468 18244 10513 18272
rect 10468 18232 10474 18244
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 10686 18232 10692 18284
rect 10744 18232 10750 18284
rect 10827 18275 10885 18281
rect 10827 18241 10839 18275
rect 10873 18272 10885 18275
rect 10962 18272 10968 18284
rect 10873 18244 10968 18272
rect 10873 18241 10885 18244
rect 10827 18235 10885 18241
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18272 14519 18275
rect 14550 18272 14556 18284
rect 14507 18244 14556 18272
rect 14507 18241 14519 18244
rect 14461 18235 14519 18241
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 15528 18244 17049 18272
rect 15528 18232 15534 18244
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18173 7527 18207
rect 7469 18167 7527 18173
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 12710 18204 12716 18216
rect 7791 18176 12716 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 7484 18136 7512 18167
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 8570 18136 8576 18148
rect 7484 18108 8576 18136
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 16206 18096 16212 18148
rect 16264 18136 16270 18148
rect 16574 18136 16580 18148
rect 16264 18108 16580 18136
rect 16264 18096 16270 18108
rect 16574 18096 16580 18108
rect 16632 18096 16638 18148
rect 17052 18136 17080 18235
rect 17126 18232 17132 18284
rect 17184 18232 17190 18284
rect 17310 18232 17316 18284
rect 17368 18281 17374 18284
rect 17368 18275 17397 18281
rect 17385 18241 17397 18275
rect 17368 18235 17397 18241
rect 17368 18232 17374 18235
rect 17512 18213 17540 18380
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 22373 18411 22431 18417
rect 22373 18408 22385 18411
rect 20128 18380 22385 18408
rect 20128 18368 20134 18380
rect 22373 18377 22385 18380
rect 22419 18377 22431 18411
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 22373 18371 22431 18377
rect 22480 18380 25421 18408
rect 18417 18343 18475 18349
rect 18417 18309 18429 18343
rect 18463 18340 18475 18343
rect 20622 18340 20628 18352
rect 18463 18312 20628 18340
rect 18463 18309 18475 18312
rect 18417 18303 18475 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 21358 18300 21364 18352
rect 21416 18340 21422 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21416 18312 22017 18340
rect 21416 18300 21422 18312
rect 22005 18309 22017 18312
rect 22051 18309 22063 18343
rect 22005 18303 22063 18309
rect 22094 18300 22100 18352
rect 22152 18340 22158 18352
rect 22205 18343 22263 18349
rect 22205 18340 22217 18343
rect 22152 18312 22217 18340
rect 22152 18300 22158 18312
rect 22205 18309 22217 18312
rect 22251 18309 22263 18343
rect 22205 18303 22263 18309
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 18012 18244 18061 18272
rect 18012 18232 18018 18244
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 18138 18232 18144 18284
rect 18196 18232 18202 18284
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 18288 18244 18337 18272
rect 18288 18232 18294 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 18555 18275 18613 18281
rect 18555 18241 18567 18275
rect 18601 18272 18613 18275
rect 18601 18244 19196 18272
rect 18601 18241 18613 18244
rect 18555 18235 18613 18241
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 19168 18204 19196 18244
rect 19242 18232 19248 18284
rect 19300 18232 19306 18284
rect 19334 18232 19340 18284
rect 19392 18232 19398 18284
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 22480 18272 22508 18380
rect 25409 18377 25421 18380
rect 25455 18377 25467 18411
rect 25409 18371 25467 18377
rect 23284 18343 23342 18349
rect 23284 18309 23296 18343
rect 23330 18340 23342 18343
rect 23474 18340 23480 18352
rect 23330 18312 23480 18340
rect 23330 18309 23342 18312
rect 23284 18303 23342 18309
rect 23474 18300 23480 18312
rect 23532 18340 23538 18352
rect 23842 18340 23848 18352
rect 23532 18312 23848 18340
rect 23532 18300 23538 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 24762 18300 24768 18352
rect 24820 18340 24826 18352
rect 25041 18343 25099 18349
rect 25041 18340 25053 18343
rect 24820 18312 25053 18340
rect 24820 18300 24826 18312
rect 25041 18309 25053 18312
rect 25087 18309 25099 18343
rect 25041 18303 25099 18309
rect 25133 18343 25191 18349
rect 25133 18309 25145 18343
rect 25179 18340 25191 18343
rect 26878 18340 26884 18352
rect 25179 18312 26884 18340
rect 25179 18309 25191 18312
rect 25133 18303 25191 18309
rect 26878 18300 26884 18312
rect 26936 18300 26942 18352
rect 21140 18244 22508 18272
rect 21140 18232 21146 18244
rect 24854 18232 24860 18284
rect 24912 18232 24918 18284
rect 25225 18275 25283 18281
rect 25225 18241 25237 18275
rect 25271 18241 25283 18275
rect 25225 18235 25283 18241
rect 19168 18176 19564 18204
rect 17497 18167 17555 18173
rect 17402 18136 17408 18148
rect 17052 18108 17408 18136
rect 17402 18096 17408 18108
rect 17460 18096 17466 18148
rect 9217 18071 9275 18077
rect 9217 18068 9229 18071
rect 6604 18040 9229 18068
rect 6604 18028 6610 18040
rect 9217 18037 9229 18040
rect 9263 18068 9275 18071
rect 9674 18068 9680 18080
rect 9263 18040 9680 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 13446 18068 13452 18080
rect 10192 18040 13452 18068
rect 10192 18028 10198 18040
rect 13446 18028 13452 18040
rect 13504 18068 13510 18080
rect 14642 18068 14648 18080
rect 13504 18040 14648 18068
rect 13504 18028 13510 18040
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 15841 18071 15899 18077
rect 15841 18037 15853 18071
rect 15887 18068 15899 18071
rect 15930 18068 15936 18080
rect 15887 18040 15936 18068
rect 15887 18037 15899 18040
rect 15841 18031 15899 18037
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16853 18071 16911 18077
rect 16853 18037 16865 18071
rect 16899 18068 16911 18071
rect 17678 18068 17684 18080
rect 16899 18040 17684 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 19536 18077 19564 18176
rect 23014 18164 23020 18216
rect 23072 18164 23078 18216
rect 24118 18164 24124 18216
rect 24176 18204 24182 18216
rect 25240 18204 25268 18235
rect 24176 18176 25268 18204
rect 24176 18164 24182 18176
rect 18693 18071 18751 18077
rect 18693 18068 18705 18071
rect 18012 18040 18705 18068
rect 18012 18028 18018 18040
rect 18693 18037 18705 18040
rect 18739 18037 18751 18071
rect 18693 18031 18751 18037
rect 19521 18071 19579 18077
rect 19521 18037 19533 18071
rect 19567 18068 19579 18071
rect 20438 18068 20444 18080
rect 19567 18040 20444 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 22189 18071 22247 18077
rect 22189 18037 22201 18071
rect 22235 18068 22247 18071
rect 23934 18068 23940 18080
rect 22235 18040 23940 18068
rect 22235 18037 22247 18040
rect 22189 18031 22247 18037
rect 23934 18028 23940 18040
rect 23992 18028 23998 18080
rect 24394 18028 24400 18080
rect 24452 18028 24458 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 2682 17824 2688 17876
rect 2740 17864 2746 17876
rect 2869 17867 2927 17873
rect 2869 17864 2881 17867
rect 2740 17836 2881 17864
rect 2740 17824 2746 17836
rect 2869 17833 2881 17836
rect 2915 17833 2927 17867
rect 2869 17827 2927 17833
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3200 17836 3341 17864
rect 3200 17824 3206 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 5718 17824 5724 17876
rect 5776 17824 5782 17876
rect 5905 17867 5963 17873
rect 5905 17833 5917 17867
rect 5951 17864 5963 17867
rect 6362 17864 6368 17876
rect 5951 17836 6368 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7282 17864 7288 17876
rect 7239 17836 7288 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 10870 17864 10876 17876
rect 10183 17836 10876 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10870 17824 10876 17836
rect 10928 17864 10934 17876
rect 12345 17867 12403 17873
rect 10928 17836 11468 17864
rect 10928 17824 10934 17836
rect 6457 17799 6515 17805
rect 6457 17765 6469 17799
rect 6503 17796 6515 17799
rect 10410 17796 10416 17808
rect 6503 17768 10416 17796
rect 6503 17765 6515 17768
rect 6457 17759 6515 17765
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 1670 17688 1676 17740
rect 1728 17728 1734 17740
rect 3053 17731 3111 17737
rect 3053 17728 3065 17731
rect 1728 17700 3065 17728
rect 1728 17688 1734 17700
rect 3053 17697 3065 17700
rect 3099 17728 3111 17731
rect 4246 17728 4252 17740
rect 3099 17700 4252 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 4246 17688 4252 17700
rect 4304 17728 4310 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4304 17700 4445 17728
rect 4304 17688 4310 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17728 4583 17731
rect 4798 17728 4804 17740
rect 4571 17700 4804 17728
rect 4571 17697 4583 17700
rect 4525 17691 4583 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 5718 17688 5724 17740
rect 5776 17728 5782 17740
rect 5776 17700 6684 17728
rect 5776 17688 5782 17700
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 2832 17632 3985 17660
rect 2832 17620 2838 17632
rect 3973 17629 3985 17632
rect 4019 17660 4031 17663
rect 4982 17660 4988 17672
rect 4019 17632 4988 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4982 17620 4988 17632
rect 5040 17660 5046 17672
rect 6656 17669 6684 17700
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 6972 17700 7512 17728
rect 6972 17688 6978 17700
rect 7484 17672 7512 17700
rect 6641 17663 6699 17669
rect 5040 17632 5764 17660
rect 5040 17620 5046 17632
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 2648 17564 5396 17592
rect 2648 17552 2654 17564
rect 4157 17527 4215 17533
rect 4157 17493 4169 17527
rect 4203 17524 4215 17527
rect 5074 17524 5080 17536
rect 4203 17496 5080 17524
rect 4203 17493 4215 17496
rect 4157 17487 4215 17493
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 5368 17524 5396 17564
rect 5442 17552 5448 17604
rect 5500 17592 5506 17604
rect 5736 17601 5764 17632
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17660 6791 17663
rect 6822 17660 6828 17672
rect 6779 17632 6828 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 6822 17620 6828 17632
rect 6880 17660 6886 17672
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 6880 17632 7389 17660
rect 6880 17620 6886 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7466 17620 7472 17672
rect 7524 17620 7530 17672
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 8202 17660 8208 17672
rect 7791 17632 8208 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 5537 17595 5595 17601
rect 5537 17592 5549 17595
rect 5500 17564 5549 17592
rect 5500 17552 5506 17564
rect 5537 17561 5549 17564
rect 5583 17561 5595 17595
rect 5537 17555 5595 17561
rect 5721 17595 5779 17601
rect 5721 17561 5733 17595
rect 5767 17561 5779 17595
rect 5721 17555 5779 17561
rect 6454 17552 6460 17604
rect 6512 17592 6518 17604
rect 7760 17592 7788 17623
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8343 17632 9536 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 9508 17604 9536 17632
rect 9950 17620 9956 17672
rect 10008 17620 10014 17672
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 10100 17632 10793 17660
rect 10100 17620 10106 17632
rect 10781 17629 10793 17632
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 6512 17564 7788 17592
rect 6512 17552 6518 17564
rect 9306 17552 9312 17604
rect 9364 17552 9370 17604
rect 9490 17552 9496 17604
rect 9548 17552 9554 17604
rect 6914 17524 6920 17536
rect 5368 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 8478 17484 8484 17536
rect 8536 17484 8542 17536
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 9582 17524 9588 17536
rect 9180 17496 9588 17524
rect 9180 17484 9186 17496
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10134 17524 10140 17536
rect 9732 17496 10140 17524
rect 9732 17484 9738 17496
rect 10134 17484 10140 17496
rect 10192 17524 10198 17536
rect 11072 17524 11100 17623
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11204 17632 11345 17660
rect 11204 17620 11210 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11440 17660 11468 17836
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 12434 17864 12440 17876
rect 12391 17836 12440 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 14182 17824 14188 17876
rect 14240 17864 14246 17876
rect 14277 17867 14335 17873
rect 14277 17864 14289 17867
rect 14240 17836 14289 17864
rect 14240 17824 14246 17836
rect 14277 17833 14289 17836
rect 14323 17833 14335 17867
rect 14277 17827 14335 17833
rect 18417 17867 18475 17873
rect 18417 17833 18429 17867
rect 18463 17864 18475 17867
rect 18690 17864 18696 17876
rect 18463 17836 18696 17864
rect 18463 17833 18475 17836
rect 18417 17827 18475 17833
rect 18690 17824 18696 17836
rect 18748 17864 18754 17876
rect 19610 17864 19616 17876
rect 18748 17836 19616 17864
rect 18748 17824 18754 17836
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 22888 17836 22937 17864
rect 22888 17824 22894 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 13725 17799 13783 17805
rect 11532 17768 13676 17796
rect 11532 17737 11560 17768
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 12250 17728 12256 17740
rect 11839 17700 12256 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 12544 17700 13216 17728
rect 12544 17660 12572 17700
rect 11440 17632 12572 17660
rect 11333 17623 11391 17629
rect 12618 17620 12624 17672
rect 12676 17620 12682 17672
rect 12894 17620 12900 17672
rect 12952 17660 12958 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12952 17632 13093 17660
rect 12952 17620 12958 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13188 17660 13216 17700
rect 13446 17688 13452 17740
rect 13504 17688 13510 17740
rect 13648 17660 13676 17768
rect 13725 17765 13737 17799
rect 13771 17796 13783 17799
rect 17034 17796 17040 17808
rect 13771 17768 17040 17796
rect 13771 17765 13783 17768
rect 13725 17759 13783 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 20809 17799 20867 17805
rect 20809 17765 20821 17799
rect 20855 17796 20867 17799
rect 24854 17796 24860 17808
rect 20855 17768 24860 17796
rect 20855 17765 20867 17768
rect 20809 17759 20867 17765
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 18932 17700 19564 17728
rect 18932 17688 18938 17700
rect 13188 17632 13609 17660
rect 13648 17632 14412 17660
rect 13081 17623 13139 17629
rect 12342 17552 12348 17604
rect 12400 17552 12406 17604
rect 12636 17592 12664 17620
rect 13170 17592 13176 17604
rect 12636 17564 13176 17592
rect 13170 17552 13176 17564
rect 13228 17552 13234 17604
rect 13581 17601 13609 17632
rect 13566 17595 13624 17601
rect 13566 17561 13578 17595
rect 13612 17592 13624 17595
rect 14182 17592 14188 17604
rect 13612 17564 14188 17592
rect 13612 17561 13624 17564
rect 13566 17555 13624 17561
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 14384 17592 14412 17632
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14608 17632 14749 17660
rect 14608 17620 14614 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17037 17663 17095 17669
rect 17037 17660 17049 17663
rect 16908 17632 17049 17660
rect 16908 17620 16914 17632
rect 17037 17629 17049 17632
rect 17083 17660 17095 17663
rect 18966 17660 18972 17672
rect 17083 17632 18972 17660
rect 17083 17629 17095 17632
rect 17037 17623 17095 17629
rect 18966 17620 18972 17632
rect 19024 17660 19030 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19024 17632 19441 17660
rect 19024 17620 19030 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19536 17660 19564 17700
rect 26970 17688 26976 17740
rect 27028 17688 27034 17740
rect 20622 17660 20628 17672
rect 19536 17632 20628 17660
rect 19429 17623 19487 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 23014 17620 23020 17672
rect 23072 17660 23078 17672
rect 25041 17663 25099 17669
rect 25041 17660 25053 17663
rect 23072 17632 25053 17660
rect 23072 17620 23078 17632
rect 25041 17629 25053 17632
rect 25087 17660 25099 17663
rect 25866 17660 25872 17672
rect 25087 17632 25872 17660
rect 25087 17629 25099 17632
rect 25041 17623 25099 17629
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 14384 17564 16436 17592
rect 12529 17527 12587 17533
rect 12529 17524 12541 17527
rect 10192 17496 12541 17524
rect 10192 17484 10198 17496
rect 12529 17493 12541 17496
rect 12575 17493 12587 17527
rect 12529 17487 12587 17493
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 13998 17524 14004 17536
rect 13403 17496 14004 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14366 17484 14372 17536
rect 14424 17524 14430 17536
rect 14645 17527 14703 17533
rect 14645 17524 14657 17527
rect 14424 17496 14657 17524
rect 14424 17484 14430 17496
rect 14645 17493 14657 17496
rect 14691 17524 14703 17527
rect 16022 17524 16028 17536
rect 14691 17496 16028 17524
rect 14691 17493 14703 17496
rect 14645 17487 14703 17493
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 16408 17524 16436 17564
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 17282 17595 17340 17601
rect 17282 17592 17294 17595
rect 16540 17564 17294 17592
rect 16540 17552 16546 17564
rect 17282 17561 17294 17564
rect 17328 17561 17340 17595
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 17282 17555 17340 17561
rect 17512 17564 19686 17592
rect 16666 17524 16672 17536
rect 16408 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 16942 17484 16948 17536
rect 17000 17524 17006 17536
rect 17402 17524 17408 17536
rect 17000 17496 17408 17524
rect 17000 17484 17006 17496
rect 17402 17484 17408 17496
rect 17460 17524 17466 17536
rect 17512 17524 17540 17564
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 19674 17555 19732 17561
rect 20162 17552 20168 17604
rect 20220 17592 20226 17604
rect 22094 17592 22100 17604
rect 20220 17564 22100 17592
rect 20220 17552 20226 17564
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22462 17552 22468 17604
rect 22520 17592 22526 17604
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22520 17564 22753 17592
rect 22520 17552 22526 17564
rect 22741 17561 22753 17564
rect 22787 17561 22799 17595
rect 22741 17555 22799 17561
rect 23934 17552 23940 17604
rect 23992 17592 23998 17604
rect 25286 17595 25344 17601
rect 25286 17592 25298 17595
rect 23992 17564 25298 17592
rect 23992 17552 23998 17564
rect 25286 17561 25298 17564
rect 25332 17561 25344 17595
rect 27218 17595 27276 17601
rect 27218 17592 27230 17595
rect 25286 17555 25344 17561
rect 26436 17564 27230 17592
rect 26436 17536 26464 17564
rect 27218 17561 27230 17564
rect 27264 17561 27276 17595
rect 27218 17555 27276 17561
rect 17460 17496 17540 17524
rect 17460 17484 17466 17496
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 20898 17524 20904 17536
rect 18012 17496 20904 17524
rect 18012 17484 18018 17496
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 22941 17527 22999 17533
rect 22941 17524 22953 17527
rect 21048 17496 22953 17524
rect 21048 17484 21054 17496
rect 22941 17493 22953 17496
rect 22987 17493 22999 17527
rect 22941 17487 22999 17493
rect 23109 17527 23167 17533
rect 23109 17493 23121 17527
rect 23155 17524 23167 17527
rect 24026 17524 24032 17536
rect 23155 17496 24032 17524
rect 23155 17493 23167 17496
rect 23109 17487 23167 17493
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 26418 17484 26424 17536
rect 26476 17484 26482 17536
rect 27522 17484 27528 17536
rect 27580 17524 27586 17536
rect 28353 17527 28411 17533
rect 28353 17524 28365 17527
rect 27580 17496 28365 17524
rect 27580 17484 27586 17496
rect 28353 17493 28365 17496
rect 28399 17493 28411 17527
rect 28353 17487 28411 17493
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 3050 17320 3056 17332
rect 2731 17292 3056 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3234 17280 3240 17332
rect 3292 17280 3298 17332
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 5997 17323 6055 17329
rect 3384 17292 4752 17320
rect 3384 17280 3390 17292
rect 4617 17255 4675 17261
rect 4617 17252 4629 17255
rect 2792 17224 4629 17252
rect 1670 17144 1676 17196
rect 1728 17144 1734 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2590 17184 2596 17196
rect 2547 17156 2596 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 2792 17193 2820 17224
rect 4617 17221 4629 17224
rect 4663 17221 4675 17255
rect 4617 17215 4675 17221
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 2924 17156 3433 17184
rect 2924 17144 2930 17156
rect 3421 17153 3433 17156
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3568 17156 3648 17184
rect 3568 17144 3574 17156
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 3620 17116 3648 17156
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 4433 17187 4491 17193
rect 4304 17156 4384 17184
rect 4304 17144 4310 17156
rect 1811 17088 3648 17116
rect 4356 17116 4384 17156
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4724 17184 4752 17292
rect 5997 17289 6009 17323
rect 6043 17320 6055 17323
rect 7006 17320 7012 17332
rect 6043 17292 7012 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8202 17320 8208 17332
rect 7484 17292 8208 17320
rect 5074 17212 5080 17264
rect 5132 17252 5138 17264
rect 5537 17255 5595 17261
rect 5537 17252 5549 17255
rect 5132 17224 5549 17252
rect 5132 17212 5138 17224
rect 5537 17221 5549 17224
rect 5583 17252 5595 17255
rect 6086 17252 6092 17264
rect 5583 17224 6092 17252
rect 5583 17221 5595 17224
rect 5537 17215 5595 17221
rect 6086 17212 6092 17224
rect 6144 17212 6150 17264
rect 7484 17252 7512 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 10042 17320 10048 17332
rect 8404 17292 10048 17320
rect 6932 17224 7512 17252
rect 6932 17196 6960 17224
rect 7558 17212 7564 17264
rect 7616 17252 7622 17264
rect 8113 17255 8171 17261
rect 8113 17252 8125 17255
rect 7616 17224 8125 17252
rect 7616 17212 7622 17224
rect 8113 17221 8125 17224
rect 8159 17221 8171 17255
rect 8113 17215 8171 17221
rect 5813 17187 5871 17193
rect 4479 17156 5488 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4798 17116 4804 17128
rect 4356 17088 4804 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 5460 17116 5488 17156
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5994 17184 6000 17196
rect 5859 17156 6000 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 5721 17119 5779 17125
rect 5460 17088 5580 17116
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 2740 17020 3709 17048
rect 2740 17008 2746 17020
rect 3697 17017 3709 17020
rect 3743 17048 3755 17051
rect 5442 17048 5448 17060
rect 3743 17020 5448 17048
rect 3743 17017 3755 17020
rect 3697 17011 3755 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 1946 16940 1952 16992
rect 2004 16980 2010 16992
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 2004 16952 2329 16980
rect 2004 16940 2010 16952
rect 2317 16949 2329 16952
rect 2363 16949 2375 16983
rect 2317 16943 2375 16949
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 5074 16980 5080 16992
rect 3844 16952 5080 16980
rect 3844 16940 3850 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5552 16989 5580 17088
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 6270 17116 6276 17128
rect 5767 17088 6276 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 6270 17076 6276 17088
rect 6328 17076 6334 17128
rect 7208 17048 7236 17147
rect 7282 17076 7288 17128
rect 7340 17076 7346 17128
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 8404 17116 8432 17292
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 12253 17323 12311 17329
rect 12253 17320 12265 17323
rect 10376 17292 12265 17320
rect 10376 17280 10382 17292
rect 12253 17289 12265 17292
rect 12299 17289 12311 17323
rect 12253 17283 12311 17289
rect 12710 17280 12716 17332
rect 12768 17280 12774 17332
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14734 17320 14740 17332
rect 14240 17292 14740 17320
rect 14240 17280 14246 17292
rect 14734 17280 14740 17292
rect 14792 17320 14798 17332
rect 14829 17323 14887 17329
rect 14829 17320 14841 17323
rect 14792 17292 14841 17320
rect 14792 17280 14798 17292
rect 14829 17289 14841 17292
rect 14875 17289 14887 17323
rect 14829 17283 14887 17289
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 19245 17323 19303 17329
rect 19245 17320 19257 17323
rect 17644 17292 19257 17320
rect 17644 17280 17650 17292
rect 19245 17289 19257 17292
rect 19291 17289 19303 17323
rect 22278 17320 22284 17332
rect 19245 17283 19303 17289
rect 20272 17292 22284 17320
rect 9208 17255 9266 17261
rect 9208 17221 9220 17255
rect 9254 17252 9266 17255
rect 10962 17252 10968 17264
rect 9254 17224 10968 17252
rect 9254 17221 9266 17224
rect 9208 17215 9266 17221
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 11882 17212 11888 17264
rect 11940 17212 11946 17264
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12268 17224 13093 17252
rect 12268 17196 12296 17224
rect 13081 17221 13093 17224
rect 13127 17221 13139 17255
rect 13081 17215 13139 17221
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 15013 17255 15071 17261
rect 15013 17252 15025 17255
rect 14056 17224 15025 17252
rect 14056 17212 14062 17224
rect 15013 17221 15025 17224
rect 15059 17221 15071 17255
rect 15013 17215 15071 17221
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18049 17255 18107 17261
rect 18049 17252 18061 17255
rect 18012 17224 18061 17252
rect 18012 17212 18018 17224
rect 18049 17221 18061 17224
rect 18095 17221 18107 17255
rect 18249 17255 18307 17261
rect 18249 17252 18261 17255
rect 18049 17215 18107 17221
rect 18156 17224 18261 17252
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 9490 17184 9496 17196
rect 8536 17156 9496 17184
rect 8536 17144 8542 17156
rect 9490 17144 9496 17156
rect 9548 17184 9554 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 9548 17156 10793 17184
rect 9548 17144 9554 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 7616 17088 8432 17116
rect 8941 17119 8999 17125
rect 7616 17076 7622 17088
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 8941 17079 8999 17085
rect 8478 17048 8484 17060
rect 7208 17020 8484 17048
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 5537 16983 5595 16989
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 5718 16980 5724 16992
rect 5583 16952 5724 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 8956 16980 8984 17079
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 12084 17116 12112 17147
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12400 17156 12909 17184
rect 12400 17144 12406 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 10008 17088 12112 17116
rect 12912 17116 12940 17147
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 14734 17184 14740 17196
rect 13228 17156 14740 17184
rect 13228 17144 13234 17156
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17770 17184 17776 17196
rect 17092 17156 17776 17184
rect 17092 17144 17098 17156
rect 17770 17144 17776 17156
rect 17828 17184 17834 17196
rect 18156 17184 18184 17224
rect 18249 17221 18261 17224
rect 18295 17221 18307 17255
rect 18249 17215 18307 17221
rect 18690 17212 18696 17264
rect 18748 17252 18754 17264
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 18748 17224 18889 17252
rect 18748 17212 18754 17224
rect 18877 17221 18889 17224
rect 18923 17221 18935 17255
rect 19077 17255 19135 17261
rect 19077 17252 19089 17255
rect 18877 17215 18935 17221
rect 18984 17224 19089 17252
rect 17828 17156 18184 17184
rect 17828 17144 17834 17156
rect 14458 17116 14464 17128
rect 12912 17088 14464 17116
rect 10008 17076 10014 17088
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17116 14611 17119
rect 14642 17116 14648 17128
rect 14599 17088 14648 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 10321 17051 10379 17057
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 11698 17048 11704 17060
rect 10367 17020 11704 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 14366 17008 14372 17060
rect 14424 17048 14430 17060
rect 14568 17048 14596 17079
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14752 17088 14933 17116
rect 14424 17020 14596 17048
rect 14424 17008 14430 17020
rect 10965 16983 11023 16989
rect 10965 16980 10977 16983
rect 8956 16952 10977 16980
rect 10965 16949 10977 16952
rect 11011 16980 11023 16983
rect 11238 16980 11244 16992
rect 11011 16952 11244 16980
rect 11011 16949 11023 16952
rect 10965 16943 11023 16949
rect 11238 16940 11244 16952
rect 11296 16980 11302 16992
rect 11974 16980 11980 16992
rect 11296 16952 11980 16980
rect 11296 16940 11302 16952
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 14752 16980 14780 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 16114 17076 16120 17128
rect 16172 17116 16178 17128
rect 18984 17116 19012 17224
rect 19077 17221 19089 17224
rect 19123 17252 19135 17255
rect 19334 17252 19340 17264
rect 19123 17224 19340 17252
rect 19123 17221 19135 17224
rect 19077 17215 19135 17221
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 20272 17261 20300 17292
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 20257 17255 20315 17261
rect 20257 17221 20269 17255
rect 20303 17221 20315 17255
rect 23290 17252 23296 17264
rect 20257 17215 20315 17221
rect 20640 17224 23296 17252
rect 20162 17144 20168 17196
rect 20220 17144 20226 17196
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 16172 17088 19012 17116
rect 20364 17116 20392 17147
rect 20438 17144 20444 17196
rect 20496 17193 20502 17196
rect 20640 17193 20668 17224
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 24946 17212 24952 17264
rect 25004 17252 25010 17264
rect 25492 17255 25550 17261
rect 25492 17252 25504 17255
rect 25004 17224 25504 17252
rect 25004 17212 25010 17224
rect 25492 17221 25504 17224
rect 25538 17252 25550 17255
rect 26142 17252 26148 17264
rect 25538 17224 26148 17252
rect 25538 17221 25550 17224
rect 25492 17215 25550 17221
rect 26142 17212 26148 17224
rect 26200 17212 26206 17264
rect 20496 17187 20525 17193
rect 20513 17153 20525 17187
rect 20496 17147 20525 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20496 17144 20502 17147
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 21048 17156 21281 17184
rect 21048 17144 21054 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 22272 17187 22330 17193
rect 22272 17153 22284 17187
rect 22318 17184 22330 17187
rect 23658 17184 23664 17196
rect 22318 17156 23664 17184
rect 22318 17153 22330 17156
rect 22272 17147 22330 17153
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25866 17184 25872 17196
rect 25271 17156 25872 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25866 17144 25872 17156
rect 25924 17144 25930 17196
rect 20364 17088 20668 17116
rect 16172 17076 16178 17088
rect 20640 17060 20668 17088
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20956 17088 21097 17116
rect 20956 17076 20962 17088
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 21085 17079 21143 17085
rect 21634 17076 21640 17128
rect 21692 17116 21698 17128
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21692 17088 22017 17116
rect 21692 17076 21698 17088
rect 22005 17085 22017 17088
rect 22051 17085 22063 17119
rect 22005 17079 22063 17085
rect 18046 17008 18052 17060
rect 18104 17048 18110 17060
rect 18417 17051 18475 17057
rect 18417 17048 18429 17051
rect 18104 17020 18429 17048
rect 18104 17008 18110 17020
rect 18417 17017 18429 17020
rect 18463 17017 18475 17051
rect 19886 17048 19892 17060
rect 18417 17011 18475 17017
rect 18984 17020 19892 17048
rect 14332 16952 14780 16980
rect 15197 16983 15255 16989
rect 14332 16940 14338 16952
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 17218 16980 17224 16992
rect 15243 16952 17224 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16980 18291 16983
rect 18984 16980 19012 17020
rect 19886 17008 19892 17020
rect 19944 17008 19950 17060
rect 20622 17008 20628 17060
rect 20680 17008 20686 17060
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 24486 17048 24492 17060
rect 23348 17020 24492 17048
rect 23348 17008 23354 17020
rect 24486 17008 24492 17020
rect 24544 17008 24550 17060
rect 18279 16952 19012 16980
rect 19061 16983 19119 16989
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 19150 16980 19156 16992
rect 19107 16952 19156 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19392 16952 19993 16980
rect 19392 16940 19398 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 21453 16983 21511 16989
rect 21453 16949 21465 16983
rect 21499 16980 21511 16983
rect 23014 16980 23020 16992
rect 21499 16952 23020 16980
rect 21499 16949 21511 16952
rect 21453 16943 21511 16949
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 23385 16983 23443 16989
rect 23385 16980 23397 16983
rect 23164 16952 23397 16980
rect 23164 16940 23170 16952
rect 23385 16949 23397 16952
rect 23431 16949 23443 16983
rect 23385 16943 23443 16949
rect 26605 16983 26663 16989
rect 26605 16949 26617 16983
rect 26651 16980 26663 16983
rect 26878 16980 26884 16992
rect 26651 16952 26884 16980
rect 26651 16949 26663 16952
rect 26605 16943 26663 16949
rect 26878 16940 26884 16952
rect 26936 16940 26942 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1765 16779 1823 16785
rect 1765 16776 1777 16779
rect 1728 16748 1777 16776
rect 1728 16736 1734 16748
rect 1765 16745 1777 16748
rect 1811 16745 1823 16779
rect 1765 16739 1823 16745
rect 5718 16736 5724 16788
rect 5776 16776 5782 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 5776 16748 5825 16776
rect 5776 16736 5782 16748
rect 5813 16745 5825 16748
rect 5859 16745 5871 16779
rect 5813 16739 5871 16745
rect 5997 16779 6055 16785
rect 5997 16745 6009 16779
rect 6043 16776 6055 16779
rect 6178 16776 6184 16788
rect 6043 16748 6184 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6178 16736 6184 16748
rect 6236 16776 6242 16788
rect 6730 16776 6736 16788
rect 6236 16748 6736 16776
rect 6236 16736 6242 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 10318 16776 10324 16788
rect 8260 16748 10324 16776
rect 8260 16736 8266 16748
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11330 16776 11336 16788
rect 11204 16748 11336 16776
rect 11204 16736 11210 16748
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 17126 16736 17132 16788
rect 17184 16776 17190 16788
rect 18782 16776 18788 16788
rect 17184 16748 18788 16776
rect 17184 16736 17190 16748
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 18874 16736 18880 16788
rect 18932 16776 18938 16788
rect 19702 16776 19708 16788
rect 18932 16748 19708 16776
rect 18932 16736 18938 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20438 16776 20444 16788
rect 20088 16748 20444 16776
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 2648 16680 4384 16708
rect 2648 16668 2654 16680
rect 4356 16652 4384 16680
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 7098 16708 7104 16720
rect 4764 16680 7104 16708
rect 4764 16668 4770 16680
rect 7098 16668 7104 16680
rect 7156 16668 7162 16720
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 9122 16708 9128 16720
rect 7331 16680 9128 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 2958 16640 2964 16652
rect 2731 16612 2964 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 4338 16600 4344 16652
rect 4396 16600 4402 16652
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 7300 16640 7328 16671
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 9493 16711 9551 16717
rect 9493 16708 9505 16711
rect 9488 16677 9505 16708
rect 9539 16677 9551 16711
rect 9488 16671 9551 16677
rect 9488 16640 9516 16671
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 9766 16708 9772 16720
rect 9640 16680 9772 16708
rect 9640 16668 9646 16680
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 12526 16708 12532 16720
rect 11256 16680 12532 16708
rect 10226 16640 10232 16652
rect 5316 16612 7328 16640
rect 7392 16612 9516 16640
rect 9600 16612 10232 16640
rect 5316 16600 5322 16612
rect 658 16532 664 16584
rect 716 16572 722 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 716 16544 1593 16572
rect 716 16532 722 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 2222 16532 2228 16584
rect 2280 16572 2286 16584
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2280 16544 2421 16572
rect 2280 16532 2286 16544
rect 2409 16541 2421 16544
rect 2455 16572 2467 16575
rect 2590 16572 2596 16584
rect 2455 16544 2596 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 3326 16532 3332 16584
rect 3384 16532 3390 16584
rect 3418 16532 3424 16584
rect 3476 16572 3482 16584
rect 4246 16572 4252 16584
rect 3476 16544 4252 16572
rect 3476 16532 3482 16544
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16572 4859 16575
rect 6178 16572 6184 16584
rect 4847 16544 6184 16572
rect 4847 16541 4859 16544
rect 4801 16535 4859 16541
rect 3142 16464 3148 16516
rect 3200 16464 3206 16516
rect 4632 16504 4660 16535
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16572 6515 16575
rect 7098 16572 7104 16584
rect 6503 16544 7104 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 3252 16476 4660 16504
rect 3252 16445 3280 16476
rect 5626 16464 5632 16516
rect 5684 16504 5690 16516
rect 5994 16504 6000 16516
rect 5684 16476 6000 16504
rect 5684 16464 5690 16476
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 7392 16504 7420 16612
rect 9600 16584 9628 16612
rect 10226 16600 10232 16612
rect 10284 16640 10290 16652
rect 10284 16612 10456 16640
rect 10284 16600 10290 16612
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7558 16572 7564 16584
rect 7515 16544 7564 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 9217 16575 9275 16581
rect 9217 16572 9229 16575
rect 8720 16544 9229 16572
rect 8720 16532 8726 16544
rect 9217 16541 9229 16544
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 6420 16476 7420 16504
rect 6420 16464 6426 16476
rect 8294 16464 8300 16516
rect 8352 16464 8358 16516
rect 8938 16504 8944 16516
rect 8680 16476 8944 16504
rect 3243 16439 3301 16445
rect 3243 16405 3255 16439
rect 3289 16405 3301 16439
rect 3243 16399 3301 16405
rect 4522 16396 4528 16448
rect 4580 16396 4586 16448
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 5829 16439 5887 16445
rect 5829 16436 5841 16439
rect 4856 16408 5841 16436
rect 4856 16396 4862 16408
rect 5829 16405 5841 16408
rect 5875 16405 5887 16439
rect 5829 16399 5887 16405
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6822 16436 6828 16448
rect 6687 16408 6828 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6822 16396 6828 16408
rect 6880 16436 6886 16448
rect 7006 16436 7012 16448
rect 6880 16408 7012 16436
rect 6880 16396 6886 16408
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 8395 16439 8453 16445
rect 8395 16436 8407 16439
rect 7616 16408 8407 16436
rect 7616 16396 7622 16408
rect 8395 16405 8407 16408
rect 8441 16405 8453 16439
rect 8395 16399 8453 16405
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16436 8539 16439
rect 8680 16436 8708 16476
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 8527 16408 8708 16436
rect 9232 16436 9260 16535
rect 9306 16532 9312 16584
rect 9364 16582 9370 16584
rect 9364 16581 9536 16582
rect 9364 16575 9551 16581
rect 9364 16554 9505 16575
rect 9364 16532 9370 16554
rect 9493 16541 9505 16554
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 9582 16532 9588 16584
rect 9640 16532 9646 16584
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 10428 16581 10456 16612
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16541 10471 16575
rect 10413 16535 10471 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10686 16572 10692 16584
rect 10551 16544 10692 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11057 16575 11115 16581
rect 11057 16541 11069 16575
rect 11103 16572 11115 16575
rect 11256 16572 11284 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 17218 16668 17224 16720
rect 17276 16708 17282 16720
rect 19150 16708 19156 16720
rect 17276 16680 19156 16708
rect 17276 16668 17282 16680
rect 19150 16668 19156 16680
rect 19208 16668 19214 16720
rect 19352 16680 19841 16708
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 12250 16640 12256 16652
rect 11563 16612 12256 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 14792 16612 15025 16640
rect 14792 16600 14798 16612
rect 15013 16609 15025 16612
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16172 16612 17080 16640
rect 16172 16600 16178 16612
rect 11103 16544 11284 16572
rect 11103 16541 11115 16544
rect 11057 16535 11115 16541
rect 11256 16436 11284 16544
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11624 16504 11652 16535
rect 11790 16532 11796 16584
rect 11848 16532 11854 16584
rect 16850 16532 16856 16584
rect 16908 16532 16914 16584
rect 17052 16581 17080 16612
rect 17862 16600 17868 16652
rect 17920 16600 17926 16652
rect 18233 16643 18291 16649
rect 18233 16609 18245 16643
rect 18279 16640 18291 16643
rect 19352 16640 19380 16680
rect 18279 16612 19380 16640
rect 18279 16609 18291 16612
rect 18233 16603 18291 16609
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17828 16544 18061 16572
rect 17828 16532 17834 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 19518 16532 19524 16584
rect 19576 16581 19582 16584
rect 19813 16582 19841 16680
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 20088 16708 20116 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 20806 16736 20812 16788
rect 20864 16736 20870 16788
rect 24210 16776 24216 16788
rect 22480 16748 24216 16776
rect 19944 16680 20116 16708
rect 19944 16668 19950 16680
rect 20088 16640 20116 16680
rect 20165 16711 20223 16717
rect 20165 16677 20177 16711
rect 20211 16708 20223 16711
rect 20211 16680 20944 16708
rect 20211 16677 20223 16680
rect 20165 16671 20223 16677
rect 20916 16649 20944 16680
rect 20901 16643 20959 16649
rect 20088 16612 20576 16640
rect 19576 16535 19586 16581
rect 19614 16575 19672 16581
rect 19614 16541 19626 16575
rect 19660 16541 19672 16575
rect 19813 16572 19932 16582
rect 20027 16575 20085 16581
rect 20027 16572 20039 16575
rect 19813 16554 20039 16572
rect 19904 16544 20039 16554
rect 19614 16535 19672 16541
rect 20027 16541 20039 16544
rect 20073 16572 20085 16575
rect 20438 16572 20444 16584
rect 20073 16544 20444 16572
rect 20073 16541 20085 16544
rect 20027 16535 20085 16541
rect 19576 16532 19582 16535
rect 11882 16504 11888 16516
rect 11624 16476 11888 16504
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 15280 16507 15338 16513
rect 15280 16473 15292 16507
rect 15326 16504 15338 16507
rect 15838 16504 15844 16516
rect 15326 16476 15844 16504
rect 15326 16473 15338 16476
rect 15280 16467 15338 16473
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 18874 16504 18880 16516
rect 17328 16476 18880 16504
rect 17328 16448 17356 16476
rect 18874 16464 18880 16476
rect 18932 16464 18938 16516
rect 9232 16408 11284 16436
rect 8527 16405 8539 16408
rect 8481 16399 8539 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 12066 16436 12072 16448
rect 11848 16408 12072 16436
rect 11848 16396 11854 16408
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 16298 16436 16304 16448
rect 15712 16408 16304 16436
rect 15712 16396 15718 16408
rect 16298 16396 16304 16408
rect 16356 16436 16362 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 16356 16408 16405 16436
rect 16356 16396 16362 16408
rect 16393 16405 16405 16408
rect 16439 16405 16451 16439
rect 16393 16399 16451 16405
rect 17221 16439 17279 16445
rect 17221 16405 17233 16439
rect 17267 16436 17279 16439
rect 17310 16436 17316 16448
rect 17267 16408 17316 16436
rect 17267 16405 17279 16408
rect 17221 16399 17279 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 19629 16436 19657 16535
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 20548 16572 20576 16612
rect 20901 16609 20913 16643
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 21008 16612 21211 16640
rect 21008 16572 21036 16612
rect 20548 16544 21036 16572
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 21183 16572 21211 16612
rect 22281 16575 22339 16581
rect 21183 16544 22248 16572
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 19797 16507 19855 16513
rect 19797 16504 19809 16507
rect 19760 16476 19809 16504
rect 19760 16464 19766 16476
rect 19797 16473 19809 16476
rect 19843 16473 19855 16507
rect 19797 16467 19855 16473
rect 19889 16507 19947 16513
rect 19889 16473 19901 16507
rect 19935 16504 19947 16507
rect 20714 16504 20720 16516
rect 19935 16476 20720 16504
rect 19935 16473 19947 16476
rect 19889 16467 19947 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 20809 16507 20867 16513
rect 20809 16473 20821 16507
rect 20855 16504 20867 16507
rect 22094 16504 22100 16516
rect 20855 16476 22100 16504
rect 20855 16473 20867 16476
rect 20809 16467 20867 16473
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 22220 16504 22248 16544
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22370 16572 22376 16584
rect 22327 16544 22376 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 22480 16581 22508 16748
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 22554 16668 22560 16720
rect 22612 16668 22618 16720
rect 23750 16668 23756 16720
rect 23808 16708 23814 16720
rect 23845 16711 23903 16717
rect 23845 16708 23857 16711
rect 23808 16680 23857 16708
rect 23808 16668 23814 16680
rect 23845 16677 23857 16680
rect 23891 16677 23903 16711
rect 23845 16671 23903 16677
rect 22572 16581 22600 16668
rect 23198 16600 23204 16652
rect 23256 16640 23262 16652
rect 23256 16612 23704 16640
rect 23256 16600 23262 16612
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22649 16575 22707 16581
rect 22649 16541 22661 16575
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22655 16504 22683 16535
rect 23290 16532 23296 16584
rect 23348 16532 23354 16584
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 23676 16581 23704 16612
rect 26970 16600 26976 16652
rect 27028 16600 27034 16652
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 23440 16544 23489 16572
rect 23440 16532 23446 16544
rect 23477 16541 23489 16544
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 24302 16572 24308 16584
rect 23707 16544 24308 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 24302 16532 24308 16544
rect 24360 16532 24366 16584
rect 24578 16532 24584 16584
rect 24636 16532 24642 16584
rect 25130 16572 25136 16584
rect 24780 16544 25136 16572
rect 22220 16476 22683 16504
rect 23569 16507 23627 16513
rect 23569 16473 23581 16507
rect 23615 16504 23627 16507
rect 24780 16504 24808 16544
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 24854 16513 24860 16516
rect 23615 16476 24808 16504
rect 23615 16473 23627 16476
rect 23569 16467 23627 16473
rect 24848 16467 24860 16513
rect 24912 16504 24918 16516
rect 24912 16476 24948 16504
rect 24854 16464 24860 16467
rect 24912 16464 24918 16476
rect 26234 16464 26240 16516
rect 26292 16504 26298 16516
rect 27218 16507 27276 16513
rect 27218 16504 27230 16507
rect 26292 16476 27230 16504
rect 26292 16464 26298 16476
rect 27218 16473 27230 16476
rect 27264 16473 27276 16507
rect 27218 16467 27276 16473
rect 19484 16408 19657 16436
rect 19484 16396 19490 16408
rect 21266 16396 21272 16448
rect 21324 16396 21330 16448
rect 22830 16396 22836 16448
rect 22888 16396 22894 16448
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 25961 16439 26019 16445
rect 25961 16436 25973 16439
rect 23348 16408 25973 16436
rect 23348 16396 23354 16408
rect 25961 16405 25973 16408
rect 26007 16405 26019 16439
rect 25961 16399 26019 16405
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 28353 16439 28411 16445
rect 28353 16436 28365 16439
rect 27120 16408 28365 16436
rect 27120 16396 27126 16408
rect 28353 16405 28365 16408
rect 28399 16405 28411 16439
rect 28353 16399 28411 16405
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 1912 16204 3893 16232
rect 1912 16192 1918 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4801 16235 4859 16241
rect 4801 16201 4813 16235
rect 4847 16232 4859 16235
rect 5810 16232 5816 16244
rect 4847 16204 5816 16232
rect 4847 16201 4859 16204
rect 4801 16195 4859 16201
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 8481 16235 8539 16241
rect 5951 16204 8432 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 5442 16164 5448 16176
rect 5276 16136 5448 16164
rect 1854 16056 1860 16108
rect 1912 16056 1918 16108
rect 2590 16056 2596 16108
rect 2648 16056 2654 16108
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 4982 16096 4988 16108
rect 2832 16068 4988 16096
rect 2832 16056 2838 16068
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5074 16056 5080 16108
rect 5132 16056 5138 16108
rect 5276 16105 5304 16136
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 6178 16164 6184 16176
rect 5828 16136 6184 16164
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 5828 16105 5856 16136
rect 6178 16124 6184 16136
rect 6236 16124 6242 16176
rect 7558 16164 7564 16176
rect 6748 16136 7564 16164
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6086 16096 6092 16108
rect 6043 16068 6092 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 6270 16096 6276 16108
rect 6144 16068 6276 16096
rect 6144 16056 6150 16068
rect 6270 16056 6276 16068
rect 6328 16056 6334 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6748 16105 6776 16136
rect 7558 16124 7564 16136
rect 7616 16124 7622 16176
rect 6697 16099 6776 16105
rect 6697 16065 6709 16099
rect 6743 16068 6776 16099
rect 6825 16099 6883 16105
rect 6743 16065 6755 16068
rect 6697 16059 6755 16065
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 6840 16028 6868 16059
rect 6914 16056 6920 16108
rect 6972 16056 6978 16108
rect 7006 16056 7012 16108
rect 7064 16105 7070 16108
rect 7064 16099 7113 16105
rect 7064 16065 7067 16099
rect 7101 16096 7113 16099
rect 8202 16096 8208 16108
rect 7101 16068 8208 16096
rect 7101 16065 7113 16068
rect 7064 16059 7113 16065
rect 7064 16056 7070 16059
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16065 8355 16099
rect 8297 16059 8355 16065
rect 5592 16000 6868 16028
rect 5592 15988 5598 16000
rect 8110 15988 8116 16040
rect 8168 15988 8174 16040
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 2774 15960 2780 15972
rect 2087 15932 2780 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 3142 15920 3148 15972
rect 3200 15960 3206 15972
rect 5626 15960 5632 15972
rect 3200 15932 5632 15960
rect 3200 15920 3206 15932
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 8312 15960 8340 16059
rect 8404 16028 8432 16204
rect 8481 16201 8493 16235
rect 8527 16232 8539 16235
rect 9674 16232 9680 16244
rect 8527 16204 9680 16232
rect 8527 16201 8539 16204
rect 8481 16195 8539 16201
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10686 16232 10692 16244
rect 10376 16204 10692 16232
rect 10376 16192 10382 16204
rect 10686 16192 10692 16204
rect 10744 16232 10750 16244
rect 10744 16204 11928 16232
rect 10744 16192 10750 16204
rect 8846 16124 8852 16176
rect 8904 16164 8910 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 8904 16136 9321 16164
rect 8904 16124 8910 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 9309 16127 9367 16133
rect 9401 16167 9459 16173
rect 9401 16133 9413 16167
rect 9447 16164 9459 16167
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 9447 16136 11805 16164
rect 9447 16133 9459 16136
rect 9401 16127 9459 16133
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 11900 16164 11928 16204
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 14734 16232 14740 16244
rect 12032 16204 14740 16232
rect 12032 16192 12038 16204
rect 12342 16164 12348 16176
rect 11900 16136 12348 16164
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9030 16096 9036 16108
rect 8812 16068 9036 16096
rect 8812 16056 8818 16068
rect 9030 16056 9036 16068
rect 9088 16096 9094 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 9088 16068 9229 16096
rect 9088 16056 9094 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9766 16096 9772 16108
rect 9723 16068 9772 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 10100 16068 10149 16096
rect 10100 16056 10106 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 9306 16028 9312 16040
rect 8404 16000 9312 16028
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 10152 16028 10180 16059
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 10284 16068 10425 16096
rect 10284 16056 10290 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 10686 16056 10692 16108
rect 10744 16056 10750 16108
rect 11330 16096 11336 16108
rect 11164 16068 11336 16096
rect 10152 16000 10456 16028
rect 10428 15972 10456 16000
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 6236 15932 8340 15960
rect 6236 15920 6242 15932
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9585 15963 9643 15969
rect 9585 15960 9597 15963
rect 9272 15932 9597 15960
rect 9272 15920 9278 15932
rect 9585 15929 9597 15932
rect 9631 15929 9643 15963
rect 9585 15923 9643 15929
rect 10410 15920 10416 15972
rect 10468 15920 10474 15972
rect 11164 15969 11192 16068
rect 11330 16056 11336 16068
rect 11388 16096 11394 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11388 16068 11713 16096
rect 11388 16056 11394 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 6546 15892 6552 15904
rect 5776 15864 6552 15892
rect 5776 15852 5782 15864
rect 6546 15852 6552 15864
rect 6604 15892 6610 15904
rect 6822 15892 6828 15904
rect 6604 15864 6828 15892
rect 6604 15852 6610 15864
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7190 15852 7196 15904
rect 7248 15852 7254 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 8941 15895 8999 15901
rect 8941 15892 8953 15895
rect 8904 15864 8953 15892
rect 8904 15852 8910 15864
rect 8941 15861 8953 15864
rect 8987 15861 8999 15895
rect 8941 15855 8999 15861
rect 10226 15852 10232 15904
rect 10284 15892 10290 15904
rect 11164 15892 11192 15923
rect 10284 15864 11192 15892
rect 11808 15892 11836 16127
rect 11900 16105 11928 16136
rect 12342 16124 12348 16136
rect 12400 16124 12406 16176
rect 12452 16105 12480 16204
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 17954 16232 17960 16244
rect 15672 16204 17960 16232
rect 13722 16124 13728 16176
rect 13780 16164 13786 16176
rect 14277 16167 14335 16173
rect 14277 16164 14289 16167
rect 13780 16136 14289 16164
rect 13780 16124 13786 16136
rect 14277 16133 14289 16136
rect 14323 16133 14335 16167
rect 14277 16127 14335 16133
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 15672 16173 15700 16204
rect 17954 16192 17960 16204
rect 18012 16232 18018 16244
rect 18598 16232 18604 16244
rect 18012 16204 18604 16232
rect 18012 16192 18018 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 22370 16232 22376 16244
rect 19576 16204 22376 16232
rect 19576 16192 19582 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 26326 16232 26332 16244
rect 22520 16204 26332 16232
rect 22520 16192 22526 16204
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 15657 16167 15715 16173
rect 14608 16136 14780 16164
rect 14608 16124 14614 16136
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 12704 16099 12762 16105
rect 12704 16065 12716 16099
rect 12750 16096 12762 16099
rect 12750 16068 14412 16096
rect 12750 16065 12762 16068
rect 12704 16059 12762 16065
rect 14384 16028 14412 16068
rect 14458 16056 14464 16108
rect 14516 16056 14522 16108
rect 14642 16056 14648 16108
rect 14700 16056 14706 16108
rect 14752 16105 14780 16136
rect 15657 16133 15669 16167
rect 15703 16133 15715 16167
rect 18138 16164 18144 16176
rect 15657 16127 15715 16133
rect 15887 16133 15945 16139
rect 15887 16130 15899 16133
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 15872 16099 15899 16130
rect 15933 16099 15945 16133
rect 15872 16096 15945 16099
rect 15436 16093 15945 16096
rect 17144 16136 18144 16164
rect 15436 16068 15900 16093
rect 15436 16056 15442 16068
rect 17144 16028 17172 16136
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 19058 16124 19064 16176
rect 19116 16164 19122 16176
rect 19245 16167 19303 16173
rect 19245 16164 19257 16167
rect 19116 16136 19257 16164
rect 19116 16124 19122 16136
rect 19245 16133 19257 16136
rect 19291 16133 19303 16167
rect 19245 16127 19303 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19392 16136 19437 16164
rect 19392 16124 19398 16136
rect 19978 16124 19984 16176
rect 20036 16164 20042 16176
rect 20073 16167 20131 16173
rect 20073 16164 20085 16167
rect 20036 16136 20085 16164
rect 20036 16124 20042 16136
rect 20073 16133 20085 16136
rect 20119 16133 20131 16167
rect 20073 16127 20131 16133
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 17770 16096 17776 16108
rect 17727 16068 17776 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18690 16096 18696 16108
rect 18064 16068 18696 16096
rect 14384 16000 17172 16028
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17276 16000 17509 16028
rect 17276 15988 17282 16000
rect 17497 15997 17509 16000
rect 17543 16028 17555 16031
rect 18064 16028 18092 16068
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19150 16056 19156 16108
rect 19208 16086 19214 16108
rect 19455 16099 19513 16105
rect 19208 16058 19243 16086
rect 19455 16065 19467 16099
rect 19501 16065 19513 16099
rect 19455 16059 19513 16065
rect 19208 16056 19214 16058
rect 19154 16055 19166 16056
rect 19200 16055 19212 16056
rect 19154 16049 19212 16055
rect 19470 16028 19498 16059
rect 19610 16056 19616 16108
rect 19668 16056 19674 16108
rect 20088 16096 20116 16127
rect 20162 16124 20168 16176
rect 20220 16164 20226 16176
rect 20273 16167 20331 16173
rect 20273 16164 20285 16167
rect 20220 16136 20285 16164
rect 20220 16124 20226 16136
rect 20273 16133 20285 16136
rect 20319 16133 20331 16167
rect 20273 16127 20331 16133
rect 20898 16124 20904 16176
rect 20956 16124 20962 16176
rect 20990 16124 20996 16176
rect 21048 16164 21054 16176
rect 21101 16167 21159 16173
rect 21101 16164 21113 16167
rect 21048 16136 21113 16164
rect 21048 16124 21054 16136
rect 21101 16133 21113 16136
rect 21147 16133 21159 16167
rect 25492 16167 25550 16173
rect 21101 16127 21159 16133
rect 22020 16136 23980 16164
rect 21358 16096 21364 16108
rect 20088 16068 21364 16096
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 22020 16105 22048 16136
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21692 16068 22017 16096
rect 21692 16056 21698 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22261 16099 22319 16105
rect 22261 16096 22273 16099
rect 22005 16059 22063 16065
rect 22112 16068 22273 16096
rect 17543 16000 18092 16028
rect 19260 16000 19498 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 19260 15960 19288 16000
rect 21082 15988 21088 16040
rect 21140 16028 21146 16040
rect 22112 16028 22140 16068
rect 22261 16065 22273 16068
rect 22307 16065 22319 16099
rect 22261 16059 22319 16065
rect 23474 16056 23480 16108
rect 23532 16096 23538 16108
rect 23845 16099 23903 16105
rect 23845 16096 23857 16099
rect 23532 16068 23857 16096
rect 23532 16056 23538 16068
rect 23845 16065 23857 16068
rect 23891 16065 23903 16099
rect 23952 16096 23980 16136
rect 25492 16133 25504 16167
rect 25538 16164 25550 16167
rect 25590 16164 25596 16176
rect 25538 16136 25596 16164
rect 25538 16133 25550 16136
rect 25492 16127 25550 16133
rect 25590 16124 25596 16136
rect 25648 16124 25654 16176
rect 24578 16096 24584 16108
rect 23952 16068 24584 16096
rect 23845 16059 23903 16065
rect 24578 16056 24584 16068
rect 24636 16096 24642 16108
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 24636 16068 25237 16096
rect 24636 16056 24642 16068
rect 25225 16065 25237 16068
rect 25271 16096 25283 16099
rect 25866 16096 25872 16108
rect 25271 16068 25872 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 25866 16056 25872 16068
rect 25924 16096 25930 16108
rect 26970 16096 26976 16108
rect 25924 16068 26976 16096
rect 25924 16056 25930 16068
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 21140 16000 22140 16028
rect 21140 15988 21146 16000
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 24762 16028 24768 16040
rect 23072 16000 24768 16028
rect 23072 15988 23078 16000
rect 24762 15988 24768 16000
rect 24820 16028 24826 16040
rect 25130 16028 25136 16040
rect 24820 16000 25136 16028
rect 24820 15988 24826 16000
rect 25130 15988 25136 16000
rect 25188 15988 25194 16040
rect 18156 15932 19288 15960
rect 18156 15904 18184 15932
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 20441 15963 20499 15969
rect 20441 15960 20453 15963
rect 19392 15932 20453 15960
rect 19392 15920 19398 15932
rect 20441 15929 20453 15932
rect 20487 15929 20499 15963
rect 20441 15923 20499 15929
rect 12618 15892 12624 15904
rect 11808 15864 12624 15892
rect 10284 15852 10290 15864
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 13814 15852 13820 15904
rect 13872 15852 13878 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 15841 15895 15899 15901
rect 15841 15892 15853 15895
rect 15804 15864 15853 15892
rect 15804 15852 15810 15864
rect 15841 15861 15853 15864
rect 15887 15861 15899 15895
rect 15841 15855 15899 15861
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 17770 15892 17776 15904
rect 16071 15864 17776 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18138 15892 18144 15904
rect 17911 15864 18144 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15892 19027 15895
rect 20162 15892 20168 15904
rect 19015 15864 20168 15892
rect 19015 15861 19027 15864
rect 18969 15855 19027 15861
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 20257 15895 20315 15901
rect 20257 15861 20269 15895
rect 20303 15892 20315 15895
rect 20346 15892 20352 15904
rect 20303 15864 20352 15892
rect 20303 15861 20315 15864
rect 20257 15855 20315 15861
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20990 15892 20996 15904
rect 20680 15864 20996 15892
rect 20680 15852 20686 15864
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15892 21143 15895
rect 21174 15892 21180 15904
rect 21131 15864 21180 15892
rect 21131 15861 21143 15864
rect 21085 15855 21143 15861
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 23014 15852 23020 15904
rect 23072 15892 23078 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 23072 15864 23397 15892
rect 23072 15852 23078 15864
rect 23385 15861 23397 15864
rect 23431 15892 23443 15895
rect 23934 15892 23940 15904
rect 23431 15864 23940 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24029 15895 24087 15901
rect 24029 15861 24041 15895
rect 24075 15892 24087 15895
rect 24578 15892 24584 15904
rect 24075 15864 24584 15892
rect 24075 15861 24087 15864
rect 24029 15855 24087 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 26602 15852 26608 15904
rect 26660 15852 26666 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 1820 15660 2881 15688
rect 1820 15648 1826 15660
rect 2869 15657 2881 15660
rect 2915 15688 2927 15691
rect 3970 15688 3976 15700
rect 2915 15660 3976 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4157 15691 4215 15697
rect 4157 15657 4169 15691
rect 4203 15688 4215 15691
rect 4890 15688 4896 15700
rect 4203 15660 4896 15688
rect 4203 15657 4215 15660
rect 4157 15651 4215 15657
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 6546 15688 6552 15700
rect 5583 15660 6552 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 8297 15691 8355 15697
rect 6880 15660 7696 15688
rect 6880 15648 6886 15660
rect 1949 15623 2007 15629
rect 1949 15589 1961 15623
rect 1995 15620 2007 15623
rect 4341 15623 4399 15629
rect 1995 15592 2774 15620
rect 1995 15589 2007 15592
rect 1949 15583 2007 15589
rect 2746 15552 2774 15592
rect 4341 15589 4353 15623
rect 4387 15620 4399 15623
rect 7098 15620 7104 15632
rect 4387 15592 7104 15620
rect 4387 15589 4399 15592
rect 4341 15583 4399 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 7668 15620 7696 15660
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8386 15688 8392 15700
rect 8343 15660 8392 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 9214 15688 9220 15700
rect 8536 15660 9220 15688
rect 8536 15648 8542 15660
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 10042 15688 10048 15700
rect 9508 15660 10048 15688
rect 9508 15620 9536 15660
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10134 15648 10140 15700
rect 10192 15648 10198 15700
rect 12713 15691 12771 15697
rect 11348 15660 12434 15688
rect 7668 15592 9536 15620
rect 9585 15623 9643 15629
rect 5626 15552 5632 15564
rect 2746 15524 5632 15552
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 5718 15512 5724 15564
rect 5776 15512 5782 15564
rect 7466 15552 7472 15564
rect 6012 15524 6592 15552
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15453 1823 15487
rect 1765 15447 1823 15453
rect 1780 15416 1808 15447
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2464 15456 2513 15484
rect 2464 15444 2470 15456
rect 2501 15453 2513 15456
rect 2547 15484 2559 15487
rect 2547 15456 4108 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 1780 15388 3096 15416
rect 2869 15351 2927 15357
rect 2869 15317 2881 15351
rect 2915 15348 2927 15351
rect 2958 15348 2964 15360
rect 2915 15320 2964 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3068 15357 3096 15388
rect 3970 15376 3976 15428
rect 4028 15376 4034 15428
rect 4080 15416 4108 15456
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5132 15456 5457 15484
rect 5132 15444 5138 15456
rect 5445 15453 5457 15456
rect 5491 15484 5503 15487
rect 6012 15484 6040 15524
rect 5491 15456 6040 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6564 15493 6592 15524
rect 6748 15524 7472 15552
rect 6748 15493 6776 15524
rect 7466 15512 7472 15524
rect 7524 15512 7530 15564
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 6144 15456 6469 15484
rect 6144 15444 6150 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 6822 15444 6828 15496
rect 6880 15444 6886 15496
rect 7668 15493 7696 15592
rect 9585 15589 9597 15623
rect 9631 15620 9643 15623
rect 11348 15620 11376 15660
rect 9631 15592 11376 15620
rect 12406 15620 12434 15660
rect 12713 15657 12725 15691
rect 12759 15688 12771 15691
rect 15838 15688 15844 15700
rect 12759 15660 15844 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 17494 15688 17500 15700
rect 16991 15660 17500 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 20622 15688 20628 15700
rect 19444 15660 20628 15688
rect 13354 15620 13360 15632
rect 12406 15592 13360 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 14366 15580 14372 15632
rect 14424 15580 14430 15632
rect 16666 15580 16672 15632
rect 16724 15620 16730 15632
rect 19444 15620 19472 15660
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 20809 15691 20867 15697
rect 20809 15688 20821 15691
rect 20772 15660 20821 15688
rect 20772 15648 20778 15660
rect 20809 15657 20821 15660
rect 20855 15657 20867 15691
rect 20809 15651 20867 15657
rect 22370 15648 22376 15700
rect 22428 15648 22434 15700
rect 26418 15688 26424 15700
rect 24504 15660 26424 15688
rect 16724 15592 19472 15620
rect 16724 15580 16730 15592
rect 8036 15524 10180 15552
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 7801 15487 7859 15493
rect 7801 15453 7813 15487
rect 7847 15484 7859 15487
rect 8036 15484 8064 15524
rect 7847 15456 8064 15484
rect 8159 15487 8217 15493
rect 7847 15453 7859 15456
rect 7801 15447 7859 15453
rect 8159 15453 8171 15487
rect 8205 15484 8217 15487
rect 8294 15484 8300 15496
rect 8205 15456 8300 15484
rect 8205 15453 8217 15456
rect 8159 15447 8217 15453
rect 8294 15444 8300 15456
rect 8352 15484 8358 15496
rect 9030 15484 9036 15496
rect 8352 15456 9036 15484
rect 8352 15444 8358 15456
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 10152 15484 10180 15524
rect 10318 15512 10324 15564
rect 10376 15512 10382 15564
rect 10502 15512 10508 15564
rect 10560 15552 10566 15564
rect 10560 15524 11468 15552
rect 10560 15512 10566 15524
rect 10152 15456 10364 15484
rect 4173 15419 4231 15425
rect 4173 15416 4185 15419
rect 4080 15388 4185 15416
rect 4173 15385 4185 15388
rect 4219 15385 4231 15419
rect 4173 15379 4231 15385
rect 6273 15419 6331 15425
rect 6273 15385 6285 15419
rect 6319 15416 6331 15419
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 6319 15388 7941 15416
rect 6319 15385 6331 15388
rect 6273 15379 6331 15385
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15385 8079 15419
rect 10137 15419 10195 15425
rect 8021 15379 8079 15385
rect 8128 15388 10088 15416
rect 3053 15351 3111 15357
rect 3053 15317 3065 15351
rect 3099 15317 3111 15351
rect 3053 15311 3111 15317
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 5810 15348 5816 15360
rect 5767 15320 5816 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 8036 15348 8064 15379
rect 8128 15360 8156 15388
rect 6052 15320 8064 15348
rect 6052 15308 6058 15320
rect 8110 15308 8116 15360
rect 8168 15308 8174 15360
rect 10060 15348 10088 15388
rect 10137 15385 10149 15419
rect 10183 15416 10195 15419
rect 10226 15416 10232 15428
rect 10183 15388 10232 15416
rect 10183 15385 10195 15388
rect 10137 15379 10195 15385
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 10336 15416 10364 15456
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10870 15484 10876 15496
rect 10468 15456 10876 15484
rect 10468 15444 10474 15456
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 11440 15484 11468 15524
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 12400 15524 17080 15552
rect 12400 15512 12406 15524
rect 11606 15493 11612 15496
rect 11589 15487 11612 15493
rect 11589 15484 11601 15487
rect 11440 15456 11601 15484
rect 11333 15447 11391 15453
rect 11589 15453 11601 15456
rect 11589 15447 11612 15453
rect 11054 15416 11060 15428
rect 10336 15388 11060 15416
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 11348 15416 11376 15447
rect 11606 15444 11612 15447
rect 11664 15444 11670 15496
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14921 15487 14979 15493
rect 14921 15484 14933 15487
rect 14240 15456 14933 15484
rect 14240 15444 14246 15456
rect 14921 15453 14933 15456
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 16298 15484 16304 15496
rect 15795 15456 16304 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16850 15444 16856 15496
rect 16908 15444 16914 15496
rect 17052 15493 17080 15524
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 18230 15552 18236 15564
rect 17460 15524 17816 15552
rect 17460 15512 17466 15524
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15453 17095 15487
rect 17037 15447 17095 15453
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 17310 15484 17316 15496
rect 17267 15456 17316 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 17678 15444 17684 15496
rect 17736 15444 17742 15496
rect 17788 15493 17816 15524
rect 18161 15524 18236 15552
rect 18161 15493 18189 15524
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 18966 15512 18972 15564
rect 19024 15552 19030 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19024 15524 19441 15552
rect 19024 15512 19030 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20772 15524 21864 15552
rect 20772 15512 20778 15524
rect 17774 15487 17832 15493
rect 17774 15453 17786 15487
rect 17820 15453 17832 15487
rect 18146 15487 18204 15493
rect 18146 15484 18158 15487
rect 17774 15447 17832 15453
rect 17880 15456 18158 15484
rect 11974 15416 11980 15428
rect 11348 15388 11980 15416
rect 11974 15376 11980 15388
rect 12032 15376 12038 15428
rect 14274 15376 14280 15428
rect 14332 15416 14338 15428
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 14332 15388 14381 15416
rect 14332 15376 14338 15388
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14369 15379 14427 15385
rect 15933 15419 15991 15425
rect 15933 15385 15945 15419
rect 15979 15416 15991 15419
rect 17880 15416 17908 15456
rect 18146 15453 18158 15456
rect 18192 15453 18204 15487
rect 18146 15447 18204 15453
rect 19628 15456 19840 15484
rect 15979 15388 17908 15416
rect 17957 15419 18015 15425
rect 15979 15385 15991 15388
rect 15933 15379 15991 15385
rect 17957 15385 17969 15419
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 18049 15419 18107 15425
rect 18049 15385 18061 15419
rect 18095 15416 18107 15419
rect 19628 15416 19656 15456
rect 19812 15428 19840 15456
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 21082 15484 21088 15496
rect 20312 15456 21088 15484
rect 20312 15444 20318 15456
rect 21082 15444 21088 15456
rect 21140 15484 21146 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 21140 15456 21465 15484
rect 21140 15444 21146 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 21542 15444 21548 15496
rect 21600 15444 21606 15496
rect 21836 15484 21864 15524
rect 21910 15512 21916 15564
rect 21968 15512 21974 15564
rect 22922 15552 22928 15564
rect 22572 15524 22928 15552
rect 22572 15496 22600 15524
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 23017 15555 23075 15561
rect 23017 15521 23029 15555
rect 23063 15552 23075 15555
rect 24504 15552 24532 15660
rect 26418 15648 26424 15660
rect 26476 15648 26482 15700
rect 23063 15524 24532 15552
rect 23063 15521 23075 15524
rect 23017 15515 23075 15521
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 21836 15456 21956 15484
rect 18095 15388 19656 15416
rect 19696 15419 19754 15425
rect 18095 15385 18107 15388
rect 18049 15379 18107 15385
rect 19696 15385 19708 15419
rect 19742 15385 19754 15419
rect 19696 15379 19754 15385
rect 10502 15348 10508 15360
rect 10060 15320 10508 15348
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 10597 15351 10655 15357
rect 10597 15317 10609 15351
rect 10643 15348 10655 15351
rect 11698 15348 11704 15360
rect 10643 15320 11704 15348
rect 10643 15317 10655 15320
rect 10597 15311 10655 15317
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 13998 15308 14004 15360
rect 14056 15348 14062 15360
rect 14550 15348 14556 15360
rect 14056 15320 14556 15348
rect 14056 15308 14062 15320
rect 14550 15308 14556 15320
rect 14608 15348 14614 15360
rect 14829 15351 14887 15357
rect 14829 15348 14841 15351
rect 14608 15320 14841 15348
rect 14608 15308 14614 15320
rect 14829 15317 14841 15320
rect 14875 15317 14887 15351
rect 14829 15311 14887 15317
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 16114 15348 16120 15360
rect 15151 15320 16120 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 17862 15348 17868 15360
rect 16531 15320 17868 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 17972 15348 18000 15379
rect 18230 15348 18236 15360
rect 17972 15320 18236 15348
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 18322 15308 18328 15360
rect 18380 15308 18386 15360
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 19720 15348 19748 15379
rect 19794 15376 19800 15428
rect 19852 15376 19858 15428
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 21269 15419 21327 15425
rect 21269 15416 21281 15419
rect 20772 15388 21281 15416
rect 20772 15376 20778 15388
rect 21269 15385 21281 15388
rect 21315 15385 21327 15419
rect 21637 15419 21695 15425
rect 21637 15416 21649 15419
rect 21269 15379 21327 15385
rect 21376 15388 21649 15416
rect 19668 15320 19748 15348
rect 19668 15308 19674 15320
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 21376 15348 21404 15388
rect 21637 15385 21649 15388
rect 21683 15385 21695 15419
rect 21637 15379 21695 15385
rect 21726 15376 21732 15428
rect 21784 15425 21790 15428
rect 21784 15419 21813 15425
rect 21801 15385 21813 15419
rect 21784 15379 21813 15385
rect 21784 15376 21790 15379
rect 20956 15320 21404 15348
rect 21928 15348 21956 15456
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22554 15484 22560 15496
rect 22428 15456 22560 15484
rect 22428 15444 22434 15456
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15484 22707 15487
rect 25774 15484 25780 15496
rect 22695 15456 24532 15484
rect 22695 15453 22707 15456
rect 22649 15447 22707 15453
rect 22738 15376 22744 15428
rect 22796 15376 22802 15428
rect 22879 15419 22937 15425
rect 22879 15385 22891 15419
rect 22925 15416 22937 15419
rect 23198 15416 23204 15428
rect 22925 15388 23204 15416
rect 22925 15385 22937 15388
rect 22879 15379 22937 15385
rect 23198 15376 23204 15388
rect 23256 15416 23262 15428
rect 23382 15416 23388 15428
rect 23256 15388 23388 15416
rect 23256 15376 23262 15388
rect 23382 15376 23388 15388
rect 23440 15376 23446 15428
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 23569 15419 23627 15425
rect 23569 15416 23581 15419
rect 23532 15388 23581 15416
rect 23532 15376 23538 15388
rect 23569 15385 23581 15388
rect 23615 15385 23627 15419
rect 23569 15379 23627 15385
rect 23753 15419 23811 15425
rect 23753 15385 23765 15419
rect 23799 15416 23811 15419
rect 24394 15416 24400 15428
rect 23799 15388 24400 15416
rect 23799 15385 23811 15388
rect 23753 15379 23811 15385
rect 24394 15376 24400 15388
rect 24452 15376 24458 15428
rect 24504 15416 24532 15456
rect 24688 15456 25780 15484
rect 24688 15416 24716 15456
rect 25774 15444 25780 15456
rect 25832 15444 25838 15496
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26973 15487 27031 15493
rect 26973 15484 26985 15487
rect 26384 15456 26985 15484
rect 26384 15444 26390 15456
rect 26973 15453 26985 15456
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 24854 15425 24860 15428
rect 24504 15388 24716 15416
rect 24848 15379 24860 15425
rect 24854 15376 24860 15379
rect 24912 15376 24918 15428
rect 26142 15416 26148 15428
rect 25516 15388 26148 15416
rect 22278 15348 22284 15360
rect 21928 15320 22284 15348
rect 20956 15308 20962 15320
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 23400 15348 23428 15376
rect 25516 15348 25544 15388
rect 26142 15376 26148 15388
rect 26200 15376 26206 15428
rect 26602 15376 26608 15428
rect 26660 15416 26666 15428
rect 27218 15419 27276 15425
rect 27218 15416 27230 15419
rect 26660 15388 27230 15416
rect 26660 15376 26666 15388
rect 27218 15385 27230 15388
rect 27264 15385 27276 15419
rect 27218 15379 27276 15385
rect 23400 15320 25544 15348
rect 25590 15308 25596 15360
rect 25648 15348 25654 15360
rect 25961 15351 26019 15357
rect 25961 15348 25973 15351
rect 25648 15320 25973 15348
rect 25648 15308 25654 15320
rect 25961 15317 25973 15320
rect 26007 15317 26019 15351
rect 25961 15311 26019 15317
rect 27430 15308 27436 15360
rect 27488 15348 27494 15360
rect 28353 15351 28411 15357
rect 28353 15348 28365 15351
rect 27488 15320 28365 15348
rect 27488 15308 27494 15320
rect 28353 15317 28365 15320
rect 28399 15317 28411 15351
rect 28353 15311 28411 15317
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 1854 15104 1860 15156
rect 1912 15144 1918 15156
rect 2241 15147 2299 15153
rect 2241 15144 2253 15147
rect 1912 15116 2253 15144
rect 1912 15104 1918 15116
rect 2241 15113 2253 15116
rect 2287 15144 2299 15147
rect 2406 15144 2412 15156
rect 2287 15116 2412 15144
rect 2287 15113 2299 15116
rect 2241 15107 2299 15113
rect 2406 15104 2412 15116
rect 2464 15104 2470 15156
rect 6549 15147 6607 15153
rect 6549 15113 6561 15147
rect 6595 15144 6607 15147
rect 6638 15144 6644 15156
rect 6595 15116 6644 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7340 15116 10364 15144
rect 7340 15104 7346 15116
rect 1762 15036 1768 15088
rect 1820 15076 1826 15088
rect 2041 15079 2099 15085
rect 2041 15076 2053 15079
rect 1820 15048 2053 15076
rect 1820 15036 1826 15048
rect 2041 15045 2053 15048
rect 2087 15045 2099 15079
rect 2041 15039 2099 15045
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 6362 15076 6368 15088
rect 3844 15048 6368 15076
rect 3844 15036 3850 15048
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 7156 15048 9413 15076
rect 7156 15036 7162 15048
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 5040 14980 5089 15008
rect 5040 14968 5046 14980
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 7760 15017 7788 15048
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 5316 14980 6837 15008
rect 5316 14968 5322 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7892 14980 7941 15008
rect 7892 14968 7898 14980
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8570 15008 8576 15020
rect 8067 14980 8576 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 5350 14940 5356 14952
rect 5215 14912 5356 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 6236 14912 6745 14940
rect 6236 14900 6242 14912
rect 6733 14909 6745 14912
rect 6779 14909 6791 14943
rect 6733 14903 6791 14909
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7055 14912 7573 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 5445 14875 5503 14881
rect 5445 14841 5457 14875
rect 5491 14872 5503 14875
rect 5718 14872 5724 14884
rect 5491 14844 5724 14872
rect 5491 14841 5503 14844
rect 5445 14835 5503 14841
rect 5718 14832 5724 14844
rect 5776 14872 5782 14884
rect 6932 14872 6960 14900
rect 5776 14844 6960 14872
rect 5776 14832 5782 14844
rect 8036 14816 8064 14971
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 8684 15011 8742 15017
rect 8684 14977 8696 15011
rect 8730 14977 8742 15011
rect 8684 14971 8742 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2222 14804 2228 14816
rect 1820 14776 2228 14804
rect 1820 14764 1826 14776
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 2406 14764 2412 14816
rect 2464 14764 2470 14816
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 2648 14776 4169 14804
rect 2648 14764 2654 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 5077 14807 5135 14813
rect 5077 14804 5089 14807
rect 4948 14776 5089 14804
rect 4948 14764 4954 14776
rect 5077 14773 5089 14776
rect 5123 14773 5135 14807
rect 5077 14767 5135 14773
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 8018 14804 8024 14816
rect 6788 14776 8024 14804
rect 6788 14764 6794 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8570 14804 8576 14816
rect 8527 14776 8576 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8699 14804 8727 14971
rect 8864 14872 8892 14971
rect 8938 14968 8944 15020
rect 8996 14968 9002 15020
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 9674 14968 9680 15020
rect 9732 14968 9738 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10137 15011 10195 15017
rect 10137 15008 10149 15011
rect 10100 14980 10149 15008
rect 10100 14968 10106 14980
rect 10137 14977 10149 14980
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10230 15011 10288 15017
rect 10230 14977 10242 15011
rect 10276 14977 10288 15011
rect 10230 14971 10288 14977
rect 9473 14943 9531 14949
rect 9473 14909 9485 14943
rect 9519 14940 9531 14943
rect 10244 14940 10272 14971
rect 9519 14912 10272 14940
rect 9519 14909 9531 14912
rect 9473 14903 9531 14909
rect 9214 14872 9220 14884
rect 8864 14844 9220 14872
rect 9214 14832 9220 14844
rect 9272 14872 9278 14884
rect 9858 14872 9864 14884
rect 9272 14844 9864 14872
rect 9272 14832 9278 14844
rect 9858 14832 9864 14844
rect 9916 14872 9922 14884
rect 10226 14872 10232 14884
rect 9916 14844 10232 14872
rect 9916 14832 9922 14844
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 10336 14872 10364 15116
rect 10778 15104 10784 15156
rect 10836 15104 10842 15156
rect 11882 15104 11888 15156
rect 11940 15104 11946 15156
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 17053 15147 17111 15153
rect 17053 15144 17065 15147
rect 16172 15116 17065 15144
rect 16172 15104 16178 15116
rect 17053 15113 17065 15116
rect 17099 15144 17111 15147
rect 21358 15144 21364 15156
rect 17099 15116 21364 15144
rect 17099 15113 17111 15116
rect 17053 15107 17111 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 22554 15104 22560 15156
rect 22612 15153 22618 15156
rect 22612 15147 22631 15153
rect 22619 15113 22631 15147
rect 24302 15144 24308 15156
rect 22612 15107 22631 15113
rect 23860 15116 24308 15144
rect 22612 15104 22618 15107
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 14982 15079 15040 15085
rect 14982 15076 14994 15079
rect 13136 15048 14994 15076
rect 13136 15036 13142 15048
rect 14982 15045 14994 15048
rect 15028 15045 15040 15079
rect 14982 15039 15040 15045
rect 15746 15036 15752 15088
rect 15804 15076 15810 15088
rect 16574 15076 16580 15088
rect 15804 15048 16580 15076
rect 15804 15036 15810 15048
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 16853 15079 16911 15085
rect 16853 15076 16865 15079
rect 16816 15048 16865 15076
rect 16816 15036 16822 15048
rect 16853 15045 16865 15048
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 18693 15079 18751 15085
rect 18693 15045 18705 15079
rect 18739 15076 18751 15079
rect 19242 15076 19248 15088
rect 18739 15048 19248 15076
rect 18739 15045 18751 15048
rect 18693 15039 18751 15045
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 19886 15076 19892 15088
rect 19720 15048 19892 15076
rect 10410 14968 10416 15020
rect 10468 14968 10474 15020
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10643 15011 10701 15017
rect 10643 14977 10655 15011
rect 10689 15008 10701 15011
rect 10778 15008 10784 15020
rect 10689 14980 10784 15008
rect 10689 14977 10701 14980
rect 10643 14971 10701 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11204 14980 11805 15008
rect 11204 14968 11210 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12158 15008 12164 15020
rect 12023 14980 12164 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 14734 14968 14740 15020
rect 14792 14968 14798 15020
rect 15562 14968 15568 15020
rect 15620 15008 15626 15020
rect 15620 14980 16620 15008
rect 15620 14968 15626 14980
rect 16592 14940 16620 14980
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 16724 14980 17877 15008
rect 16724 14968 16730 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 19720 15008 19748 15048
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 20070 15085 20076 15088
rect 20064 15076 20076 15085
rect 20031 15048 20076 15076
rect 20064 15039 20076 15048
rect 20070 15036 20076 15039
rect 20128 15036 20134 15088
rect 20622 15036 20628 15088
rect 20680 15076 20686 15088
rect 23860 15085 23888 15116
rect 24302 15104 24308 15116
rect 24360 15104 24366 15156
rect 22373 15079 22431 15085
rect 22373 15076 22385 15079
rect 20680 15048 22385 15076
rect 20680 15036 20686 15048
rect 22373 15045 22385 15048
rect 22419 15045 22431 15079
rect 22373 15039 22431 15045
rect 23845 15079 23903 15085
rect 23845 15045 23857 15079
rect 23891 15045 23903 15079
rect 23845 15039 23903 15045
rect 23937 15079 23995 15085
rect 23937 15045 23949 15079
rect 23983 15076 23995 15079
rect 24946 15076 24952 15088
rect 23983 15048 24952 15076
rect 23983 15045 23995 15048
rect 23937 15039 23995 15045
rect 24946 15036 24952 15048
rect 25004 15036 25010 15088
rect 25492 15079 25550 15085
rect 25492 15045 25504 15079
rect 25538 15076 25550 15079
rect 26510 15076 26516 15088
rect 25538 15048 26516 15076
rect 25538 15045 25550 15048
rect 25492 15039 25550 15045
rect 26510 15036 26516 15048
rect 26568 15036 26574 15088
rect 22002 15008 22008 15020
rect 17865 14971 17923 14977
rect 18340 14980 19748 15008
rect 19812 14980 22008 15008
rect 16758 14940 16764 14952
rect 16592 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14940 16822 14952
rect 17678 14940 17684 14952
rect 16816 14912 17684 14940
rect 16816 14900 16822 14912
rect 17678 14900 17684 14912
rect 17736 14940 17742 14952
rect 18340 14940 18368 14980
rect 17736 14912 18368 14940
rect 17736 14900 17742 14912
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 19812 14949 19840 14980
rect 22002 14968 22008 14980
rect 22060 15008 22066 15020
rect 23474 15008 23480 15020
rect 22060 14980 23480 15008
rect 22060 14968 22066 14980
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 23566 14968 23572 15020
rect 23624 14968 23630 15020
rect 23750 15017 23756 15020
rect 23717 15011 23756 15017
rect 23717 14977 23729 15011
rect 23717 14971 23756 14977
rect 23750 14968 23756 14971
rect 23808 14968 23814 15020
rect 24118 15017 24124 15020
rect 24075 15011 24124 15017
rect 24075 14977 24087 15011
rect 24121 14977 24124 15011
rect 24075 14971 24124 14977
rect 24118 14968 24124 14971
rect 24176 14968 24182 15020
rect 24394 14968 24400 15020
rect 24452 15008 24458 15020
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 24452 14980 25237 15008
rect 24452 14968 24458 14980
rect 25225 14977 25237 14980
rect 25271 15008 25283 15011
rect 26326 15008 26332 15020
rect 25271 14980 26332 15008
rect 25271 14977 25283 14980
rect 25225 14971 25283 14977
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 19797 14943 19855 14949
rect 19797 14940 19809 14943
rect 19576 14912 19809 14940
rect 19576 14900 19582 14912
rect 19797 14909 19809 14912
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22554 14940 22560 14952
rect 22152 14912 22560 14940
rect 22152 14900 22158 14912
rect 22554 14900 22560 14912
rect 22612 14940 22618 14952
rect 23198 14940 23204 14952
rect 22612 14912 23204 14940
rect 22612 14900 22618 14912
rect 23198 14900 23204 14912
rect 23256 14900 23262 14952
rect 13630 14872 13636 14884
rect 10336 14844 13636 14872
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 18049 14875 18107 14881
rect 15672 14844 17080 14872
rect 10502 14804 10508 14816
rect 8699 14776 10508 14804
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 15672 14804 15700 14844
rect 13964 14776 15700 14804
rect 16117 14807 16175 14813
rect 13964 14764 13970 14776
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 16942 14804 16948 14816
rect 16163 14776 16948 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17052 14813 17080 14844
rect 18049 14841 18061 14875
rect 18095 14872 18107 14875
rect 18966 14872 18972 14884
rect 18095 14844 18972 14872
rect 18095 14841 18107 14844
rect 18049 14835 18107 14841
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 21634 14832 21640 14884
rect 21692 14872 21698 14884
rect 24213 14875 24271 14881
rect 24213 14872 24225 14875
rect 21692 14844 24225 14872
rect 21692 14832 21698 14844
rect 24213 14841 24225 14844
rect 24259 14841 24271 14875
rect 24213 14835 24271 14841
rect 17037 14807 17095 14813
rect 17037 14773 17049 14807
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 17221 14807 17279 14813
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17954 14804 17960 14816
rect 17267 14776 17960 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14804 18843 14807
rect 20898 14804 20904 14816
rect 18831 14776 20904 14804
rect 18831 14773 18843 14776
rect 18785 14767 18843 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21174 14764 21180 14816
rect 21232 14764 21238 14816
rect 22557 14807 22615 14813
rect 22557 14773 22569 14807
rect 22603 14804 22615 14807
rect 22646 14804 22652 14816
rect 22603 14776 22652 14804
rect 22603 14773 22615 14776
rect 22557 14767 22615 14773
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 22738 14764 22744 14816
rect 22796 14764 22802 14816
rect 26605 14807 26663 14813
rect 26605 14773 26617 14807
rect 26651 14804 26663 14807
rect 26786 14804 26792 14816
rect 26651 14776 26792 14804
rect 26651 14773 26663 14776
rect 26605 14767 26663 14773
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3016 14572 3433 14600
rect 3016 14560 3022 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 5442 14600 5448 14612
rect 4387 14572 5448 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 3436 14532 3464 14563
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 5534 14560 5540 14612
rect 5592 14560 5598 14612
rect 7837 14603 7895 14609
rect 7837 14569 7849 14603
rect 7883 14600 7895 14603
rect 10410 14600 10416 14612
rect 7883 14572 10416 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 10652 14572 11713 14600
rect 10652 14560 10658 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 11701 14563 11759 14569
rect 11808 14572 12541 14600
rect 4890 14532 4896 14544
rect 3436 14504 4896 14532
rect 4890 14492 4896 14504
rect 4948 14492 4954 14544
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 7374 14532 7380 14544
rect 5684 14504 7380 14532
rect 5684 14492 5690 14504
rect 7374 14492 7380 14504
rect 7432 14492 7438 14544
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 9125 14535 9183 14541
rect 9125 14532 9137 14535
rect 7708 14504 9137 14532
rect 7708 14492 7714 14504
rect 9125 14501 9137 14504
rect 9171 14501 9183 14535
rect 9125 14495 9183 14501
rect 9488 14504 9674 14532
rect 2869 14467 2927 14473
rect 2869 14464 2881 14467
rect 2746 14436 2881 14464
rect 566 14356 572 14408
rect 624 14396 630 14408
rect 1581 14399 1639 14405
rect 1581 14396 1593 14399
rect 624 14368 1593 14396
rect 624 14356 630 14368
rect 1581 14365 1593 14368
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 2746 14396 2774 14436
rect 2869 14433 2881 14436
rect 2915 14464 2927 14467
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 2915 14436 3985 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 3973 14433 3985 14436
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 6730 14464 6736 14476
rect 5040 14436 5856 14464
rect 5040 14424 5046 14436
rect 1912 14368 2774 14396
rect 3237 14399 3295 14405
rect 1912 14356 1918 14368
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 5350 14396 5356 14408
rect 3283 14368 5356 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 5828 14405 5856 14436
rect 6012 14436 6736 14464
rect 6012 14405 6040 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 6880 14436 7236 14464
rect 6880 14424 6886 14436
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5684 14368 5733 14396
rect 5684 14356 5690 14368
rect 5721 14365 5733 14368
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7006 14396 7012 14408
rect 6963 14368 7012 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4341 14331 4399 14337
rect 4341 14328 4353 14331
rect 4028 14300 4353 14328
rect 4028 14288 4034 14300
rect 4341 14297 4353 14300
rect 4387 14297 4399 14331
rect 4341 14291 4399 14297
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 6104 14328 6132 14359
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7208 14405 7236 14436
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 9488 14464 9516 14504
rect 7340 14436 8156 14464
rect 7340 14424 7346 14436
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 8128 14405 8156 14436
rect 8496 14436 9516 14464
rect 9646 14464 9674 14504
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 11808 14532 11836 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 12529 14563 12587 14569
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16945 14603 17003 14609
rect 16945 14600 16957 14603
rect 16632 14572 16957 14600
rect 16632 14560 16638 14572
rect 16945 14569 16957 14572
rect 16991 14569 17003 14603
rect 16945 14563 17003 14569
rect 17770 14560 17776 14612
rect 17828 14560 17834 14612
rect 17865 14603 17923 14609
rect 17865 14569 17877 14603
rect 17911 14600 17923 14603
rect 21266 14600 21272 14612
rect 17911 14572 21272 14600
rect 17911 14569 17923 14572
rect 17865 14563 17923 14569
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 21450 14560 21456 14612
rect 21508 14600 21514 14612
rect 22370 14600 22376 14612
rect 21508 14572 22376 14600
rect 21508 14560 21514 14572
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 11112 14504 11836 14532
rect 11112 14492 11118 14504
rect 11882 14492 11888 14544
rect 11940 14532 11946 14544
rect 13814 14532 13820 14544
rect 11940 14504 13820 14532
rect 11940 14492 11946 14504
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14532 17739 14535
rect 18046 14532 18052 14544
rect 17727 14504 18052 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 18785 14535 18843 14541
rect 18785 14501 18797 14535
rect 18831 14532 18843 14535
rect 18874 14532 18880 14544
rect 18831 14504 18880 14532
rect 18831 14501 18843 14504
rect 18785 14495 18843 14501
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 19702 14492 19708 14544
rect 19760 14492 19766 14544
rect 23753 14535 23811 14541
rect 23753 14501 23765 14535
rect 23799 14501 23811 14535
rect 23753 14495 23811 14501
rect 9646 14436 11376 14464
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7708 14368 8033 14396
rect 7708 14356 7714 14368
rect 8021 14365 8033 14368
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8294 14356 8300 14408
rect 8352 14356 8358 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 5592 14300 6132 14328
rect 5592 14288 5598 14300
rect 6362 14288 6368 14340
rect 6420 14328 6426 14340
rect 8404 14328 8432 14359
rect 6420 14300 8432 14328
rect 6420 14288 6426 14300
rect 3053 14263 3111 14269
rect 3053 14229 3065 14263
rect 3099 14260 3111 14263
rect 3234 14260 3240 14272
rect 3099 14232 3240 14260
rect 3099 14229 3111 14232
rect 3053 14223 3111 14229
rect 3234 14220 3240 14232
rect 3292 14220 3298 14272
rect 4522 14220 4528 14272
rect 4580 14220 4586 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 6052 14232 6745 14260
rect 6052 14220 6058 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 6733 14223 6791 14229
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 8496 14260 8524 14436
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 9088 14368 9137 14396
rect 9088 14356 9094 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9324 14368 9413 14396
rect 6880 14232 8524 14260
rect 9324 14260 9352 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 9490 14356 9496 14408
rect 9548 14356 9554 14408
rect 11238 14405 11244 14408
rect 9613 14399 9671 14405
rect 9613 14365 9625 14399
rect 9659 14396 9671 14399
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 9659 14365 9674 14396
rect 9613 14359 9674 14365
rect 9646 14340 9674 14359
rect 10888 14368 11069 14396
rect 9646 14300 9680 14340
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 10888 14328 10916 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11205 14399 11244 14405
rect 11205 14365 11217 14399
rect 11205 14359 11244 14365
rect 11238 14356 11244 14359
rect 11296 14356 11302 14408
rect 11348 14405 11376 14436
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 14734 14464 14740 14476
rect 14424 14436 14740 14464
rect 14424 14424 14430 14436
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 21266 14464 21272 14476
rect 16816 14436 21272 14464
rect 16816 14424 16822 14436
rect 21266 14424 21272 14436
rect 21324 14464 21330 14476
rect 22278 14464 22284 14476
rect 21324 14436 22284 14464
rect 21324 14424 21330 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 11561 14399 11619 14405
rect 11561 14365 11573 14399
rect 11607 14396 11619 14399
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 11607 14368 12817 14396
rect 11607 14365 11619 14368
rect 11561 14359 11619 14365
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 14292 14396 14320 14424
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14292 14368 14565 14396
rect 12805 14359 12863 14365
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14396 15623 14399
rect 16666 14396 16672 14408
rect 15611 14368 16672 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 11578 14328 11606 14359
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17460 14368 18153 14396
rect 17460 14356 17466 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14396 18659 14399
rect 19702 14396 19708 14408
rect 18647 14368 19708 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 21174 14356 21180 14408
rect 21232 14396 21238 14408
rect 21453 14399 21511 14405
rect 21453 14396 21465 14399
rect 21232 14368 21465 14396
rect 21232 14356 21238 14368
rect 21453 14365 21465 14368
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14365 21695 14399
rect 22094 14396 22100 14408
rect 21637 14359 21695 14365
rect 10836 14300 10916 14328
rect 10980 14300 11606 14328
rect 12529 14331 12587 14337
rect 10836 14288 10842 14300
rect 9582 14260 9588 14272
rect 9324 14232 9588 14260
rect 6880 14220 6886 14232
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 9692 14260 9720 14288
rect 10502 14260 10508 14272
rect 9692 14232 10508 14260
rect 10502 14220 10508 14232
rect 10560 14260 10566 14272
rect 10980 14260 11008 14300
rect 12529 14297 12541 14331
rect 12575 14297 12587 14331
rect 12529 14291 12587 14297
rect 10560 14232 11008 14260
rect 10560 14220 10566 14232
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 12544 14260 12572 14291
rect 14182 14288 14188 14340
rect 14240 14328 14246 14340
rect 14277 14331 14335 14337
rect 14277 14328 14289 14331
rect 14240 14300 14289 14328
rect 14240 14288 14246 14300
rect 14277 14297 14289 14300
rect 14323 14297 14335 14331
rect 14277 14291 14335 14297
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 15832 14331 15890 14337
rect 14424 14300 14964 14328
rect 14424 14288 14430 14300
rect 11664 14232 12572 14260
rect 11664 14220 11670 14232
rect 12710 14220 12716 14272
rect 12768 14220 12774 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14550 14260 14556 14272
rect 13872 14232 14556 14260
rect 13872 14220 13878 14232
rect 14550 14220 14556 14232
rect 14608 14260 14614 14272
rect 14936 14269 14964 14300
rect 15832 14297 15844 14331
rect 15878 14328 15890 14331
rect 15930 14328 15936 14340
rect 15878 14300 15936 14328
rect 15878 14297 15890 14300
rect 15832 14291 15890 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14328 19579 14331
rect 20530 14328 20536 14340
rect 19567 14300 20536 14328
rect 19567 14297 19579 14300
rect 19521 14291 19579 14297
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 21082 14288 21088 14340
rect 21140 14328 21146 14340
rect 21652 14328 21680 14359
rect 21140 14300 21680 14328
rect 22066 14356 22100 14396
rect 22152 14356 22158 14408
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14396 22431 14399
rect 22419 14368 22600 14396
rect 22419 14365 22431 14368
rect 22373 14359 22431 14365
rect 21140 14288 21146 14300
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14608 14232 14657 14260
rect 14608 14220 14614 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 14645 14223 14703 14229
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14260 14979 14263
rect 16758 14260 16764 14272
rect 14967 14232 16764 14260
rect 14967 14229 14979 14232
rect 14921 14223 14979 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17405 14263 17463 14269
rect 17405 14260 17417 14263
rect 17092 14232 17417 14260
rect 17092 14220 17098 14232
rect 17405 14229 17417 14232
rect 17451 14229 17463 14263
rect 17405 14223 17463 14229
rect 18046 14220 18052 14272
rect 18104 14220 18110 14272
rect 18322 14220 18328 14272
rect 18380 14260 18386 14272
rect 20990 14260 20996 14272
rect 18380 14232 20996 14260
rect 18380 14220 18386 14232
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21821 14263 21879 14269
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 22066 14260 22094 14356
rect 21867 14232 22094 14260
rect 22572 14260 22600 14368
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23768 14396 23796 14495
rect 26510 14464 26516 14476
rect 25148 14436 26516 14464
rect 23256 14368 23796 14396
rect 23256 14356 23262 14368
rect 24118 14356 24124 14408
rect 24176 14396 24182 14408
rect 24394 14396 24400 14408
rect 24176 14368 24400 14396
rect 24176 14356 24182 14368
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 25148 14405 25176 14436
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 26970 14424 26976 14476
rect 27028 14424 27034 14476
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14365 25191 14399
rect 25133 14359 25191 14365
rect 25222 14356 25228 14408
rect 25280 14396 25286 14408
rect 25501 14399 25559 14405
rect 25501 14396 25513 14399
rect 25280 14368 25513 14396
rect 25280 14356 25286 14368
rect 25501 14365 25513 14368
rect 25547 14365 25559 14399
rect 25501 14359 25559 14365
rect 22646 14337 22652 14340
rect 22640 14291 22652 14337
rect 22704 14328 22710 14340
rect 23290 14328 23296 14340
rect 22704 14300 23296 14328
rect 22646 14288 22652 14291
rect 22704 14288 22710 14300
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 24302 14288 24308 14340
rect 24360 14328 24366 14340
rect 25317 14331 25375 14337
rect 25317 14328 25329 14331
rect 24360 14300 25329 14328
rect 24360 14288 24366 14300
rect 25317 14297 25329 14300
rect 25363 14297 25375 14331
rect 25317 14291 25375 14297
rect 25409 14331 25467 14337
rect 25409 14297 25421 14331
rect 25455 14328 25467 14331
rect 26050 14328 26056 14340
rect 25455 14300 26056 14328
rect 25455 14297 25467 14300
rect 25409 14291 25467 14297
rect 26050 14288 26056 14300
rect 26108 14288 26114 14340
rect 27062 14288 27068 14340
rect 27120 14328 27126 14340
rect 27218 14331 27276 14337
rect 27218 14328 27230 14331
rect 27120 14300 27230 14328
rect 27120 14288 27126 14300
rect 27218 14297 27230 14300
rect 27264 14297 27276 14331
rect 27218 14291 27276 14297
rect 23658 14260 23664 14272
rect 22572 14232 23664 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 24394 14220 24400 14272
rect 24452 14260 24458 14272
rect 25685 14263 25743 14269
rect 25685 14260 25697 14263
rect 24452 14232 25697 14260
rect 24452 14220 24458 14232
rect 25685 14229 25697 14232
rect 25731 14229 25743 14263
rect 25685 14223 25743 14229
rect 28350 14220 28356 14272
rect 28408 14220 28414 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5258 14056 5264 14068
rect 4755 14028 5264 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5960 14028 6009 14056
rect 5960 14016 5966 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 8294 14056 8300 14068
rect 5997 14019 6055 14025
rect 7116 14028 8300 14056
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 7116 13988 7144 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11790 14056 11796 14068
rect 11011 14028 11796 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11790 14016 11796 14028
rect 11848 14056 11854 14068
rect 12342 14056 12348 14068
rect 11848 14028 12348 14056
rect 11848 14016 11854 14028
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 13081 14059 13139 14065
rect 13081 14056 13093 14059
rect 12860 14028 13093 14056
rect 12860 14016 12866 14028
rect 13081 14025 13093 14028
rect 13127 14056 13139 14059
rect 13446 14056 13452 14068
rect 13127 14028 13452 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13630 14016 13636 14068
rect 13688 14016 13694 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 14608 14028 16313 14056
rect 14608 14016 14614 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 16758 14056 16764 14068
rect 16301 14019 16359 14025
rect 16592 14028 16764 14056
rect 4580 13960 7144 13988
rect 4580 13948 4586 13960
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 2464 13892 3525 13920
rect 2464 13880 2470 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4120 13892 5089 13920
rect 4120 13880 4126 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5718 13880 5724 13932
rect 5776 13880 5782 13932
rect 7116 13929 7144 13960
rect 8386 13948 8392 14000
rect 8444 13948 8450 14000
rect 9852 13991 9910 13997
rect 9852 13957 9864 13991
rect 9898 13988 9910 13991
rect 11882 13988 11888 14000
rect 9898 13960 11888 13988
rect 9898 13957 9910 13960
rect 9852 13951 9910 13957
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 13538 13948 13544 14000
rect 13596 13948 13602 14000
rect 13648 13988 13676 14016
rect 13757 13991 13815 13997
rect 13757 13988 13769 13991
rect 13648 13960 13769 13988
rect 13757 13957 13769 13960
rect 13803 13988 13815 13991
rect 13803 13960 14780 13988
rect 13803 13957 13815 13960
rect 13757 13951 13815 13957
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 8113 13923 8171 13929
rect 8113 13920 8125 13923
rect 7800 13892 8125 13920
rect 7800 13880 7806 13892
rect 8113 13889 8125 13892
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 8478 13880 8484 13932
rect 8536 13929 8542 13932
rect 8536 13923 8591 13929
rect 8536 13889 8545 13923
rect 8579 13920 8591 13923
rect 8938 13920 8944 13932
rect 8579 13892 8944 13920
rect 8579 13889 8591 13892
rect 8536 13883 8591 13889
rect 8536 13880 8542 13883
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9030 13880 9036 13932
rect 9088 13920 9094 13932
rect 10778 13920 10784 13932
rect 9088 13892 10784 13920
rect 9088 13880 9094 13892
rect 10778 13880 10784 13892
rect 10836 13920 10842 13932
rect 11606 13920 11612 13932
rect 10836 13892 11612 13920
rect 10836 13880 10842 13892
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11968 13923 12026 13929
rect 11968 13889 11980 13923
rect 12014 13920 12026 13923
rect 12434 13920 12440 13932
rect 12014 13892 12440 13920
rect 12014 13889 12026 13892
rect 11968 13883 12026 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14752 13920 14780 13960
rect 14826 13948 14832 14000
rect 14884 13988 14890 14000
rect 14946 13991 15004 13997
rect 14946 13988 14958 13991
rect 14884 13960 14958 13988
rect 14884 13948 14890 13960
rect 14946 13957 14958 13960
rect 14992 13957 15004 13991
rect 14946 13951 15004 13957
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15804 13960 15945 13988
rect 15804 13948 15810 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 16149 13991 16207 13997
rect 16149 13957 16161 13991
rect 16195 13988 16207 13991
rect 16592 13988 16620 14028
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 17000 14028 18245 14056
rect 17000 14016 17006 14028
rect 18233 14025 18245 14028
rect 18279 14056 18291 14059
rect 18322 14056 18328 14068
rect 18279 14028 18328 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 18506 14016 18512 14068
rect 18564 14056 18570 14068
rect 19334 14056 19340 14068
rect 18564 14028 19340 14056
rect 18564 14016 18570 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 20404 14028 20821 14056
rect 20404 14016 20410 14028
rect 20809 14025 20821 14028
rect 20855 14056 20867 14059
rect 20855 14028 22324 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 16195 13960 16620 13988
rect 16195 13957 16207 13960
rect 16149 13951 16207 13957
rect 17954 13948 17960 14000
rect 18012 13988 18018 14000
rect 19518 13988 19524 14000
rect 18012 13954 18032 13988
rect 18800 13960 19524 13988
rect 18012 13948 18092 13954
rect 16298 13920 16304 13932
rect 14332 13892 14587 13920
rect 14752 13892 16304 13920
rect 14332 13880 14338 13892
rect 4246 13812 4252 13864
rect 4304 13852 4310 13864
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 4304 13824 4905 13852
rect 4304 13812 4310 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13821 5043 13855
rect 4985 13815 5043 13821
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5258 13852 5264 13864
rect 5215 13824 5264 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5000 13784 5028 13815
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5994 13812 6000 13864
rect 6052 13812 6058 13864
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6604 13824 8708 13852
rect 6604 13812 6610 13824
rect 5442 13784 5448 13796
rect 5000 13756 5448 13784
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 5810 13744 5816 13796
rect 5868 13744 5874 13796
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 8680 13793 8708 13824
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9548 13824 9597 13852
rect 9548 13812 9554 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11204 13824 11713 13852
rect 11204 13812 11210 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 13596 13824 14412 13852
rect 13596 13812 13602 13824
rect 7285 13787 7343 13793
rect 7285 13784 7297 13787
rect 6788 13756 7297 13784
rect 6788 13744 6794 13756
rect 7285 13753 7297 13756
rect 7331 13753 7343 13787
rect 7285 13747 7343 13753
rect 8665 13787 8723 13793
rect 8665 13753 8677 13787
rect 8711 13753 8723 13787
rect 8665 13747 8723 13753
rect 13262 13744 13268 13796
rect 13320 13784 13326 13796
rect 14274 13784 14280 13796
rect 13320 13756 14280 13784
rect 13320 13744 13326 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 3697 13719 3755 13725
rect 3697 13685 3709 13719
rect 3743 13716 3755 13719
rect 4982 13716 4988 13728
rect 3743 13688 4988 13716
rect 3743 13685 3755 13688
rect 3697 13679 3755 13685
rect 4982 13676 4988 13688
rect 5040 13716 5046 13728
rect 5258 13716 5264 13728
rect 5040 13688 5264 13716
rect 5040 13676 5046 13688
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 13722 13676 13728 13728
rect 13780 13676 13786 13728
rect 13906 13676 13912 13728
rect 13964 13676 13970 13728
rect 14384 13716 14412 13824
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 14559 13852 14587 13892
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 18004 13929 18092 13948
rect 18004 13926 18107 13929
rect 18049 13923 18107 13926
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18322 13880 18328 13932
rect 18380 13880 18386 13932
rect 18690 13880 18696 13932
rect 18748 13920 18754 13932
rect 18800 13929 18828 13960
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 22005 13991 22063 13997
rect 22005 13988 22017 13991
rect 21192 13960 22017 13988
rect 18785 13923 18843 13929
rect 18785 13920 18797 13923
rect 18748 13892 18797 13920
rect 18748 13880 18754 13892
rect 18785 13889 18797 13892
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 18874 13880 18880 13932
rect 18932 13880 18938 13932
rect 19052 13923 19110 13929
rect 19052 13889 19064 13923
rect 19098 13920 19110 13923
rect 20254 13920 20260 13932
rect 19098 13892 20260 13920
rect 19098 13889 19110 13892
rect 19052 13883 19110 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 20622 13880 20628 13932
rect 20680 13880 20686 13932
rect 14734 13852 14740 13864
rect 14559 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 14826 13812 14832 13864
rect 14884 13812 14890 13864
rect 18892 13852 18920 13880
rect 15120 13824 18920 13852
rect 14476 13784 14504 13812
rect 15010 13784 15016 13796
rect 14476 13756 15016 13784
rect 15010 13744 15016 13756
rect 15068 13744 15074 13796
rect 15120 13793 15148 13824
rect 19886 13812 19892 13864
rect 19944 13852 19950 13864
rect 21192 13852 21220 13960
rect 22005 13957 22017 13960
rect 22051 13957 22063 13991
rect 22005 13951 22063 13957
rect 22205 13991 22263 13997
rect 22205 13957 22217 13991
rect 22251 13957 22263 13991
rect 22296 13988 22324 14028
rect 22370 14016 22376 14068
rect 22428 14016 22434 14068
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 24854 14056 24860 14068
rect 22888 14028 24860 14056
rect 22888 14016 22894 14028
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 25501 14059 25559 14065
rect 25501 14025 25513 14059
rect 25547 14056 25559 14059
rect 25774 14056 25780 14068
rect 25547 14028 25780 14056
rect 25547 14025 25559 14028
rect 25501 14019 25559 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 26513 14059 26571 14065
rect 26513 14025 26525 14059
rect 26559 14056 26571 14059
rect 26694 14056 26700 14068
rect 26559 14028 26700 14056
rect 26559 14025 26571 14028
rect 26513 14019 26571 14025
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 22462 13988 22468 14000
rect 22296 13960 22468 13988
rect 22205 13951 22263 13957
rect 22220 13920 22248 13951
rect 22462 13948 22468 13960
rect 22520 13988 22526 14000
rect 23290 13988 23296 14000
rect 22520 13960 23296 13988
rect 22520 13948 22526 13960
rect 23290 13948 23296 13960
rect 23348 13948 23354 14000
rect 23523 13957 23581 13963
rect 23523 13954 23535 13957
rect 19944 13824 21220 13852
rect 21376 13892 22248 13920
rect 23508 13923 23535 13954
rect 23569 13923 23581 13957
rect 26142 13948 26148 14000
rect 26200 13948 26206 14000
rect 26234 13948 26240 14000
rect 26292 13948 26298 14000
rect 23508 13917 23581 13923
rect 19944 13812 19950 13824
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13753 15163 13787
rect 15105 13747 15163 13753
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 17770 13784 17776 13796
rect 17276 13756 17776 13784
rect 17276 13744 17282 13756
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 17865 13787 17923 13793
rect 17865 13753 17877 13787
rect 17911 13784 17923 13787
rect 18506 13784 18512 13796
rect 17911 13756 18512 13784
rect 17911 13753 17923 13756
rect 17865 13747 17923 13753
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 20990 13744 20996 13796
rect 21048 13784 21054 13796
rect 21376 13784 21404 13892
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 23508 13852 23536 13917
rect 23658 13880 23664 13932
rect 23716 13920 23722 13932
rect 24118 13920 24124 13932
rect 23716 13892 24124 13920
rect 23716 13880 23722 13892
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 24377 13923 24435 13929
rect 24377 13920 24389 13923
rect 24268 13892 24389 13920
rect 24268 13880 24274 13892
rect 24377 13889 24389 13892
rect 24423 13889 24435 13923
rect 24377 13883 24435 13889
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 21508 13824 23536 13852
rect 25976 13852 26004 13883
rect 26326 13880 26332 13932
rect 26384 13880 26390 13932
rect 27522 13852 27528 13864
rect 25976 13824 27528 13852
rect 21508 13812 21514 13824
rect 27522 13812 27528 13824
rect 27580 13812 27586 13864
rect 27062 13784 27068 13796
rect 21048 13756 21404 13784
rect 23492 13756 24164 13784
rect 21048 13744 21054 13756
rect 15562 13716 15568 13728
rect 14384 13688 15568 13716
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 16117 13719 16175 13725
rect 16117 13685 16129 13719
rect 16163 13716 16175 13719
rect 16390 13716 16396 13728
rect 16163 13688 16396 13716
rect 16163 13685 16175 13688
rect 16117 13679 16175 13685
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 17589 13719 17647 13725
rect 17589 13716 17601 13719
rect 17368 13688 17601 13716
rect 17368 13676 17374 13688
rect 17589 13685 17601 13688
rect 17635 13685 17647 13719
rect 17589 13679 17647 13685
rect 17957 13719 18015 13725
rect 17957 13685 17969 13719
rect 18003 13716 18015 13719
rect 19518 13716 19524 13728
rect 18003 13688 19524 13716
rect 18003 13685 18015 13688
rect 17957 13679 18015 13685
rect 19518 13676 19524 13688
rect 19576 13676 19582 13728
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 20128 13688 20177 13716
rect 20128 13676 20134 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 20165 13679 20223 13685
rect 20898 13676 20904 13728
rect 20956 13716 20962 13728
rect 21358 13716 21364 13728
rect 20956 13688 21364 13716
rect 20956 13676 20962 13688
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22189 13719 22247 13725
rect 22189 13685 22201 13719
rect 22235 13716 22247 13719
rect 23382 13716 23388 13728
rect 22235 13688 23388 13716
rect 22235 13685 22247 13688
rect 22189 13679 22247 13685
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 23492 13725 23520 13756
rect 23477 13719 23535 13725
rect 23477 13685 23489 13719
rect 23523 13685 23535 13719
rect 23477 13679 23535 13685
rect 23658 13676 23664 13728
rect 23716 13676 23722 13728
rect 23750 13676 23756 13728
rect 23808 13716 23814 13728
rect 24026 13716 24032 13728
rect 23808 13688 24032 13716
rect 23808 13676 23814 13688
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24136 13716 24164 13756
rect 25424 13756 27068 13784
rect 25424 13716 25452 13756
rect 27062 13744 27068 13756
rect 27120 13744 27126 13796
rect 24136 13688 25452 13716
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 3973 13515 4031 13521
rect 3973 13481 3985 13515
rect 4019 13512 4031 13515
rect 5718 13512 5724 13524
rect 4019 13484 5724 13512
rect 4019 13481 4031 13484
rect 3973 13475 4031 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 6822 13512 6828 13524
rect 6687 13484 6828 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 8662 13512 8668 13524
rect 7432 13484 8668 13512
rect 7432 13472 7438 13484
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 9640 13484 10609 13512
rect 9640 13472 9646 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 10597 13475 10655 13481
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 10870 13512 10876 13524
rect 10744 13484 10876 13512
rect 10744 13472 10750 13484
rect 10870 13472 10876 13484
rect 10928 13512 10934 13524
rect 10928 13484 13860 13512
rect 10928 13472 10934 13484
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 9214 13444 9220 13456
rect 5675 13416 9220 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 11238 13444 11244 13456
rect 9447 13416 11244 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 4798 13376 4804 13388
rect 4663 13348 4804 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5718 13336 5724 13388
rect 5776 13376 5782 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5776 13348 5825 13376
rect 5776 13336 5782 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 5813 13339 5871 13345
rect 6748 13348 6837 13376
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 3292 13280 4261 13308
rect 3292 13268 3298 13280
rect 4249 13277 4261 13280
rect 4295 13308 4307 13311
rect 4522 13308 4528 13320
rect 4295 13280 4528 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 4982 13308 4988 13320
rect 4755 13280 4988 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5905 13311 5963 13317
rect 5905 13308 5917 13311
rect 5500 13280 5917 13308
rect 5500 13268 5506 13280
rect 5905 13277 5917 13280
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 5460 13240 5488 13268
rect 4479 13212 5488 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4304 13144 4353 13172
rect 4304 13132 4310 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 5258 13132 5264 13184
rect 5316 13172 5322 13184
rect 5810 13172 5816 13184
rect 5316 13144 5816 13172
rect 5316 13132 5322 13144
rect 5810 13132 5816 13144
rect 5868 13172 5874 13184
rect 6104 13172 6132 13271
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6748 13308 6776 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7282 13376 7288 13388
rect 6963 13348 7288 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 11440 13385 11468 13484
rect 13832 13456 13860 13484
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 14148 13484 14473 13512
rect 14148 13472 14154 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 14461 13475 14519 13481
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 16172 13484 16313 13512
rect 16172 13472 16178 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 16485 13515 16543 13521
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 16850 13512 16856 13524
rect 16531 13484 16856 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 17644 13484 17693 13512
rect 17644 13472 17650 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 17681 13475 17739 13481
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 23566 13512 23572 13524
rect 18564 13484 23572 13512
rect 18564 13472 18570 13484
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 23658 13472 23664 13524
rect 23716 13472 23722 13524
rect 26053 13515 26111 13521
rect 26053 13481 26065 13515
rect 26099 13512 26111 13515
rect 26234 13512 26240 13524
rect 26099 13484 26240 13512
rect 26099 13481 26111 13484
rect 26053 13475 26111 13481
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 12894 13444 12900 13456
rect 11900 13416 12900 13444
rect 11425 13379 11483 13385
rect 8588 13348 11284 13376
rect 6512 13280 6776 13308
rect 6512 13268 6518 13280
rect 7006 13268 7012 13320
rect 7064 13268 7070 13320
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7190 13308 7196 13320
rect 7147 13280 7196 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7116 13240 7144 13271
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7616 13280 7757 13308
rect 7616 13268 7622 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13308 7895 13311
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 7883 13280 8401 13308
rect 7883 13277 7895 13280
rect 7837 13271 7895 13277
rect 8389 13277 8401 13280
rect 8435 13308 8447 13311
rect 8478 13308 8484 13320
rect 8435 13280 8484 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8588 13317 8616 13348
rect 11256 13320 11284 13348
rect 11425 13345 11437 13379
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 8573 13271 8631 13277
rect 8680 13280 9597 13308
rect 8680 13240 8708 13280
rect 9585 13277 9597 13280
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 7116 13212 8708 13240
rect 7116 13172 7144 13212
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9364 13212 9413 13240
rect 9364 13200 9370 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9600 13240 9628 13271
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 9824 13280 10885 13308
rect 9824 13268 9830 13280
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11900 13308 11928 13416
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 13722 13444 13728 13456
rect 13464 13416 13728 13444
rect 13262 13376 13268 13388
rect 11992 13348 13268 13376
rect 11992 13317 12020 13348
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 11296 13280 11928 13308
rect 11977 13311 12035 13317
rect 11296 13268 11302 13280
rect 11977 13277 11989 13311
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 13464 13308 13492 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14642 13444 14648 13456
rect 13872 13416 14648 13444
rect 13872 13404 13878 13416
rect 14642 13404 14648 13416
rect 14700 13444 14706 13456
rect 15105 13447 15163 13453
rect 15105 13444 15117 13447
rect 14700 13416 15117 13444
rect 14700 13404 14706 13416
rect 15105 13413 15117 13416
rect 15151 13413 15163 13447
rect 15105 13407 15163 13413
rect 17954 13404 17960 13456
rect 18012 13444 18018 13456
rect 20070 13444 20076 13456
rect 18012 13416 20076 13444
rect 18012 13404 18018 13416
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 22738 13404 22744 13456
rect 22796 13444 22802 13456
rect 23753 13447 23811 13453
rect 23753 13444 23765 13447
rect 22796 13416 23765 13444
rect 22796 13404 22802 13416
rect 23753 13413 23765 13416
rect 23799 13413 23811 13447
rect 23753 13407 23811 13413
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 20254 13376 20260 13388
rect 15703 13348 20260 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 20254 13336 20260 13348
rect 20312 13336 20318 13388
rect 23952 13348 24808 13376
rect 14182 13308 14188 13320
rect 12115 13280 13492 13308
rect 13556 13280 14188 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 9600 13212 10272 13240
rect 9401 13203 9459 13209
rect 5868 13144 7144 13172
rect 5868 13132 5874 13144
rect 8478 13132 8484 13184
rect 8536 13132 8542 13184
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 9628 13172 9634 13184
rect 8628 13144 9634 13172
rect 8628 13132 8634 13144
rect 9628 13132 9634 13144
rect 9686 13132 9692 13184
rect 10244 13172 10272 13212
rect 10502 13200 10508 13252
rect 10560 13240 10566 13252
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 10560 13212 10609 13240
rect 10560 13200 10566 13212
rect 10597 13209 10609 13212
rect 10643 13209 10655 13243
rect 12161 13243 12219 13249
rect 12161 13240 12173 13243
rect 10597 13203 10655 13209
rect 10888 13212 12173 13240
rect 10888 13184 10916 13212
rect 12161 13209 12173 13212
rect 12207 13240 12219 13243
rect 13556 13240 13584 13280
rect 14182 13268 14188 13280
rect 14240 13308 14246 13320
rect 14826 13308 14832 13320
rect 14240 13280 14832 13308
rect 14240 13268 14246 13280
rect 14826 13268 14832 13280
rect 14884 13308 14890 13320
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 14884 13280 15301 13308
rect 14884 13268 14890 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16850 13308 16856 13320
rect 15804 13280 16856 13308
rect 15804 13268 15810 13280
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18138 13308 18144 13320
rect 18003 13280 18144 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18138 13268 18144 13280
rect 18196 13308 18202 13320
rect 19058 13308 19064 13320
rect 18196 13280 19064 13308
rect 18196 13268 18202 13280
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13308 19579 13311
rect 20346 13308 20352 13320
rect 19567 13280 20352 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 22002 13308 22008 13320
rect 21039 13280 22008 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 23566 13268 23572 13320
rect 23624 13268 23630 13320
rect 23658 13268 23664 13320
rect 23716 13308 23722 13320
rect 23952 13308 23980 13348
rect 23716 13280 23980 13308
rect 24029 13311 24087 13317
rect 23716 13268 23722 13280
rect 24029 13277 24041 13311
rect 24075 13308 24087 13311
rect 24486 13308 24492 13320
rect 24075 13280 24492 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 12207 13212 13584 13240
rect 14277 13243 14335 13249
rect 12207 13209 12219 13212
rect 12161 13203 12219 13209
rect 14277 13209 14289 13243
rect 14323 13209 14335 13243
rect 14277 13203 14335 13209
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10244 13144 10793 13172
rect 10781 13141 10793 13144
rect 10827 13141 10839 13175
rect 10781 13135 10839 13141
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 11606 13132 11612 13184
rect 11664 13132 11670 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 14292 13172 14320 13203
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 15381 13243 15439 13249
rect 15381 13240 15393 13243
rect 14792 13212 15393 13240
rect 14792 13200 14798 13212
rect 15381 13209 15393 13212
rect 15427 13209 15439 13243
rect 15381 13203 15439 13209
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 15620 13212 16129 13240
rect 15620 13200 15626 13212
rect 16117 13209 16129 13212
rect 16163 13209 16175 13243
rect 16117 13203 16175 13209
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 16540 13212 20029 13240
rect 16540 13200 16546 13212
rect 13412 13144 14320 13172
rect 13412 13132 13418 13144
rect 14458 13132 14464 13184
rect 14516 13181 14522 13184
rect 14516 13175 14535 13181
rect 14523 13141 14535 13175
rect 14516 13135 14535 13141
rect 14516 13132 14522 13135
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 15068 13144 15485 13172
rect 15068 13132 15074 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 16317 13175 16375 13181
rect 16317 13172 16329 13175
rect 16080 13144 16329 13172
rect 16080 13132 16086 13144
rect 16317 13141 16329 13144
rect 16363 13141 16375 13175
rect 16317 13135 16375 13141
rect 17218 13132 17224 13184
rect 17276 13132 17282 13184
rect 17865 13175 17923 13181
rect 17865 13141 17877 13175
rect 17911 13172 17923 13175
rect 18506 13172 18512 13184
rect 17911 13144 18512 13172
rect 17911 13141 17923 13144
rect 17865 13135 17923 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19242 13132 19248 13184
rect 19300 13172 19306 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19300 13144 19625 13172
rect 19300 13132 19306 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 20001 13172 20029 13212
rect 20806 13200 20812 13252
rect 20864 13240 20870 13252
rect 21238 13243 21296 13249
rect 21238 13240 21250 13243
rect 20864 13212 21250 13240
rect 20864 13200 20870 13212
rect 21238 13209 21250 13212
rect 21284 13209 21296 13243
rect 24044 13240 24072 13271
rect 24486 13268 24492 13280
rect 24544 13268 24550 13320
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24780 13308 24808 13348
rect 26418 13336 26424 13388
rect 26476 13376 26482 13388
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26476 13348 26525 13376
rect 26476 13336 26482 13348
rect 26513 13345 26525 13348
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 24780 13280 26464 13308
rect 24673 13271 24731 13277
rect 21238 13203 21296 13209
rect 22020 13212 24072 13240
rect 22020 13172 22048 13212
rect 24118 13200 24124 13252
rect 24176 13240 24182 13252
rect 24688 13240 24716 13271
rect 24762 13240 24768 13252
rect 24176 13212 24768 13240
rect 24176 13200 24182 13212
rect 24762 13200 24768 13212
rect 24820 13200 24826 13252
rect 24946 13249 24952 13252
rect 24940 13203 24952 13249
rect 24946 13200 24952 13203
rect 25004 13200 25010 13252
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 26436 13240 26464 13280
rect 26602 13240 26608 13252
rect 25096 13212 26004 13240
rect 26436 13212 26608 13240
rect 25096 13200 25102 13212
rect 20001 13144 22048 13172
rect 19613 13135 19671 13141
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 22738 13172 22744 13184
rect 22428 13144 22744 13172
rect 22428 13132 22434 13144
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 22830 13132 22836 13184
rect 22888 13172 22894 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22888 13144 23305 13172
rect 22888 13132 22894 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 23937 13175 23995 13181
rect 23937 13141 23949 13175
rect 23983 13172 23995 13175
rect 25866 13172 25872 13184
rect 23983 13144 25872 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 25976 13172 26004 13212
rect 26602 13200 26608 13212
rect 26660 13200 26666 13252
rect 26780 13243 26838 13249
rect 26780 13209 26792 13243
rect 26826 13240 26838 13243
rect 27798 13240 27804 13252
rect 26826 13212 27804 13240
rect 26826 13209 26838 13212
rect 26780 13203 26838 13209
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 27893 13175 27951 13181
rect 27893 13172 27905 13175
rect 25976 13144 27905 13172
rect 27893 13141 27905 13144
rect 27939 13141 27951 13175
rect 27893 13135 27951 13141
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5534 12968 5540 12980
rect 4755 12940 5540 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6086 12968 6092 12980
rect 5951 12940 6092 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 7650 12968 7656 12980
rect 6656 12940 7656 12968
rect 4522 12860 4528 12912
rect 4580 12900 4586 12912
rect 5074 12900 5080 12912
rect 4580 12872 5080 12900
rect 4580 12860 4586 12872
rect 4908 12841 4936 12872
rect 5074 12860 5080 12872
rect 5132 12900 5138 12912
rect 6656 12909 6684 12940
rect 7650 12928 7656 12940
rect 7708 12968 7714 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7708 12940 7941 12968
rect 7708 12928 7714 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 12158 12968 12164 12980
rect 9272 12940 12164 12968
rect 9272 12928 9278 12940
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13814 12968 13820 12980
rect 13127 12940 13820 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 14277 12971 14335 12977
rect 13955 12940 14228 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 6641 12903 6699 12909
rect 5132 12872 6132 12900
rect 5132 12860 5138 12872
rect 6104 12844 6132 12872
rect 6641 12869 6653 12903
rect 6687 12869 6699 12903
rect 6841 12903 6899 12909
rect 6841 12900 6853 12903
rect 6641 12863 6699 12869
rect 6840 12869 6853 12900
rect 6887 12869 6899 12903
rect 8662 12900 8668 12912
rect 6840 12863 6899 12869
rect 7668 12872 8668 12900
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 4304 12736 5181 12764
rect 4304 12724 4310 12736
rect 5169 12733 5181 12736
rect 5215 12764 5227 12767
rect 5644 12764 5672 12795
rect 6086 12792 6092 12844
rect 6144 12792 6150 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6546 12832 6552 12844
rect 6328 12804 6552 12832
rect 6328 12792 6334 12804
rect 6546 12792 6552 12804
rect 6604 12832 6610 12844
rect 6840 12832 6868 12863
rect 7668 12841 7696 12872
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 11020 12872 12541 12900
rect 11020 12860 11026 12872
rect 12529 12869 12541 12872
rect 12575 12869 12587 12903
rect 12529 12863 12587 12869
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 14093 12903 14151 12909
rect 14093 12900 14105 12903
rect 12768 12872 14105 12900
rect 12768 12860 12774 12872
rect 14093 12869 14105 12872
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 6604 12804 6868 12832
rect 7653 12835 7711 12841
rect 6604 12792 6610 12804
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 5215 12736 5672 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 5902 12724 5908 12776
rect 5960 12724 5966 12776
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8294 12764 8300 12776
rect 7975 12736 8300 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8294 12724 8300 12736
rect 8352 12764 8358 12776
rect 8478 12764 8484 12776
rect 8352 12736 8484 12764
rect 8352 12724 8358 12736
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 5736 12696 5764 12724
rect 6914 12696 6920 12708
rect 5736 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 8386 12696 8392 12708
rect 7791 12668 8392 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8588 12696 8616 12795
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9640 12804 9781 12832
rect 9640 12792 9646 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 12802 12832 12808 12844
rect 11664 12804 12808 12832
rect 11664 12792 11670 12804
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13722 12832 13728 12844
rect 13412 12804 13728 12832
rect 13412 12792 13418 12804
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 9916 12736 13001 12764
rect 9916 12724 9922 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 14016 12764 14044 12795
rect 12989 12727 13047 12733
rect 13096 12736 14044 12764
rect 10134 12696 10140 12708
rect 8588 12668 10140 12696
rect 10134 12656 10140 12668
rect 10192 12696 10198 12708
rect 12529 12699 12587 12705
rect 12529 12696 12541 12699
rect 10192 12668 12541 12696
rect 10192 12656 10198 12668
rect 12529 12665 12541 12668
rect 12575 12696 12587 12699
rect 12618 12696 12624 12708
rect 12575 12668 12624 12696
rect 12575 12665 12587 12668
rect 12529 12659 12587 12665
rect 12618 12656 12624 12668
rect 12676 12696 12682 12708
rect 13096 12696 13124 12736
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14200 12764 14228 12940
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 16482 12968 16488 12980
rect 14323 12940 16488 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 17644 12940 18153 12968
rect 17644 12928 17650 12940
rect 18141 12937 18153 12940
rect 18187 12937 18199 12971
rect 18141 12931 18199 12937
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18748 12940 18889 12968
rect 18748 12928 18754 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 21082 12968 21088 12980
rect 19300 12940 21088 12968
rect 19300 12928 19306 12940
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 25130 12968 25136 12980
rect 22296 12940 25136 12968
rect 15933 12903 15991 12909
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 16206 12900 16212 12912
rect 15979 12872 16212 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 17770 12900 17776 12912
rect 17604 12872 17776 12900
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 15838 12841 15844 12844
rect 15805 12835 15844 12841
rect 15805 12801 15817 12835
rect 15805 12795 15844 12801
rect 15838 12792 15844 12795
rect 15896 12792 15902 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 14148 12736 14228 12764
rect 14148 12724 14154 12736
rect 12676 12668 13124 12696
rect 12676 12656 12682 12668
rect 13446 12656 13452 12708
rect 13504 12696 13510 12708
rect 16040 12696 16068 12795
rect 16114 12792 16120 12844
rect 16172 12841 16178 12844
rect 16172 12832 16180 12841
rect 16172 12804 16217 12832
rect 16172 12795 16180 12804
rect 16172 12792 16178 12795
rect 16298 12792 16304 12844
rect 16356 12832 16362 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16356 12804 17049 12832
rect 16356 12792 16362 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17604 12832 17632 12872
rect 17770 12860 17776 12872
rect 17828 12860 17834 12912
rect 17989 12903 18047 12909
rect 17989 12869 18001 12903
rect 18035 12900 18047 12903
rect 18322 12900 18328 12912
rect 18035 12872 18328 12900
rect 18035 12869 18047 12872
rect 17989 12863 18047 12869
rect 18322 12860 18328 12872
rect 18380 12900 18386 12912
rect 19150 12900 19156 12912
rect 18380 12872 19156 12900
rect 18380 12860 18386 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19426 12860 19432 12912
rect 19484 12860 19490 12912
rect 20622 12900 20628 12912
rect 19628 12872 20628 12900
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 17604 12804 18705 12832
rect 16850 12724 16856 12776
rect 16908 12724 16914 12776
rect 17604 12696 17632 12804
rect 18693 12801 18705 12804
rect 18739 12832 18751 12835
rect 19628 12832 19656 12872
rect 20622 12860 20628 12872
rect 20680 12860 20686 12912
rect 18739 12804 19656 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 17920 12736 19533 12764
rect 17920 12724 17926 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 13504 12668 16068 12696
rect 16224 12668 17632 12696
rect 13504 12656 13510 12668
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5166 12628 5172 12640
rect 5123 12600 5172 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5166 12588 5172 12600
rect 5224 12628 5230 12640
rect 5721 12631 5779 12637
rect 5721 12628 5733 12631
rect 5224 12600 5733 12628
rect 5224 12588 5230 12600
rect 5721 12597 5733 12600
rect 5767 12597 5779 12631
rect 5721 12591 5779 12597
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6604 12600 6837 12628
rect 6604 12588 6610 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7190 12628 7196 12640
rect 7055 12600 7196 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 8478 12588 8484 12640
rect 8536 12588 8542 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12628 9919 12631
rect 11882 12628 11888 12640
rect 9907 12600 11888 12628
rect 9907 12597 9919 12600
rect 9861 12591 9919 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12628 13323 12631
rect 13630 12628 13636 12640
rect 13311 12600 13636 12628
rect 13311 12597 13323 12600
rect 13265 12591 13323 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 16224 12628 16252 12668
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 19150 12696 19156 12708
rect 17736 12668 19156 12696
rect 17736 12656 17742 12668
rect 19150 12656 19156 12668
rect 19208 12656 19214 12708
rect 19628 12696 19656 12804
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12832 19763 12835
rect 19886 12832 19892 12844
rect 19751 12804 19892 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 22296 12841 22324 12940
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 22649 12903 22707 12909
rect 22649 12869 22661 12903
rect 22695 12900 22707 12903
rect 24670 12900 24676 12912
rect 22695 12872 24676 12900
rect 22695 12869 22707 12872
rect 22649 12863 22707 12869
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 22428 12804 22473 12832
rect 22428 12792 22434 12804
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 22738 12792 22744 12844
rect 22796 12841 22802 12844
rect 22796 12832 22804 12841
rect 22796 12804 22841 12832
rect 22796 12795 22804 12804
rect 22796 12792 22802 12795
rect 24026 12792 24032 12844
rect 24084 12792 24090 12844
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 23569 12767 23627 12773
rect 23569 12764 23581 12767
rect 19444 12668 19656 12696
rect 19812 12736 23581 12764
rect 19444 12640 19472 12668
rect 13780 12600 16252 12628
rect 13780 12588 13786 12600
rect 16298 12588 16304 12640
rect 16356 12588 16362 12640
rect 17221 12631 17279 12637
rect 17221 12597 17233 12631
rect 17267 12628 17279 12631
rect 17586 12628 17592 12640
rect 17267 12600 17592 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17954 12588 17960 12640
rect 18012 12588 18018 12640
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 18322 12628 18328 12640
rect 18104 12600 18328 12628
rect 18104 12588 18110 12600
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 19426 12588 19432 12640
rect 19484 12588 19490 12640
rect 19705 12631 19763 12637
rect 19705 12597 19717 12631
rect 19751 12628 19763 12631
rect 19812 12628 19840 12736
rect 23569 12733 23581 12736
rect 23615 12733 23627 12767
rect 23569 12727 23627 12733
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 23937 12767 23995 12773
rect 23937 12764 23949 12767
rect 23716 12736 23949 12764
rect 23716 12724 23722 12736
rect 23937 12733 23949 12736
rect 23983 12733 23995 12767
rect 24136 12764 24164 12795
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 24854 12832 24860 12844
rect 24412 12804 24860 12832
rect 24412 12764 24440 12804
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25032 12835 25090 12841
rect 25032 12801 25044 12835
rect 25078 12832 25090 12835
rect 26878 12832 26884 12844
rect 25078 12804 26884 12832
rect 25078 12801 25090 12804
rect 25032 12795 25090 12801
rect 24136 12736 24440 12764
rect 23937 12727 23995 12733
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 23845 12699 23903 12705
rect 23845 12665 23857 12699
rect 23891 12696 23903 12699
rect 24578 12696 24584 12708
rect 23891 12668 24584 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 24578 12656 24584 12668
rect 24636 12656 24642 12708
rect 19751 12600 19840 12628
rect 19751 12597 19763 12600
rect 19705 12591 19763 12597
rect 19886 12588 19892 12640
rect 19944 12588 19950 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22925 12631 22983 12637
rect 22925 12628 22937 12631
rect 22336 12600 22937 12628
rect 22336 12588 22342 12600
rect 22925 12597 22937 12600
rect 22971 12597 22983 12631
rect 22925 12591 22983 12597
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 25792 12628 25820 12804
rect 26878 12792 26884 12804
rect 26936 12792 26942 12844
rect 23532 12600 25820 12628
rect 23532 12588 23538 12600
rect 26142 12588 26148 12640
rect 26200 12588 26206 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4246 12424 4252 12436
rect 4019 12396 4252 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5261 12427 5319 12433
rect 5261 12393 5273 12427
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 5166 12356 5172 12368
rect 4856 12328 5172 12356
rect 4856 12316 4862 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 5276 12356 5304 12387
rect 5442 12384 5448 12436
rect 5500 12384 5506 12436
rect 5994 12424 6000 12436
rect 5552 12396 6000 12424
rect 5552 12356 5580 12396
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 7098 12424 7104 12436
rect 6604 12396 7104 12424
rect 6604 12384 6610 12396
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7466 12384 7472 12436
rect 7524 12384 7530 12436
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 10962 12424 10968 12436
rect 10376 12396 10968 12424
rect 10376 12384 10382 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 11664 12396 12081 12424
rect 11664 12384 11670 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 14090 12424 14096 12436
rect 12069 12387 12127 12393
rect 12406 12396 14096 12424
rect 5276 12328 5580 12356
rect 9677 12359 9735 12365
rect 9677 12325 9689 12359
rect 9723 12356 9735 12359
rect 10870 12356 10876 12368
rect 9723 12328 10876 12356
rect 9723 12325 9735 12328
rect 9677 12319 9735 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11974 12356 11980 12368
rect 11296 12328 11980 12356
rect 11296 12316 11302 12328
rect 11974 12316 11980 12328
rect 12032 12316 12038 12368
rect 1854 12248 1860 12300
rect 1912 12248 1918 12300
rect 4982 12288 4988 12300
rect 4356 12260 4988 12288
rect 750 12180 756 12232
rect 808 12220 814 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 808 12192 1593 12220
rect 808 12180 814 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4028 12192 4169 12220
rect 4028 12180 4034 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4172 12084 4200 12183
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4356 12229 4384 12260
rect 4982 12248 4988 12260
rect 5040 12288 5046 12300
rect 7282 12288 7288 12300
rect 5040 12260 7288 12288
rect 5040 12248 5046 12260
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 4304 12192 4353 12220
rect 4304 12180 4310 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4706 12220 4712 12232
rect 4479 12192 4712 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12220 5319 12223
rect 5350 12220 5356 12232
rect 5307 12192 5356 12220
rect 5307 12189 5319 12192
rect 5261 12183 5319 12189
rect 4908 12152 4936 12183
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 6638 12220 6644 12232
rect 5552 12192 6644 12220
rect 5074 12152 5080 12164
rect 4908 12124 5080 12152
rect 5074 12112 5080 12124
rect 5132 12152 5138 12164
rect 5442 12152 5448 12164
rect 5132 12124 5448 12152
rect 5132 12112 5138 12124
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 5552 12084 5580 12192
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6748 12229 6776 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 8444 12260 8493 12288
rect 8444 12248 8450 12260
rect 8481 12257 8493 12260
rect 8527 12288 8539 12291
rect 9306 12288 9312 12300
rect 8527 12260 9312 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10686 12288 10692 12300
rect 10275 12260 10692 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 12406 12288 12434 12396
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 16758 12424 16764 12436
rect 16448 12396 16764 12424
rect 16448 12384 16454 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 17000 12396 17049 12424
rect 17000 12384 17006 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17037 12387 17095 12393
rect 17126 12384 17132 12436
rect 17184 12384 17190 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 20254 12424 20260 12436
rect 19659 12396 20260 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 21174 12424 21180 12436
rect 20456 12396 21180 12424
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 17494 12356 17500 12368
rect 16724 12328 17500 12356
rect 16724 12316 16730 12328
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 17920 12328 20300 12356
rect 17920 12316 17926 12328
rect 11900 12260 12434 12288
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 6454 12112 6460 12164
rect 6512 12152 6518 12164
rect 6840 12152 6868 12183
rect 6512 12124 6868 12152
rect 7024 12152 7052 12183
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7466 12220 7472 12232
rect 7156 12192 7472 12220
rect 7156 12180 7162 12192
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 7668 12152 7696 12183
rect 8294 12180 8300 12232
rect 8352 12180 8358 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8662 12220 8668 12232
rect 8619 12192 8668 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8662 12180 8668 12192
rect 8720 12220 8726 12232
rect 9766 12220 9772 12232
rect 8720 12192 9772 12220
rect 8720 12180 8726 12192
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 11146 12220 11152 12232
rect 10468 12192 11152 12220
rect 10468 12180 10474 12192
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11756 12192 11805 12220
rect 11756 12180 11762 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 7024 12124 7696 12152
rect 9677 12155 9735 12161
rect 6512 12112 6518 12124
rect 4172 12056 5580 12084
rect 6086 12044 6092 12096
rect 6144 12084 6150 12096
rect 7024 12084 7052 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 9858 12152 9864 12164
rect 9723 12124 9864 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 11900 12152 11928 12260
rect 16206 12248 16212 12300
rect 16264 12288 16270 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 16264 12260 18337 12288
rect 16264 12248 16270 12260
rect 18325 12257 18337 12260
rect 18371 12288 18383 12291
rect 19242 12288 19248 12300
rect 18371 12260 19248 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 20272 12297 20300 12328
rect 20257 12291 20315 12297
rect 20257 12257 20269 12291
rect 20303 12288 20315 12291
rect 20456 12288 20484 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 21542 12424 21548 12436
rect 21499 12396 21548 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 21542 12384 21548 12396
rect 21600 12424 21606 12436
rect 23382 12424 23388 12436
rect 21600 12396 23388 12424
rect 21600 12384 21606 12396
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23474 12384 23480 12436
rect 23532 12384 23538 12436
rect 23566 12384 23572 12436
rect 23624 12424 23630 12436
rect 23661 12427 23719 12433
rect 23661 12424 23673 12427
rect 23624 12396 23673 12424
rect 23624 12384 23630 12396
rect 23661 12393 23673 12396
rect 23707 12393 23719 12427
rect 23661 12387 23719 12393
rect 25406 12384 25412 12436
rect 25464 12424 25470 12436
rect 27338 12424 27344 12436
rect 25464 12396 27344 12424
rect 25464 12384 25470 12396
rect 27338 12384 27344 12396
rect 27396 12384 27402 12436
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12356 20683 12359
rect 22462 12356 22468 12368
rect 20671 12328 22468 12356
rect 20671 12325 20683 12328
rect 20625 12319 20683 12325
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 20303 12260 20484 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 21284 12260 23428 12288
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 17184 12192 17233 12220
rect 17184 12180 17190 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 17402 12180 17408 12232
rect 17460 12180 17466 12232
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17678 12220 17684 12232
rect 17543 12192 17684 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 14544 12155 14602 12161
rect 10008 12124 12020 12152
rect 10008 12112 10014 12124
rect 11992 12096 12020 12124
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 16482 12152 16488 12164
rect 14590 12124 16488 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17420 12152 17448 12180
rect 17586 12152 17592 12164
rect 17000 12124 17592 12152
rect 17000 12112 17006 12124
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 18064 12152 18092 12183
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 18196 12192 20453 12220
rect 18196 12180 18202 12192
rect 19659 12189 19717 12192
rect 18598 12152 18604 12164
rect 18064 12124 18604 12152
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 19429 12155 19487 12161
rect 19429 12121 19441 12155
rect 19475 12152 19487 12155
rect 19518 12152 19524 12164
rect 19475 12124 19524 12152
rect 19475 12121 19487 12124
rect 19429 12115 19487 12121
rect 19518 12112 19524 12124
rect 19576 12112 19582 12164
rect 19659 12155 19671 12189
rect 19705 12155 19717 12189
rect 20441 12189 20453 12192
rect 20487 12220 20499 12223
rect 20990 12220 20996 12232
rect 20487 12192 20996 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21284 12229 21312 12260
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21232 12192 21281 12220
rect 21232 12180 21238 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 22189 12223 22247 12229
rect 22189 12220 22201 12223
rect 21269 12183 21327 12189
rect 22066 12192 22201 12220
rect 19659 12149 19717 12155
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 22066 12152 22094 12192
rect 22189 12189 22201 12192
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 22337 12223 22395 12229
rect 22337 12189 22349 12223
rect 22383 12220 22395 12223
rect 22383 12189 22416 12220
rect 22337 12183 22416 12189
rect 20220 12124 22094 12152
rect 22388 12152 22416 12183
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 22554 12180 22560 12232
rect 22612 12180 22618 12232
rect 22646 12180 22652 12232
rect 22704 12229 22710 12232
rect 22704 12220 22712 12229
rect 22704 12192 22749 12220
rect 22704 12183 22712 12192
rect 22704 12180 22710 12183
rect 22388 12124 22968 12152
rect 20220 12112 20226 12124
rect 6144 12056 7052 12084
rect 6144 12044 6150 12056
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 7156 12056 8125 12084
rect 7156 12044 7162 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10318 12084 10324 12096
rect 10192 12056 10324 12084
rect 10192 12044 10198 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10413 12087 10471 12093
rect 10413 12053 10425 12087
rect 10459 12084 10471 12087
rect 11146 12084 11152 12096
rect 10459 12056 11152 12084
rect 10459 12053 10471 12056
rect 10413 12047 10471 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11974 12044 11980 12096
rect 12032 12044 12038 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15344 12056 15669 12084
rect 15344 12044 15350 12056
rect 15657 12053 15669 12056
rect 15703 12053 15715 12087
rect 15657 12047 15715 12053
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 16724 12056 16773 12084
rect 16724 12044 16730 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 16761 12047 16819 12053
rect 17402 12044 17408 12096
rect 17460 12044 17466 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 18748 12056 19809 12084
rect 18748 12044 18754 12056
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 19797 12047 19855 12053
rect 22278 12044 22284 12096
rect 22336 12084 22342 12096
rect 22833 12087 22891 12093
rect 22833 12084 22845 12087
rect 22336 12056 22845 12084
rect 22336 12044 22342 12056
rect 22833 12053 22845 12056
rect 22879 12053 22891 12087
rect 22940 12084 22968 12124
rect 23014 12112 23020 12164
rect 23072 12152 23078 12164
rect 23290 12152 23296 12164
rect 23072 12124 23296 12152
rect 23072 12112 23078 12124
rect 23290 12112 23296 12124
rect 23348 12112 23354 12164
rect 23400 12152 23428 12260
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 25133 12223 25191 12229
rect 25133 12220 25145 12223
rect 24820 12192 25145 12220
rect 24820 12180 24826 12192
rect 25133 12189 25145 12192
rect 25179 12220 25191 12223
rect 26973 12223 27031 12229
rect 26973 12220 26985 12223
rect 25179 12192 26985 12220
rect 25179 12189 25191 12192
rect 25133 12183 25191 12189
rect 26973 12189 26985 12192
rect 27019 12189 27031 12223
rect 26973 12183 27031 12189
rect 28350 12180 28356 12232
rect 28408 12180 28414 12232
rect 25406 12161 25412 12164
rect 23493 12155 23551 12161
rect 23493 12152 23505 12155
rect 23400 12124 23505 12152
rect 23493 12121 23505 12124
rect 23539 12121 23551 12155
rect 23493 12115 23551 12121
rect 25400 12115 25412 12161
rect 25406 12112 25412 12115
rect 25464 12112 25470 12164
rect 25498 12112 25504 12164
rect 25556 12152 25562 12164
rect 27218 12155 27276 12161
rect 27218 12152 27230 12155
rect 25556 12124 27230 12152
rect 25556 12112 25562 12124
rect 27218 12121 27230 12124
rect 27264 12152 27276 12155
rect 28368 12152 28396 12180
rect 27264 12124 28396 12152
rect 27264 12121 27276 12124
rect 27218 12115 27276 12121
rect 25590 12084 25596 12096
rect 22940 12056 25596 12084
rect 22833 12047 22891 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 26510 12044 26516 12096
rect 26568 12044 26574 12096
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 28353 12087 28411 12093
rect 28353 12084 28365 12087
rect 26660 12056 28365 12084
rect 26660 12044 26666 12056
rect 28353 12053 28365 12056
rect 28399 12053 28411 12087
rect 28353 12047 28411 12053
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 5997 11883 6055 11889
rect 2746 11852 5948 11880
rect 1762 11568 1768 11620
rect 1820 11608 1826 11620
rect 2746 11608 2774 11852
rect 4249 11815 4307 11821
rect 4249 11781 4261 11815
rect 4295 11812 4307 11815
rect 4338 11812 4344 11824
rect 4295 11784 4344 11812
rect 4295 11781 4307 11784
rect 4249 11775 4307 11781
rect 4338 11772 4344 11784
rect 4396 11772 4402 11824
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5442 11744 5448 11756
rect 5215 11716 5448 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 3896 11676 3924 11707
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 5920 11744 5948 11852
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6178 11880 6184 11892
rect 6043 11852 6184 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6914 11840 6920 11892
rect 6972 11840 6978 11892
rect 8205 11883 8263 11889
rect 8205 11849 8217 11883
rect 8251 11880 8263 11883
rect 10134 11880 10140 11892
rect 8251 11852 10140 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 11756 11852 14136 11880
rect 11756 11840 11762 11852
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 6512 11784 6561 11812
rect 6512 11772 6518 11784
rect 6549 11781 6561 11784
rect 6595 11781 6607 11815
rect 6549 11775 6607 11781
rect 6730 11772 6736 11824
rect 6788 11772 6794 11824
rect 9760 11815 9818 11821
rect 9760 11781 9772 11815
rect 9806 11812 9818 11815
rect 14108 11812 14136 11852
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14734 11880 14740 11892
rect 14240 11852 14740 11880
rect 14240 11840 14246 11852
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 19426 11880 19432 11892
rect 15611 11852 19432 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19644 11852 20029 11880
rect 9806 11784 12112 11812
rect 14108 11784 14412 11812
rect 9806 11781 9818 11784
rect 9760 11775 9818 11781
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5920 11716 6009 11744
rect 5997 11713 6009 11716
rect 6043 11744 6055 11747
rect 7558 11744 7564 11756
rect 6043 11716 7564 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 7558 11704 7564 11716
rect 7616 11744 7622 11756
rect 8297 11747 8355 11753
rect 7616 11716 8156 11744
rect 7616 11704 7622 11716
rect 4246 11676 4252 11688
rect 3896 11648 4252 11676
rect 4246 11636 4252 11648
rect 4304 11676 4310 11688
rect 4890 11676 4896 11688
rect 4304 11648 4896 11676
rect 4304 11636 4310 11648
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 4982 11636 4988 11688
rect 5040 11636 5046 11688
rect 5074 11636 5080 11688
rect 5132 11636 5138 11688
rect 5258 11636 5264 11688
rect 5316 11636 5322 11688
rect 8128 11676 8156 11716
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 9398 11744 9404 11756
rect 8343 11716 9404 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 10318 11744 10324 11756
rect 9539 11716 10324 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 11957 11747 12015 11753
rect 11957 11744 11969 11747
rect 11848 11716 11969 11744
rect 11848 11704 11854 11716
rect 11957 11713 11969 11716
rect 12003 11713 12015 11747
rect 12084 11744 12112 11784
rect 14090 11744 14096 11756
rect 12084 11716 14096 11744
rect 11957 11707 12015 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14384 11753 14412 11784
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 16206 11812 16212 11824
rect 15252 11784 16212 11812
rect 15252 11772 15258 11784
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 18966 11812 18972 11824
rect 16776 11784 18972 11812
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14826 11744 14832 11756
rect 14415 11716 14832 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8128 11648 8401 11676
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 1820 11580 2774 11608
rect 1820 11568 1826 11580
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 4764 11580 4936 11608
rect 4764 11568 4770 11580
rect 4908 11552 4936 11580
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 6546 11608 6552 11620
rect 5776 11580 6552 11608
rect 5776 11568 5782 11580
rect 6546 11568 6552 11580
rect 6604 11608 6610 11620
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 6604 11580 7849 11608
rect 6604 11568 6610 11580
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7837 11571 7895 11577
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3970 11540 3976 11552
rect 3476 11512 3976 11540
rect 3476 11500 3482 11512
rect 3970 11500 3976 11512
rect 4028 11540 4034 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4028 11512 4813 11540
rect 4028 11500 4034 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 7558 11540 7564 11552
rect 4948 11512 7564 11540
rect 4948 11500 4954 11512
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8404 11540 8432 11639
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 10744 11648 11713 11676
rect 10744 11636 10750 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 14200 11676 14228 11707
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15286 11704 15292 11756
rect 15344 11704 15350 11756
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11744 15439 11747
rect 15654 11744 15660 11756
rect 15427 11716 15660 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 15654 11704 15660 11716
rect 15712 11744 15718 11756
rect 16776 11744 16804 11784
rect 18966 11772 18972 11784
rect 19024 11772 19030 11824
rect 19058 11772 19064 11824
rect 19116 11812 19122 11824
rect 19644 11812 19672 11852
rect 19116 11784 19672 11812
rect 19116 11772 19122 11784
rect 19702 11772 19708 11824
rect 19760 11812 19766 11824
rect 19889 11815 19947 11821
rect 19889 11812 19901 11815
rect 19760 11784 19901 11812
rect 19760 11772 19766 11784
rect 19889 11781 19901 11784
rect 19935 11781 19947 11815
rect 19889 11775 19947 11781
rect 15712 11716 16804 11744
rect 15712 11704 15718 11716
rect 16850 11704 16856 11756
rect 16908 11704 16914 11756
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17954 11753 17960 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17552 11716 17693 11744
rect 17552 11704 17558 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17948 11744 17960 11753
rect 17915 11716 17960 11744
rect 17681 11707 17739 11713
rect 17948 11707 17960 11716
rect 17954 11704 17960 11707
rect 18012 11704 18018 11756
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 15930 11676 15936 11688
rect 13964 11648 15936 11676
rect 13964 11636 13970 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16540 11648 17264 11676
rect 16540 11636 16546 11648
rect 14461 11611 14519 11617
rect 14461 11577 14473 11611
rect 14507 11577 14519 11611
rect 14461 11571 14519 11577
rect 9214 11540 9220 11552
rect 8404 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11540 9278 11552
rect 9858 11540 9864 11552
rect 9272 11512 9864 11540
rect 9272 11500 9278 11512
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10836 11512 10885 11540
rect 10836 11500 10842 11512
rect 10873 11509 10885 11512
rect 10919 11540 10931 11543
rect 11238 11540 11244 11552
rect 10919 11512 11244 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13078 11540 13084 11552
rect 12860 11512 13084 11540
rect 12860 11500 12866 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 14476 11540 14504 11571
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 17126 11608 17132 11620
rect 14976 11580 17132 11608
rect 14976 11568 14982 11580
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 17236 11608 17264 11648
rect 19536 11608 19564 11707
rect 19610 11704 19616 11756
rect 19668 11744 19674 11756
rect 20001 11753 20029 11852
rect 21082 11840 21088 11892
rect 21140 11840 21146 11892
rect 22646 11840 22652 11892
rect 22704 11880 22710 11892
rect 23014 11880 23020 11892
rect 22704 11852 23020 11880
rect 22704 11840 22710 11852
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 24210 11880 24216 11892
rect 23624 11852 24216 11880
rect 23624 11840 23630 11852
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 25038 11840 25044 11892
rect 25096 11840 25102 11892
rect 26602 11880 26608 11892
rect 25148 11852 26608 11880
rect 20530 11812 20536 11824
rect 20180 11784 20536 11812
rect 19797 11747 19855 11753
rect 19668 11716 19713 11744
rect 19668 11704 19674 11716
rect 19797 11713 19809 11747
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 19986 11747 20044 11753
rect 19986 11713 19998 11747
rect 20032 11713 20044 11747
rect 19986 11707 20044 11713
rect 19812 11676 19840 11707
rect 20180 11688 20208 11784
rect 20530 11772 20536 11784
rect 20588 11772 20594 11824
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 21100 11753 21128 11840
rect 22554 11812 22560 11824
rect 22020 11784 22560 11812
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20312 11716 21097 11744
rect 20312 11704 20318 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21450 11744 21456 11756
rect 21315 11716 21456 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 20162 11676 20168 11688
rect 19812 11648 20168 11676
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20346 11636 20352 11688
rect 20404 11676 20410 11688
rect 22020 11676 22048 11784
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 22738 11772 22744 11824
rect 22796 11812 22802 11824
rect 22833 11815 22891 11821
rect 22833 11812 22845 11815
rect 22796 11784 22845 11812
rect 22796 11772 22802 11784
rect 22833 11781 22845 11784
rect 22879 11781 22891 11815
rect 22833 11775 22891 11781
rect 22925 11815 22983 11821
rect 22925 11781 22937 11815
rect 22971 11812 22983 11815
rect 22971 11784 23704 11812
rect 22971 11781 22983 11784
rect 22925 11775 22983 11781
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 22649 11747 22707 11753
rect 22649 11744 22661 11747
rect 22244 11716 22661 11744
rect 22244 11704 22250 11716
rect 22649 11713 22661 11716
rect 22695 11713 22707 11747
rect 22649 11707 22707 11713
rect 23014 11704 23020 11756
rect 23072 11704 23078 11756
rect 23566 11704 23572 11756
rect 23624 11704 23630 11756
rect 23676 11744 23704 11784
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 23928 11815 23986 11821
rect 23928 11812 23940 11815
rect 23808 11784 23940 11812
rect 23808 11772 23814 11784
rect 23928 11781 23940 11784
rect 23974 11812 23986 11815
rect 25148 11812 25176 11852
rect 26602 11840 26608 11852
rect 26660 11840 26666 11892
rect 27154 11840 27160 11892
rect 27212 11840 27218 11892
rect 25590 11812 25596 11824
rect 23974 11784 25176 11812
rect 25424 11784 25596 11812
rect 23974 11781 23986 11784
rect 23928 11775 23986 11781
rect 25424 11744 25452 11784
rect 25590 11772 25596 11784
rect 25648 11772 25654 11824
rect 25777 11815 25835 11821
rect 25777 11781 25789 11815
rect 25823 11812 25835 11815
rect 26786 11812 26792 11824
rect 25823 11784 26792 11812
rect 25823 11781 25835 11784
rect 25777 11775 25835 11781
rect 26786 11772 26792 11784
rect 26844 11772 26850 11824
rect 26878 11772 26884 11824
rect 26936 11812 26942 11824
rect 27172 11812 27200 11840
rect 27433 11815 27491 11821
rect 27433 11812 27445 11815
rect 26936 11784 27445 11812
rect 26936 11772 26942 11784
rect 27433 11781 27445 11784
rect 27479 11781 27491 11815
rect 27433 11775 27491 11781
rect 23676 11716 25452 11744
rect 25498 11704 25504 11756
rect 25556 11704 25562 11756
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 25869 11747 25927 11753
rect 25869 11713 25881 11747
rect 25915 11744 25927 11747
rect 26142 11744 26148 11756
rect 25915 11716 26148 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 20404 11648 22048 11676
rect 20404 11636 20410 11648
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 23584 11676 23612 11704
rect 22152 11648 23612 11676
rect 22152 11636 22158 11648
rect 23658 11636 23664 11688
rect 23716 11636 23722 11688
rect 24762 11636 24768 11688
rect 24820 11676 24826 11688
rect 25700 11676 25728 11707
rect 26142 11704 26148 11716
rect 26200 11704 26206 11756
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 27246 11744 27252 11756
rect 27203 11716 27252 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 27246 11704 27252 11716
rect 27304 11704 27310 11756
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11713 27399 11747
rect 27341 11707 27399 11713
rect 26326 11676 26332 11688
rect 24820 11648 26332 11676
rect 24820 11636 24826 11648
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27062 11636 27068 11688
rect 27120 11676 27126 11688
rect 27356 11676 27384 11707
rect 27522 11704 27528 11756
rect 27580 11704 27586 11756
rect 27120 11648 27384 11676
rect 27120 11636 27126 11648
rect 23566 11608 23572 11620
rect 17236 11580 17632 11608
rect 19536 11580 23572 11608
rect 16942 11540 16948 11552
rect 14476 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 17494 11540 17500 11552
rect 17083 11512 17500 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 17604 11540 17632 11580
rect 23566 11568 23572 11580
rect 23624 11568 23630 11620
rect 17862 11540 17868 11552
rect 17604 11512 17868 11540
rect 17862 11500 17868 11512
rect 17920 11540 17926 11552
rect 19061 11543 19119 11549
rect 19061 11540 19073 11543
rect 17920 11512 19073 11540
rect 17920 11500 17926 11512
rect 19061 11509 19073 11512
rect 19107 11509 19119 11543
rect 19061 11503 19119 11509
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 20165 11543 20223 11549
rect 20165 11540 20177 11543
rect 19760 11512 20177 11540
rect 19760 11500 19766 11512
rect 20165 11509 20177 11512
rect 20211 11509 20223 11543
rect 20165 11503 20223 11509
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 22646 11500 22652 11552
rect 22704 11540 22710 11552
rect 23201 11543 23259 11549
rect 23201 11540 23213 11543
rect 22704 11512 23213 11540
rect 22704 11500 22710 11512
rect 23201 11509 23213 11512
rect 23247 11509 23259 11543
rect 23201 11503 23259 11509
rect 23382 11500 23388 11552
rect 23440 11540 23446 11552
rect 26053 11543 26111 11549
rect 26053 11540 26065 11543
rect 23440 11512 26065 11540
rect 23440 11500 23446 11512
rect 26053 11509 26065 11512
rect 26099 11509 26111 11543
rect 26053 11503 26111 11509
rect 27706 11500 27712 11552
rect 27764 11500 27770 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 4154 11336 4160 11348
rect 4111 11308 4160 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 4154 11296 4160 11308
rect 4212 11336 4218 11348
rect 5166 11336 5172 11348
rect 4212 11308 5172 11336
rect 4212 11296 4218 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 5316 11308 5917 11336
rect 5316 11296 5322 11308
rect 5905 11305 5917 11308
rect 5951 11305 5963 11339
rect 5905 11299 5963 11305
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6420 11308 6837 11336
rect 6420 11296 6426 11308
rect 6825 11305 6837 11308
rect 6871 11336 6883 11339
rect 9582 11336 9588 11348
rect 6871 11308 9588 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9858 11296 9864 11348
rect 9916 11296 9922 11348
rect 10686 11336 10692 11348
rect 9968 11308 10692 11336
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 4617 11271 4675 11277
rect 4617 11268 4629 11271
rect 4396 11240 4629 11268
rect 4396 11228 4402 11240
rect 4617 11237 4629 11240
rect 4663 11268 4675 11271
rect 5442 11268 5448 11280
rect 4663 11240 5448 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 6086 11228 6092 11280
rect 6144 11268 6150 11280
rect 7009 11271 7067 11277
rect 7009 11268 7021 11271
rect 6144 11240 7021 11268
rect 6144 11228 6150 11240
rect 7009 11237 7021 11240
rect 7055 11237 7067 11271
rect 7009 11231 7067 11237
rect 7558 11228 7564 11280
rect 7616 11268 7622 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 7616 11240 7665 11268
rect 7616 11228 7622 11240
rect 7653 11237 7665 11240
rect 7699 11237 7711 11271
rect 7653 11231 7711 11237
rect 9309 11271 9367 11277
rect 9309 11237 9321 11271
rect 9355 11237 9367 11271
rect 9309 11231 9367 11237
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 7098 11200 7104 11212
rect 5399 11172 6132 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 4154 11092 4160 11144
rect 4212 11141 4218 11144
rect 4212 11135 4245 11141
rect 4233 11101 4245 11135
rect 4212 11095 4245 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 4212 11092 4218 11095
rect 3510 11024 3516 11076
rect 3568 11064 3574 11076
rect 4724 11064 4752 11095
rect 5258 11092 5264 11144
rect 5316 11092 5322 11144
rect 6104 11141 6132 11172
rect 6288 11172 7104 11200
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 6089 11135 6147 11141
rect 5491 11104 6040 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5810 11064 5816 11076
rect 3568 11036 4292 11064
rect 4724 11036 5816 11064
rect 3568 11024 3574 11036
rect 4264 11005 4292 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 5905 11067 5963 11073
rect 5905 11033 5917 11067
rect 5951 11033 5963 11067
rect 6012 11064 6040 11104
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6178 11092 6184 11144
rect 6236 11092 6242 11144
rect 6288 11064 6316 11172
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 9324 11200 9352 11231
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 9968 11268 9996 11308
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 12342 11336 12348 11348
rect 11204 11308 12348 11336
rect 11204 11296 11210 11308
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 15194 11336 15200 11348
rect 13504 11308 15200 11336
rect 13504 11296 13510 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 15933 11339 15991 11345
rect 15933 11305 15945 11339
rect 15979 11336 15991 11339
rect 18230 11336 18236 11348
rect 15979 11308 18236 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 9548 11240 9996 11268
rect 11793 11271 11851 11277
rect 9548 11228 9554 11240
rect 11793 11237 11805 11271
rect 11839 11268 11851 11271
rect 12250 11268 12256 11280
rect 11839 11240 12256 11268
rect 11839 11237 11851 11240
rect 11793 11231 11851 11237
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 15764 11268 15792 11299
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20622 11336 20628 11348
rect 20395 11308 20628 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 23014 11296 23020 11348
rect 23072 11336 23078 11348
rect 25038 11336 25044 11348
rect 23072 11308 25044 11336
rect 23072 11296 23078 11308
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 25130 11296 25136 11348
rect 25188 11296 25194 11348
rect 17218 11268 17224 11280
rect 15764 11240 17224 11268
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18877 11271 18935 11277
rect 18877 11237 18889 11271
rect 18923 11268 18935 11271
rect 18966 11268 18972 11280
rect 18923 11240 18972 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 20070 11228 20076 11280
rect 20128 11268 20134 11280
rect 20438 11268 20444 11280
rect 20128 11240 20444 11268
rect 20128 11228 20134 11240
rect 20438 11228 20444 11240
rect 20496 11228 20502 11280
rect 22186 11268 22192 11280
rect 21192 11240 22192 11268
rect 9508 11200 9536 11228
rect 7524 11172 9352 11200
rect 9416 11172 9536 11200
rect 7524 11160 7530 11172
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6012 11036 6316 11064
rect 6656 11064 6684 11095
rect 6822 11092 6828 11144
rect 6880 11092 6886 11144
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 9416 11132 9444 11172
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10410 11160 10416 11212
rect 10468 11160 10474 11212
rect 15286 11200 15292 11212
rect 14752 11172 15292 11200
rect 8996 11104 9444 11132
rect 9491 11135 9549 11141
rect 8996 11092 9002 11104
rect 9491 11101 9503 11135
rect 9537 11132 9549 11135
rect 10680 11135 10738 11141
rect 9537 11104 9904 11132
rect 9537 11101 9549 11104
rect 9491 11095 9549 11101
rect 6914 11064 6920 11076
rect 6656 11036 6920 11064
rect 5905 11027 5963 11033
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10965 4307 10999
rect 4249 10959 4307 10965
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 5920 10996 5948 11027
rect 6914 11024 6920 11036
rect 6972 11064 6978 11076
rect 7190 11064 7196 11076
rect 6972 11036 7196 11064
rect 6972 11024 6978 11036
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7340 11036 7941 11064
rect 7340 11024 7346 11036
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 9030 11064 9036 11076
rect 8260 11036 9036 11064
rect 8260 11024 8266 11036
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9876 11064 9904 11104
rect 10680 11101 10692 11135
rect 10726 11132 10738 11135
rect 14090 11132 14096 11144
rect 10726 11104 14096 11132
rect 10726 11101 10738 11104
rect 10680 11095 10738 11101
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14752 11141 14780 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 17310 11200 17316 11212
rect 15703 11172 17316 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17494 11160 17500 11212
rect 17552 11160 17558 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 19576 11172 19993 11200
rect 19576 11160 19582 11172
rect 19904 11144 19932 11172
rect 19981 11169 19993 11172
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15436 11104 15761 11132
rect 15436 11092 15442 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16264 11104 16681 11132
rect 16264 11092 16270 11104
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 16758 11092 16764 11144
rect 16816 11092 16822 11144
rect 16942 11092 16948 11144
rect 17000 11092 17006 11144
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11132 17095 11135
rect 17126 11132 17132 11144
rect 17083 11104 17132 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17764 11135 17822 11141
rect 17764 11132 17776 11135
rect 17696 11104 17776 11132
rect 9232 11036 9628 11064
rect 9876 11036 15148 11064
rect 5500 10968 5948 10996
rect 8113 10999 8171 11005
rect 5500 10956 5506 10968
rect 8113 10965 8125 10999
rect 8159 10996 8171 10999
rect 8570 10996 8576 11008
rect 8159 10968 8576 10996
rect 8159 10965 8171 10968
rect 8113 10959 8171 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 9232 10996 9260 11036
rect 8812 10968 9260 10996
rect 8812 10956 8818 10968
rect 9490 10956 9496 11008
rect 9548 10956 9554 11008
rect 9600 10996 9628 11036
rect 10318 10996 10324 11008
rect 9600 10968 10324 10996
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 11146 10996 11152 11008
rect 10468 10968 11152 10996
rect 10468 10956 10474 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 15120 10996 15148 11036
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 16485 11067 16543 11073
rect 16485 11033 16497 11067
rect 16531 11064 16543 11067
rect 17310 11064 17316 11076
rect 16531 11036 17316 11064
rect 16531 11033 16543 11036
rect 16485 11027 16543 11033
rect 17310 11024 17316 11036
rect 17368 11024 17374 11076
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 17696 11064 17724 11104
rect 17764 11101 17776 11104
rect 17810 11101 17822 11135
rect 17764 11095 17822 11101
rect 19886 11092 19892 11144
rect 19944 11092 19950 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 19996 11104 20177 11132
rect 19996 11076 20024 11104
rect 20165 11101 20177 11104
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 20772 11104 20913 11132
rect 20772 11092 20778 11104
rect 20901 11101 20913 11104
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 21082 11092 21088 11144
rect 21140 11092 21146 11144
rect 21192 11141 21220 11240
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 22554 11228 22560 11280
rect 22612 11268 22618 11280
rect 22612 11240 23152 11268
rect 22612 11228 22618 11240
rect 21358 11200 21364 11212
rect 21284 11172 21364 11200
rect 21284 11141 21312 11172
rect 21358 11160 21364 11172
rect 21416 11160 21422 11212
rect 21545 11203 21603 11209
rect 21545 11169 21557 11203
rect 21591 11200 21603 11203
rect 23014 11200 23020 11212
rect 21591 11172 23020 11200
rect 21591 11169 21603 11172
rect 21545 11163 21603 11169
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 23124 11200 23152 11240
rect 23658 11228 23664 11280
rect 23716 11268 23722 11280
rect 24029 11271 24087 11277
rect 24029 11268 24041 11271
rect 23716 11240 24041 11268
rect 23716 11228 23722 11240
rect 24029 11237 24041 11240
rect 24075 11268 24087 11271
rect 24854 11268 24860 11280
rect 24075 11240 24860 11268
rect 24075 11237 24087 11240
rect 24029 11231 24087 11237
rect 24854 11228 24860 11240
rect 24912 11228 24918 11280
rect 24946 11228 24952 11280
rect 25004 11268 25010 11280
rect 25958 11268 25964 11280
rect 25004 11240 25964 11268
rect 25004 11228 25010 11240
rect 25958 11228 25964 11240
rect 26016 11228 26022 11280
rect 27338 11228 27344 11280
rect 27396 11228 27402 11280
rect 23124 11172 23198 11200
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 22830 11141 22836 11144
rect 22797 11135 22836 11141
rect 22797 11101 22809 11135
rect 22797 11095 22836 11101
rect 22830 11092 22836 11095
rect 22888 11092 22894 11144
rect 23170 11141 23198 11172
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 24872 11200 24900 11228
rect 23348 11172 23520 11200
rect 24872 11172 25075 11200
rect 23348 11160 23354 11172
rect 23153 11135 23211 11141
rect 23153 11101 23165 11135
rect 23199 11101 23211 11135
rect 23492 11132 23520 11172
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23492 11104 23857 11132
rect 23153 11095 23211 11101
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 17460 11036 17724 11064
rect 17460 11024 17466 11036
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 18690 11064 18696 11076
rect 18196 11036 18696 11064
rect 18196 11024 18202 11036
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 18874 11024 18880 11076
rect 18932 11064 18938 11076
rect 19978 11064 19984 11076
rect 18932 11036 19984 11064
rect 18932 11024 18938 11036
rect 19978 11024 19984 11036
rect 20036 11024 20042 11076
rect 21450 11073 21456 11076
rect 21407 11067 21456 11073
rect 21407 11033 21419 11067
rect 21453 11033 21456 11067
rect 21407 11027 21456 11033
rect 21450 11024 21456 11027
rect 21508 11024 21514 11076
rect 22370 11024 22376 11076
rect 22428 11064 22434 11076
rect 22925 11067 22983 11073
rect 22925 11064 22937 11067
rect 22428 11036 22937 11064
rect 22428 11024 22434 11036
rect 22925 11033 22937 11036
rect 22971 11033 22983 11067
rect 22925 11027 22983 11033
rect 23017 11067 23075 11073
rect 23017 11033 23029 11067
rect 23063 11064 23075 11067
rect 24026 11064 24032 11076
rect 23063 11036 24032 11064
rect 23063 11033 23075 11036
rect 23017 11027 23075 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 24596 11064 24624 11095
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 25047 11132 25075 11172
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25280 11172 26096 11200
rect 25280 11160 25286 11172
rect 25961 11135 26019 11141
rect 25961 11132 25973 11135
rect 25047 11104 25973 11132
rect 25961 11101 25973 11104
rect 26007 11101 26019 11135
rect 26068 11132 26096 11172
rect 26217 11135 26275 11141
rect 26217 11132 26229 11135
rect 26068 11104 26229 11132
rect 25961 11095 26019 11101
rect 26217 11101 26229 11104
rect 26263 11101 26275 11135
rect 26217 11095 26275 11101
rect 24688 11064 24716 11092
rect 24596 11036 24716 11064
rect 24857 11067 24915 11073
rect 24857 11033 24869 11067
rect 24903 11064 24915 11067
rect 26050 11064 26056 11076
rect 24903 11036 26056 11064
rect 24903 11033 24915 11036
rect 24857 11027 24915 11033
rect 26050 11024 26056 11036
rect 26108 11024 26114 11076
rect 16206 10996 16212 11008
rect 15120 10968 16212 10996
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17494 10996 17500 11008
rect 16908 10968 17500 10996
rect 16908 10956 16914 10968
rect 17494 10956 17500 10968
rect 17552 10996 17558 11008
rect 20070 10996 20076 11008
rect 17552 10968 20076 10996
rect 17552 10956 17558 10968
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 23290 10956 23296 11008
rect 23348 10956 23354 11008
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 24486 10996 24492 11008
rect 24360 10968 24492 10996
rect 24360 10956 24366 10968
rect 24486 10956 24492 10968
rect 24544 10996 24550 11008
rect 24946 10996 24952 11008
rect 24544 10968 24952 10996
rect 24544 10956 24550 10968
rect 24946 10956 24952 10968
rect 25004 10996 25010 11008
rect 26142 10996 26148 11008
rect 25004 10968 26148 10996
rect 25004 10956 25010 10968
rect 26142 10956 26148 10968
rect 26200 10956 26206 11008
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 5626 10792 5632 10804
rect 5500 10764 5632 10792
rect 5500 10752 5506 10764
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5960 10764 6009 10792
rect 5960 10752 5966 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 9033 10795 9091 10801
rect 7800 10764 8984 10792
rect 7800 10752 7806 10764
rect 2590 10684 2596 10736
rect 2648 10684 2654 10736
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 7374 10724 7380 10736
rect 5123 10696 7380 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 8536 10696 8585 10724
rect 8536 10684 8542 10696
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 8956 10724 8984 10764
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9490 10792 9496 10804
rect 9079 10764 9496 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 11698 10792 11704 10804
rect 10376 10764 11704 10792
rect 10376 10752 10382 10764
rect 11698 10752 11704 10764
rect 11756 10792 11762 10804
rect 13906 10792 13912 10804
rect 11756 10764 13912 10792
rect 11756 10752 11762 10764
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 15470 10792 15476 10804
rect 14783 10764 15476 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 16172 10764 16313 10792
rect 16172 10752 16178 10764
rect 16301 10761 16313 10764
rect 16347 10792 16359 10795
rect 16390 10792 16396 10804
rect 16347 10764 16396 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 10045 10727 10103 10733
rect 10045 10724 10057 10727
rect 8956 10696 10057 10724
rect 8573 10687 8631 10693
rect 10045 10693 10057 10696
rect 10091 10693 10103 10727
rect 10045 10687 10103 10693
rect 13164 10727 13222 10733
rect 13164 10693 13176 10727
rect 13210 10724 13222 10727
rect 17770 10724 17776 10736
rect 13210 10696 17776 10724
rect 13210 10693 13222 10696
rect 13164 10687 13222 10693
rect 17770 10684 17776 10696
rect 17828 10724 17834 10736
rect 18248 10724 18276 10755
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19392 10764 19809 10792
rect 19392 10752 19398 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 21358 10792 21364 10804
rect 19797 10755 19855 10761
rect 20732 10764 21364 10792
rect 17828 10696 18276 10724
rect 17828 10684 17834 10696
rect 19150 10684 19156 10736
rect 19208 10724 19214 10736
rect 19429 10727 19487 10733
rect 19429 10724 19441 10727
rect 19208 10696 19441 10724
rect 19208 10684 19214 10696
rect 19429 10693 19441 10696
rect 19475 10693 19487 10727
rect 19429 10687 19487 10693
rect 19645 10727 19703 10733
rect 19645 10693 19657 10727
rect 19691 10724 19703 10727
rect 19978 10724 19984 10736
rect 19691 10696 19984 10724
rect 19691 10693 19703 10696
rect 19645 10687 19703 10693
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4304 10628 4813 10656
rect 4304 10616 4310 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5224 10628 5733 10656
rect 5224 10616 5230 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6236 10628 6561 10656
rect 6236 10616 6242 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6696 10628 6745 10656
rect 6696 10616 6702 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7098 10616 7104 10668
rect 7156 10616 7162 10668
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 7800 10628 8217 10656
rect 7800 10616 7806 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9582 10656 9588 10668
rect 9324 10628 9588 10656
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 3476 10560 6009 10588
rect 3476 10548 3482 10560
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 9324 10588 9352 10628
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9916 10628 10241 10656
rect 9916 10616 9922 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10376 10628 10425 10656
rect 10376 10616 10382 10628
rect 10413 10625 10425 10628
rect 10459 10656 10471 10659
rect 11606 10656 11612 10668
rect 10459 10628 11612 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12894 10616 12900 10668
rect 12952 10616 12958 10668
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 13964 10628 15301 10656
rect 13964 10616 13970 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15654 10656 15660 10668
rect 15519 10628 15660 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15654 10616 15660 10628
rect 15712 10656 15718 10668
rect 15838 10656 15844 10668
rect 15712 10628 15844 10656
rect 15712 10616 15718 10628
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 16022 10616 16028 10668
rect 16080 10656 16086 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 16080 10628 16129 10656
rect 16080 10616 16086 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 16850 10616 16856 10668
rect 16908 10616 16914 10668
rect 17120 10659 17178 10665
rect 17120 10625 17132 10659
rect 17166 10656 17178 10659
rect 17166 10628 17954 10656
rect 17166 10625 17178 10628
rect 17120 10619 17178 10625
rect 8527 10560 9352 10588
rect 9493 10591 9551 10597
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 7006 10480 7012 10532
rect 7064 10480 7070 10532
rect 9508 10520 9536 10551
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10505 10591 10563 10597
rect 10505 10588 10517 10591
rect 9732 10560 10517 10588
rect 9732 10548 9738 10560
rect 10505 10557 10517 10560
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14056 10560 15209 10588
rect 14056 10548 14062 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 8312 10492 9536 10520
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 3881 10455 3939 10461
rect 3881 10452 3893 10455
rect 1636 10424 3893 10452
rect 1636 10412 1642 10424
rect 3881 10421 3893 10424
rect 3927 10421 3939 10455
rect 3881 10415 3939 10421
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 5902 10452 5908 10464
rect 5859 10424 5908 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 8312 10452 8340 10492
rect 14090 10480 14096 10532
rect 14148 10520 14154 10532
rect 15105 10523 15163 10529
rect 15105 10520 15117 10523
rect 14148 10492 15117 10520
rect 14148 10480 14154 10492
rect 15105 10489 15117 10492
rect 15151 10489 15163 10523
rect 17926 10520 17954 10628
rect 18874 10616 18880 10668
rect 18932 10656 18938 10668
rect 18932 10628 20576 10656
rect 18932 10616 18938 10628
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19610 10588 19616 10600
rect 19208 10560 19616 10588
rect 19208 10548 19214 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 20548 10588 20576 10628
rect 20622 10616 20628 10668
rect 20680 10616 20686 10668
rect 20732 10656 20760 10764
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 23842 10792 23848 10804
rect 22112 10764 23848 10792
rect 20809 10727 20867 10733
rect 20809 10693 20821 10727
rect 20855 10724 20867 10727
rect 22002 10724 22008 10736
rect 20855 10696 22008 10724
rect 20855 10693 20867 10696
rect 20809 10687 20867 10693
rect 22002 10684 22008 10696
rect 22060 10684 22066 10736
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 20732 10628 20913 10656
rect 20901 10625 20913 10628
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 20993 10659 21051 10665
rect 20993 10625 21005 10659
rect 21039 10656 21051 10659
rect 21542 10656 21548 10668
rect 21039 10628 21548 10656
rect 21039 10625 21051 10628
rect 20993 10619 21051 10625
rect 21542 10616 21548 10628
rect 21600 10616 21606 10668
rect 22002 10588 22008 10600
rect 20548 10560 22008 10588
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 19518 10520 19524 10532
rect 17926 10492 19524 10520
rect 15105 10483 15163 10489
rect 19518 10480 19524 10492
rect 19576 10520 19582 10532
rect 21450 10520 21456 10532
rect 19576 10492 21456 10520
rect 19576 10480 19582 10492
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 7524 10424 8340 10452
rect 7524 10412 7530 10424
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9272 10424 9413 10452
rect 9272 10412 9278 10424
rect 9401 10421 9413 10424
rect 9447 10452 9459 10455
rect 10318 10452 10324 10464
rect 9447 10424 10324 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 14240 10424 14289 10452
rect 14240 10412 14246 10424
rect 14277 10421 14289 10424
rect 14323 10452 14335 10455
rect 14734 10452 14740 10464
rect 14323 10424 14740 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10452 15071 10455
rect 18506 10452 18512 10464
rect 15059 10424 18512 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 19610 10412 19616 10464
rect 19668 10412 19674 10464
rect 21174 10412 21180 10464
rect 21232 10412 21238 10464
rect 22112 10452 22140 10764
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 24118 10752 24124 10804
rect 24176 10792 24182 10804
rect 24673 10795 24731 10801
rect 24673 10792 24685 10795
rect 24176 10764 24685 10792
rect 24176 10752 24182 10764
rect 24673 10761 24685 10764
rect 24719 10761 24731 10795
rect 24673 10755 24731 10761
rect 24762 10752 24768 10804
rect 24820 10792 24826 10804
rect 25314 10792 25320 10804
rect 24820 10764 25320 10792
rect 24820 10752 24826 10764
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 25866 10752 25872 10804
rect 25924 10792 25930 10804
rect 26605 10795 26663 10801
rect 26605 10792 26617 10795
rect 25924 10764 26617 10792
rect 25924 10752 25930 10764
rect 26605 10761 26617 10764
rect 26651 10761 26663 10795
rect 26605 10755 26663 10761
rect 27522 10752 27528 10804
rect 27580 10792 27586 10804
rect 27709 10795 27767 10801
rect 27709 10792 27721 10795
rect 27580 10764 27721 10792
rect 27580 10752 27586 10764
rect 27709 10761 27721 10764
rect 27755 10761 27767 10795
rect 27709 10755 27767 10761
rect 22186 10684 22192 10736
rect 22244 10684 22250 10736
rect 22370 10684 22376 10736
rect 22428 10724 22434 10736
rect 24305 10727 24363 10733
rect 24305 10724 24317 10727
rect 22428 10696 24317 10724
rect 22428 10684 22434 10696
rect 24305 10693 24317 10696
rect 24351 10693 24363 10727
rect 24305 10687 24363 10693
rect 24394 10684 24400 10736
rect 24452 10724 24458 10736
rect 24505 10727 24563 10733
rect 24505 10724 24517 10727
rect 24452 10696 24517 10724
rect 24452 10684 24458 10696
rect 24505 10693 24517 10696
rect 24551 10693 24563 10727
rect 24505 10687 24563 10693
rect 22465 10659 22523 10665
rect 22465 10625 22477 10659
rect 22511 10656 22523 10659
rect 22830 10656 22836 10668
rect 22511 10628 22836 10656
rect 22511 10625 22523 10628
rect 22465 10619 22523 10625
rect 22830 10616 22836 10628
rect 22888 10616 22894 10668
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10656 23351 10659
rect 23382 10656 23388 10668
rect 23339 10628 23388 10656
rect 23339 10625 23351 10628
rect 23293 10619 23351 10625
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10625 23627 10659
rect 23569 10619 23627 10625
rect 22370 10548 22376 10600
rect 22428 10548 22434 10600
rect 23584 10588 23612 10619
rect 23658 10616 23664 10668
rect 23716 10616 23722 10668
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25130 10656 25136 10668
rect 24912 10628 25136 10656
rect 24912 10616 24918 10628
rect 25130 10616 25136 10628
rect 25188 10656 25194 10668
rect 25225 10659 25283 10665
rect 25225 10656 25237 10659
rect 25188 10628 25237 10656
rect 25188 10616 25194 10628
rect 25225 10625 25237 10628
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 25481 10659 25539 10665
rect 25481 10656 25493 10659
rect 25372 10628 25493 10656
rect 25372 10616 25378 10628
rect 25481 10625 25493 10628
rect 25527 10625 25539 10659
rect 25481 10619 25539 10625
rect 27154 10616 27160 10668
rect 27212 10616 27218 10668
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10625 27399 10659
rect 27341 10619 27399 10625
rect 24946 10588 24952 10600
rect 23584 10560 24952 10588
rect 24946 10548 24952 10560
rect 25004 10548 25010 10600
rect 26234 10548 26240 10600
rect 26292 10588 26298 10600
rect 27062 10588 27068 10600
rect 26292 10560 27068 10588
rect 26292 10548 26298 10560
rect 27062 10548 27068 10560
rect 27120 10588 27126 10600
rect 27356 10588 27384 10619
rect 27430 10616 27436 10668
rect 27488 10616 27494 10668
rect 27525 10659 27583 10665
rect 27525 10625 27537 10659
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27120 10560 27384 10588
rect 27120 10548 27126 10560
rect 22189 10455 22247 10461
rect 22189 10452 22201 10455
rect 22112 10424 22201 10452
rect 22189 10421 22201 10424
rect 22235 10421 22247 10455
rect 22189 10415 22247 10421
rect 22646 10412 22652 10464
rect 22704 10412 22710 10464
rect 23842 10412 23848 10464
rect 23900 10412 23906 10464
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 25038 10452 25044 10464
rect 24535 10424 25044 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25222 10412 25228 10464
rect 25280 10452 25286 10464
rect 27540 10452 27568 10619
rect 25280 10424 27568 10452
rect 25280 10412 25286 10424
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1762 10208 1768 10260
rect 1820 10208 1826 10260
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3510 10248 3516 10260
rect 2731 10220 3516 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4154 10248 4160 10260
rect 4019 10220 4160 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4856 10220 5273 10248
rect 4856 10208 4862 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 7190 10248 7196 10260
rect 6696 10220 7196 10248
rect 6696 10208 6702 10220
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 9214 10208 9220 10260
rect 9272 10208 9278 10260
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 10594 10208 10600 10260
rect 10652 10208 10658 10260
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 10704 10220 16129 10248
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 4062 10180 4068 10192
rect 3375 10152 4068 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 4341 10183 4399 10189
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 4706 10180 4712 10192
rect 4387 10152 4712 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 4706 10140 4712 10152
rect 4764 10180 4770 10192
rect 7282 10180 7288 10192
rect 4764 10152 7288 10180
rect 4764 10140 4770 10152
rect 7282 10140 7288 10152
rect 7340 10140 7346 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 10704 10180 10732 10220
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 16117 10211 16175 10217
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 17957 10251 18015 10257
rect 17957 10248 17969 10251
rect 17368 10220 17969 10248
rect 17368 10208 17374 10220
rect 17957 10217 17969 10220
rect 18003 10217 18015 10251
rect 17957 10211 18015 10217
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18196 10220 18429 10248
rect 18196 10208 18202 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18417 10211 18475 10217
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 20530 10248 20536 10260
rect 18840 10220 20536 10248
rect 18840 10208 18846 10220
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 20990 10248 20996 10260
rect 20763 10220 20996 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 21821 10251 21879 10257
rect 21821 10248 21833 10251
rect 21324 10220 21833 10248
rect 21324 10208 21330 10220
rect 21821 10217 21833 10220
rect 21867 10217 21879 10251
rect 21821 10211 21879 10217
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 23198 10248 23204 10260
rect 22060 10220 23204 10248
rect 22060 10208 22066 10220
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 23382 10208 23388 10260
rect 23440 10248 23446 10260
rect 25774 10248 25780 10260
rect 23440 10220 25780 10248
rect 23440 10208 23446 10220
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 26786 10208 26792 10260
rect 26844 10248 26850 10260
rect 28353 10251 28411 10257
rect 28353 10248 28365 10251
rect 26844 10220 28365 10248
rect 26844 10208 26850 10220
rect 28353 10217 28365 10220
rect 28399 10217 28411 10251
rect 28353 10211 28411 10217
rect 8444 10152 10732 10180
rect 12805 10183 12863 10189
rect 8444 10140 8450 10152
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 13722 10180 13728 10192
rect 12851 10152 13728 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 19334 10180 19340 10192
rect 16316 10152 19340 10180
rect 5166 10112 5172 10124
rect 2792 10084 4476 10112
rect 842 10004 848 10056
rect 900 10044 906 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 900 10016 1593 10044
rect 900 10004 906 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 2590 10004 2596 10056
rect 2648 10004 2654 10056
rect 2792 10053 2820 10084
rect 4448 10056 4476 10084
rect 4816 10084 5172 10112
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3252 9976 3280 10007
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4338 10044 4344 10056
rect 4203 10016 4344 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4816 9976 4844 10084
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 7374 10112 7380 10124
rect 5224 10084 5488 10112
rect 5224 10072 5230 10084
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5460 10053 5488 10084
rect 6380 10084 7380 10112
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 4948 10016 5273 10044
rect 4948 10004 4954 10016
rect 5261 10013 5273 10016
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6380 10053 6408 10084
rect 7374 10072 7380 10084
rect 7432 10112 7438 10124
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 7432 10084 7665 10112
rect 7432 10072 7438 10084
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 6236 10016 6377 10044
rect 6236 10004 6242 10016
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6638 10044 6644 10056
rect 6595 10016 6644 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7156 10016 7205 10044
rect 7156 10004 7162 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7282 10004 7288 10056
rect 7340 10044 7346 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7340 10016 7481 10044
rect 7340 10004 7346 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7616 10016 8309 10044
rect 7616 10004 7622 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 9122 10004 9128 10056
rect 9180 10004 9186 10056
rect 9416 10044 9444 10075
rect 10134 10072 10140 10124
rect 10192 10072 10198 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10318 10112 10324 10124
rect 10275 10084 10324 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11204 10084 11437 10112
rect 11204 10072 11210 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 9858 10053 9864 10056
rect 9849 10047 9864 10053
rect 9849 10044 9861 10047
rect 9416 10016 9861 10044
rect 9849 10013 9861 10016
rect 9849 10007 9864 10013
rect 9858 10004 9864 10007
rect 9916 10004 9922 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 3252 9948 4844 9976
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6454 9976 6460 9988
rect 5960 9948 6460 9976
rect 5960 9936 5966 9948
rect 6454 9936 6460 9948
rect 6512 9976 6518 9988
rect 8389 9979 8447 9985
rect 8389 9976 8401 9979
rect 6512 9948 8401 9976
rect 6512 9936 6518 9948
rect 8389 9945 8401 9948
rect 8435 9945 8447 9979
rect 10060 9976 10088 10007
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 13722 10044 13728 10056
rect 11532 10016 13728 10044
rect 11532 9976 11560 10016
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 11681 9979 11739 9985
rect 11681 9976 11693 9979
rect 10060 9948 11560 9976
rect 11624 9948 11693 9976
rect 8389 9939 8447 9945
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 7282 9868 7288 9920
rect 7340 9868 7346 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 11624 9908 11652 9948
rect 11681 9945 11693 9948
rect 11727 9945 11739 9979
rect 11681 9939 11739 9945
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 12894 9976 12900 9988
rect 11848 9948 12900 9976
rect 11848 9936 11854 9948
rect 12894 9936 12900 9948
rect 12952 9976 12958 9988
rect 14292 9976 14320 10072
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16316 10053 16344 10152
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 19444 10152 19565 10180
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 19444 10112 19472 10152
rect 18187 10084 19472 10112
rect 19537 10112 19565 10152
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 19668 10152 22293 10180
rect 19668 10140 19674 10152
rect 22281 10149 22293 10152
rect 22327 10149 22339 10183
rect 22281 10143 22339 10149
rect 23566 10140 23572 10192
rect 23624 10180 23630 10192
rect 23661 10183 23719 10189
rect 23661 10180 23673 10183
rect 23624 10152 23673 10180
rect 23624 10140 23630 10152
rect 23661 10149 23673 10152
rect 23707 10149 23719 10183
rect 23661 10143 23719 10149
rect 24026 10140 24032 10192
rect 24084 10180 24090 10192
rect 24670 10180 24676 10192
rect 24084 10152 24676 10180
rect 24084 10140 24090 10152
rect 24670 10140 24676 10152
rect 24728 10140 24734 10192
rect 19537 10084 21281 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 19392 10016 19441 10044
rect 19392 10004 19398 10016
rect 19429 10013 19441 10016
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 19576 10016 19621 10044
rect 19576 10004 19582 10016
rect 19886 10004 19892 10056
rect 19944 10053 19950 10056
rect 19944 10044 19952 10053
rect 20346 10044 20352 10056
rect 19944 10016 20352 10044
rect 19944 10007 19952 10016
rect 19944 10004 19950 10007
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 21082 10044 21088 10056
rect 20456 10016 21088 10044
rect 12952 9948 14320 9976
rect 12952 9936 12958 9948
rect 14474 9936 14480 9988
rect 14532 9985 14538 9988
rect 14532 9979 14580 9985
rect 14532 9945 14534 9979
rect 14568 9945 14580 9979
rect 14532 9939 14580 9945
rect 14532 9936 14538 9939
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 16758 9976 16764 9988
rect 14884 9948 16764 9976
rect 14884 9936 14890 9948
rect 16758 9936 16764 9948
rect 16816 9936 16822 9988
rect 17770 9936 17776 9988
rect 17828 9936 17834 9988
rect 18046 9936 18052 9988
rect 18104 9976 18110 9988
rect 19705 9979 19763 9985
rect 18104 9948 19288 9976
rect 18104 9936 18110 9948
rect 9732 9880 11652 9908
rect 15657 9911 15715 9917
rect 9732 9868 9738 9880
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 19150 9908 19156 9920
rect 15703 9880 19156 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19260 9908 19288 9948
rect 19705 9945 19717 9979
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 20456 9976 20484 10016
rect 21082 10004 21088 10016
rect 21140 10004 21146 10056
rect 19843 9948 20484 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 19720 9908 19748 9939
rect 20530 9936 20536 9988
rect 20588 9936 20594 9988
rect 20806 9985 20812 9988
rect 20749 9979 20812 9985
rect 20749 9945 20761 9979
rect 20795 9945 20812 9979
rect 20749 9939 20812 9945
rect 20806 9936 20812 9939
rect 20864 9936 20870 9988
rect 19260 9880 19748 9908
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 19944 9880 20085 9908
rect 19944 9868 19950 9880
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 20898 9868 20904 9920
rect 20956 9868 20962 9920
rect 21253 9908 21281 10084
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 21913 10115 21971 10121
rect 21913 10112 21925 10115
rect 21692 10084 21925 10112
rect 21692 10072 21698 10084
rect 21913 10081 21925 10084
rect 21959 10081 21971 10115
rect 21913 10075 21971 10081
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 22097 10047 22155 10053
rect 22097 10013 22109 10047
rect 22143 10044 22155 10047
rect 22278 10044 22284 10056
rect 22143 10016 22284 10044
rect 22143 10013 22155 10016
rect 22097 10007 22155 10013
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 23106 10004 23112 10056
rect 23164 10004 23170 10056
rect 23198 10004 23204 10056
rect 23256 10044 23262 10056
rect 23293 10047 23351 10053
rect 23293 10044 23305 10047
rect 23256 10016 23305 10044
rect 23256 10004 23262 10016
rect 23293 10013 23305 10016
rect 23339 10013 23351 10047
rect 23293 10007 23351 10013
rect 23474 10004 23480 10056
rect 23532 10044 23538 10056
rect 24762 10044 24768 10056
rect 23532 10016 24768 10044
rect 23532 10004 23538 10016
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 25400 10047 25458 10053
rect 25400 10013 25412 10047
rect 25446 10044 25458 10047
rect 26878 10044 26884 10056
rect 25446 10016 26884 10044
rect 25446 10013 25458 10016
rect 25400 10007 25458 10013
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 21821 9979 21879 9985
rect 21821 9945 21833 9979
rect 21867 9976 21879 9979
rect 22462 9976 22468 9988
rect 21867 9948 22468 9976
rect 21867 9945 21879 9948
rect 21821 9939 21879 9945
rect 22462 9936 22468 9948
rect 22520 9936 22526 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9945 23443 9979
rect 23385 9939 23443 9945
rect 23198 9908 23204 9920
rect 21253 9880 23204 9908
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23400 9908 23428 9939
rect 25866 9936 25872 9988
rect 25924 9976 25930 9988
rect 27218 9979 27276 9985
rect 27218 9976 27230 9979
rect 25924 9948 27230 9976
rect 25924 9936 25930 9948
rect 27218 9945 27230 9948
rect 27264 9945 27276 9979
rect 27218 9939 27276 9945
rect 26513 9911 26571 9917
rect 26513 9908 26525 9911
rect 23400 9880 26525 9908
rect 26513 9877 26525 9880
rect 26559 9908 26571 9911
rect 26878 9908 26884 9920
rect 26559 9880 26884 9908
rect 26559 9877 26571 9880
rect 26513 9871 26571 9877
rect 26878 9868 26884 9880
rect 26936 9868 26942 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 4706 9704 4712 9716
rect 2648 9676 4712 9704
rect 2648 9664 2654 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4816 9676 5212 9704
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 4816 9636 4844 9676
rect 3283 9608 4844 9636
rect 4893 9639 4951 9645
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 4893 9605 4905 9639
rect 4939 9636 4951 9639
rect 5074 9636 5080 9648
rect 4939 9608 5080 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5184 9636 5212 9676
rect 7374 9664 7380 9716
rect 7432 9713 7438 9716
rect 7432 9707 7451 9713
rect 7439 9673 7451 9707
rect 7432 9667 7451 9673
rect 7432 9664 7438 9667
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 10410 9704 10416 9716
rect 7616 9676 10416 9704
rect 7616 9664 7622 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 13906 9704 13912 9716
rect 10744 9676 13912 9704
rect 10744 9664 10750 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 15194 9664 15200 9716
rect 15252 9664 15258 9716
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 19518 9704 19524 9716
rect 17828 9676 19524 9704
rect 17828 9664 17834 9676
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 20254 9704 20260 9716
rect 20040 9676 20260 9704
rect 5184 9608 7052 9636
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 5166 9568 5172 9580
rect 4295 9540 5172 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 1854 9460 1860 9512
rect 1912 9460 1918 9512
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4488 9472 4629 9500
rect 4488 9460 4494 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 4632 9432 4660 9463
rect 4706 9460 4712 9512
rect 4764 9460 4770 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5552 9500 5580 9531
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5757 9571 5815 9577
rect 5757 9537 5769 9571
rect 5803 9568 5815 9571
rect 5902 9568 5908 9580
rect 5803 9540 5908 9568
rect 5803 9537 5815 9540
rect 5757 9531 5815 9537
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 7024 9568 7052 9608
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 7156 9608 7205 9636
rect 7156 9596 7162 9608
rect 7193 9605 7205 9608
rect 7239 9605 7251 9639
rect 9214 9636 9220 9648
rect 7193 9599 7251 9605
rect 7300 9608 9220 9636
rect 7300 9568 7328 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 9576 9639 9634 9645
rect 9576 9605 9588 9639
rect 9622 9636 9634 9639
rect 12253 9639 12311 9645
rect 9622 9608 12020 9636
rect 9622 9605 9634 9608
rect 9576 9599 9634 9605
rect 7024 9540 7328 9568
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8478 9568 8484 9580
rect 8343 9540 8484 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 11146 9568 11152 9580
rect 9364 9540 11152 9568
rect 9364 9528 9370 9540
rect 11146 9528 11152 9540
rect 11204 9568 11210 9580
rect 11790 9568 11796 9580
rect 11204 9540 11796 9568
rect 11204 9528 11210 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 5132 9472 5580 9500
rect 5132 9460 5138 9472
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6696 9472 7604 9500
rect 6696 9460 6702 9472
rect 5353 9435 5411 9441
rect 4632 9404 4752 9432
rect 4724 9364 4752 9404
rect 5353 9401 5365 9435
rect 5399 9432 5411 9435
rect 5994 9432 6000 9444
rect 5399 9404 6000 9432
rect 5399 9401 5411 9404
rect 5353 9395 5411 9401
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 7576 9441 7604 9472
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 8444 9472 8585 9500
rect 8444 9460 8450 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 11992 9500 12020 9608
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12526 9636 12532 9648
rect 12299 9608 12532 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 13072 9639 13130 9645
rect 13072 9605 13084 9639
rect 13118 9636 13130 9639
rect 13814 9636 13820 9648
rect 13118 9608 13820 9636
rect 13118 9605 13130 9608
rect 13072 9599 13130 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 16022 9636 16028 9648
rect 15212 9608 16028 9636
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12805 9571 12863 9577
rect 12115 9540 12434 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12250 9500 12256 9512
rect 11992 9472 12256 9500
rect 8573 9463 8631 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 7561 9435 7619 9441
rect 6512 9404 7512 9432
rect 6512 9392 6518 9404
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 4724 9336 6653 9364
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 7248 9336 7389 9364
rect 7248 9324 7254 9336
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 7484 9364 7512 9404
rect 7561 9401 7573 9435
rect 7607 9401 7619 9435
rect 7561 9395 7619 9401
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 7800 9404 8493 9432
rect 7800 9392 7806 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 7484 9336 8125 9364
rect 7377 9327 7435 9333
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8113 9327 8171 9333
rect 10686 9324 10692 9376
rect 10744 9324 10750 9376
rect 12406 9364 12434 9540
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 12894 9568 12900 9580
rect 12851 9540 12900 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 15212 9577 15240 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 17586 9596 17592 9648
rect 17644 9636 17650 9648
rect 18046 9636 18052 9648
rect 17644 9608 18052 9636
rect 17644 9596 17650 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 18196 9608 19840 9636
rect 18196 9596 18202 9608
rect 15197 9571 15255 9577
rect 13412 9540 13860 9568
rect 13412 9528 13418 9540
rect 13832 9500 13860 9540
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9568 15439 9571
rect 15470 9568 15476 9580
rect 15427 9540 15476 9568
rect 15427 9537 15439 9540
rect 15381 9531 15439 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 16666 9568 16672 9580
rect 15887 9540 16672 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 15580 9500 15608 9531
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 19812 9577 19840 9608
rect 19886 9596 19892 9648
rect 19944 9596 19950 9648
rect 20040 9577 20068 9676
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 22465 9707 22523 9713
rect 22465 9704 22477 9707
rect 21416 9676 22477 9704
rect 21416 9664 21422 9676
rect 22465 9673 22477 9676
rect 22511 9673 22523 9707
rect 23658 9704 23664 9716
rect 22465 9667 22523 9673
rect 22572 9676 23664 9704
rect 20099 9639 20157 9645
rect 20099 9605 20111 9639
rect 20145 9636 20157 9639
rect 22572 9636 22600 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 25056 9676 25360 9704
rect 23842 9636 23848 9648
rect 20145 9608 22600 9636
rect 22664 9608 23848 9636
rect 20145 9605 20162 9608
rect 20099 9599 20162 9605
rect 19797 9571 19855 9577
rect 17736 9540 19748 9568
rect 17736 9528 17742 9540
rect 13832 9472 15608 9500
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 18506 9500 18512 9512
rect 17276 9472 18512 9500
rect 17276 9460 17282 9472
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 14274 9432 14280 9444
rect 13740 9404 14280 9432
rect 13740 9364 13768 9404
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 16298 9432 16304 9444
rect 15528 9404 16304 9432
rect 15528 9392 15534 9404
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18690 9432 18696 9444
rect 18012 9404 18696 9432
rect 18012 9392 18018 9404
rect 18690 9392 18696 9404
rect 18748 9432 18754 9444
rect 19518 9432 19524 9444
rect 18748 9404 19524 9432
rect 18748 9392 18754 9404
rect 19518 9392 19524 9404
rect 19576 9392 19582 9444
rect 19720 9432 19748 9540
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 20006 9571 20068 9577
rect 20006 9537 20018 9571
rect 20052 9540 20068 9571
rect 20052 9537 20064 9540
rect 20006 9531 20064 9537
rect 19812 9500 19840 9531
rect 19886 9500 19892 9512
rect 19812 9472 19892 9500
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 20134 9500 20162 9599
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9568 20315 9571
rect 20901 9571 20959 9577
rect 20303 9540 20852 9568
rect 20303 9537 20315 9540
rect 20257 9531 20315 9537
rect 19996 9472 20162 9500
rect 19996 9432 20024 9472
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20717 9503 20775 9509
rect 20717 9500 20729 9503
rect 20496 9472 20729 9500
rect 20496 9460 20502 9472
rect 20717 9469 20729 9472
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 20824 9444 20852 9540
rect 20901 9537 20913 9571
rect 20947 9568 20959 9571
rect 20990 9568 20996 9580
rect 20947 9540 20996 9568
rect 20947 9537 20959 9540
rect 20901 9531 20959 9537
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9568 22431 9571
rect 22462 9568 22468 9580
rect 22419 9540 22468 9568
rect 22419 9537 22431 9540
rect 22373 9531 22431 9537
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9500 22615 9503
rect 22664 9500 22692 9608
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 24118 9596 24124 9648
rect 24176 9636 24182 9648
rect 25056 9636 25084 9676
rect 24176 9608 25084 9636
rect 25332 9636 25360 9676
rect 25498 9664 25504 9716
rect 25556 9704 25562 9716
rect 25777 9707 25835 9713
rect 25777 9704 25789 9707
rect 25556 9676 25789 9704
rect 25556 9664 25562 9676
rect 25777 9673 25789 9676
rect 25823 9673 25835 9707
rect 25777 9667 25835 9673
rect 25332 9608 25452 9636
rect 24176 9596 24182 9608
rect 22738 9528 22744 9580
rect 22796 9528 22802 9580
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 23382 9568 23388 9580
rect 23339 9540 23388 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 25424 9577 25452 9608
rect 23560 9571 23618 9577
rect 23560 9537 23572 9571
rect 23606 9568 23618 9571
rect 25133 9571 25191 9577
rect 23606 9540 25084 9568
rect 23606 9537 23618 9540
rect 23560 9531 23618 9537
rect 22603 9472 22692 9500
rect 22603 9469 22615 9472
rect 22557 9463 22615 9469
rect 19720 9404 20024 9432
rect 20806 9392 20812 9444
rect 20864 9392 20870 9444
rect 22649 9435 22707 9441
rect 22649 9401 22661 9435
rect 22695 9432 22707 9435
rect 23014 9432 23020 9444
rect 22695 9404 23020 9432
rect 22695 9401 22707 9404
rect 22649 9395 22707 9401
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 12406 9336 13768 9364
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 14366 9364 14372 9376
rect 14231 9336 14372 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16666 9364 16672 9376
rect 15344 9336 16672 9364
rect 15344 9324 15350 9336
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 19150 9324 19156 9376
rect 19208 9364 19214 9376
rect 19613 9367 19671 9373
rect 19613 9364 19625 9367
rect 19208 9336 19625 9364
rect 19208 9324 19214 9336
rect 19613 9333 19625 9336
rect 19659 9333 19671 9367
rect 19613 9327 19671 9333
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 21085 9367 21143 9373
rect 21085 9364 21097 9367
rect 20588 9336 21097 9364
rect 20588 9324 20594 9336
rect 21085 9333 21097 9336
rect 21131 9364 21143 9367
rect 22554 9364 22560 9376
rect 21131 9336 22560 9364
rect 21131 9333 21143 9336
rect 21085 9327 21143 9333
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 24673 9367 24731 9373
rect 24673 9364 24685 9367
rect 23164 9336 24685 9364
rect 23164 9324 23170 9336
rect 24673 9333 24685 9336
rect 24719 9333 24731 9367
rect 25056 9364 25084 9540
rect 25133 9537 25145 9571
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 25226 9571 25284 9577
rect 25226 9537 25238 9571
rect 25272 9537 25284 9571
rect 25226 9531 25284 9537
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25148 9432 25176 9531
rect 25240 9500 25268 9531
rect 25498 9528 25504 9580
rect 25556 9528 25562 9580
rect 25639 9571 25697 9577
rect 25639 9537 25651 9571
rect 25685 9568 25697 9571
rect 26326 9568 26332 9580
rect 25685 9540 26332 9568
rect 25685 9537 25697 9540
rect 25639 9531 25697 9537
rect 26068 9512 26096 9540
rect 26326 9528 26332 9540
rect 26384 9528 26390 9580
rect 25958 9500 25964 9512
rect 25240 9472 25964 9500
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 26050 9460 26056 9512
rect 26108 9460 26114 9512
rect 25406 9432 25412 9444
rect 25148 9404 25412 9432
rect 25406 9392 25412 9404
rect 25464 9392 25470 9444
rect 25498 9392 25504 9444
rect 25556 9432 25562 9444
rect 27890 9432 27896 9444
rect 25556 9404 27896 9432
rect 25556 9392 25562 9404
rect 27890 9392 27896 9404
rect 27948 9392 27954 9444
rect 26510 9364 26516 9376
rect 25056 9336 26516 9364
rect 24673 9327 24731 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 2961 9163 3019 9169
rect 1912 9132 2774 9160
rect 1912 9120 1918 9132
rect 2746 9092 2774 9132
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3326 9160 3332 9172
rect 3007 9132 3332 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4798 9160 4804 9172
rect 4203 9132 4804 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 5868 9132 6377 9160
rect 5868 9120 5874 9132
rect 6365 9129 6377 9132
rect 6411 9129 6423 9163
rect 6365 9123 6423 9129
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 6880 9132 7573 9160
rect 6880 9120 6886 9132
rect 7561 9129 7573 9132
rect 7607 9129 7619 9163
rect 7561 9123 7619 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9585 9163 9643 9169
rect 9585 9160 9597 9163
rect 9364 9132 9597 9160
rect 9364 9120 9370 9132
rect 9585 9129 9597 9132
rect 9631 9129 9643 9163
rect 9585 9123 9643 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 15194 9160 15200 9172
rect 9824 9132 15200 9160
rect 9824 9120 9830 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 16025 9163 16083 9169
rect 16025 9129 16037 9163
rect 16071 9160 16083 9163
rect 16850 9160 16856 9172
rect 16071 9132 16856 9160
rect 16071 9129 16083 9132
rect 16025 9123 16083 9129
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 16942 9120 16948 9172
rect 17000 9160 17006 9172
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17000 9132 17325 9160
rect 17000 9120 17006 9132
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 17313 9123 17371 9129
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 19242 9160 19248 9172
rect 18564 9132 19248 9160
rect 18564 9120 18570 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 19518 9120 19524 9172
rect 19576 9120 19582 9172
rect 23290 9160 23296 9172
rect 19720 9132 23296 9160
rect 7006 9092 7012 9104
rect 2746 9064 6316 9092
rect 1578 8984 1584 9036
rect 1636 8984 1642 9036
rect 5258 9024 5264 9036
rect 4356 8996 5264 9024
rect 4356 8965 4384 8996
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 4798 8956 4804 8968
rect 4663 8928 4804 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5718 8956 5724 8968
rect 5123 8928 5724 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 1848 8891 1906 8897
rect 1848 8857 1860 8891
rect 1894 8888 1906 8891
rect 1946 8888 1952 8900
rect 1894 8860 1952 8888
rect 1894 8857 1906 8860
rect 1848 8851 1906 8857
rect 1946 8848 1952 8860
rect 2004 8848 2010 8900
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 5224 8860 5273 8888
rect 5224 8848 5230 8860
rect 5261 8857 5273 8860
rect 5307 8857 5319 8891
rect 5261 8851 5319 8857
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 4890 8820 4896 8832
rect 4571 8792 4896 8820
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 5408 8792 5457 8820
rect 5408 8780 5414 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 6288 8820 6316 9064
rect 6564 9064 7012 9092
rect 6564 8965 6592 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 13446 9092 13452 9104
rect 11756 9064 13452 9092
rect 11756 9052 11762 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 13633 9095 13691 9101
rect 13633 9092 13645 9095
rect 13596 9064 13645 9092
rect 13596 9052 13602 9064
rect 13633 9061 13645 9064
rect 13679 9061 13691 9095
rect 13633 9055 13691 9061
rect 14642 9052 14648 9104
rect 14700 9092 14706 9104
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 14700 9064 14933 9092
rect 14700 9052 14706 9064
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 15160 9064 15884 9092
rect 15160 9052 15166 9064
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6696 8996 7052 9024
rect 6696 8984 6702 8996
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7024 8965 7052 8996
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7248 8996 7788 9024
rect 7248 8984 7254 8996
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6641 8891 6699 8897
rect 6641 8888 6653 8891
rect 6420 8860 6653 8888
rect 6420 8848 6426 8860
rect 6641 8857 6653 8860
rect 6687 8857 6699 8891
rect 6932 8888 6960 8919
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7760 8965 7788 8996
rect 11790 8984 11796 9036
rect 11848 8984 11854 9036
rect 12544 8996 13492 9024
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7432 8928 7573 8956
rect 7432 8916 7438 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8996 8928 9413 8956
rect 8996 8916 9002 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 11882 8956 11888 8968
rect 11563 8928 11888 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 11882 8916 11888 8928
rect 11940 8956 11946 8968
rect 12544 8956 12572 8996
rect 11940 8928 12572 8956
rect 11940 8916 11946 8928
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 13464 8965 13492 8996
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 14792 8996 15025 9024
rect 14792 8984 14798 8996
rect 15013 8993 15025 8996
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13998 8956 14004 8968
rect 13495 8928 14004 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14608 8928 14841 8956
rect 14608 8916 14614 8928
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 7282 8888 7288 8900
rect 6932 8860 7288 8888
rect 6641 8851 6699 8857
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 12158 8888 12164 8900
rect 10836 8860 12164 8888
rect 10836 8848 10842 8860
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12345 8891 12403 8897
rect 12345 8857 12357 8891
rect 12391 8888 12403 8891
rect 12391 8860 13492 8888
rect 12391 8857 12403 8860
rect 12345 8851 12403 8857
rect 13464 8832 13492 8860
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 14642 8888 14648 8900
rect 14516 8860 14648 8888
rect 14516 8848 14522 8860
rect 14642 8848 14648 8860
rect 14700 8888 14706 8900
rect 15120 8888 15148 8919
rect 15286 8916 15292 8968
rect 15344 8916 15350 8968
rect 14700 8860 15148 8888
rect 15749 8891 15807 8897
rect 14700 8848 14706 8860
rect 15749 8857 15761 8891
rect 15795 8857 15807 8891
rect 15856 8888 15884 9064
rect 16206 9052 16212 9104
rect 16264 9052 16270 9104
rect 16298 9052 16304 9104
rect 16356 9092 16362 9104
rect 18877 9095 18935 9101
rect 18877 9092 18889 9095
rect 16356 9064 18889 9092
rect 16356 9052 16362 9064
rect 18877 9061 18889 9064
rect 18923 9061 18935 9095
rect 19720 9092 19748 9132
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 24026 9120 24032 9172
rect 24084 9120 24090 9172
rect 25774 9120 25780 9172
rect 25832 9160 25838 9172
rect 26421 9163 26479 9169
rect 26421 9160 26433 9163
rect 25832 9132 26433 9160
rect 25832 9120 25838 9132
rect 26421 9129 26433 9132
rect 26467 9129 26479 9163
rect 26421 9123 26479 9129
rect 27246 9120 27252 9172
rect 27304 9160 27310 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 27304 9132 28273 9160
rect 27304 9120 27310 9132
rect 28261 9129 28273 9132
rect 28307 9129 28319 9163
rect 28261 9123 28319 9129
rect 18877 9055 18935 9061
rect 19536 9064 19748 9092
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 19334 9024 19340 9036
rect 15979 8996 19340 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19536 9033 19564 9064
rect 19886 9052 19892 9104
rect 19944 9092 19950 9104
rect 20714 9092 20720 9104
rect 19944 9064 20720 9092
rect 19944 9052 19950 9064
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 8993 19579 9027
rect 20438 9024 20444 9036
rect 19521 8987 19579 8993
rect 19628 8996 20444 9024
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16482 8956 16488 8968
rect 16071 8928 16488 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8956 17187 8959
rect 17218 8956 17224 8968
rect 17175 8928 17224 8956
rect 17175 8925 17187 8928
rect 17129 8919 17187 8925
rect 16776 8888 16804 8919
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 15856 8860 16804 8888
rect 16945 8891 17003 8897
rect 15749 8851 15807 8857
rect 16945 8857 16957 8891
rect 16991 8857 17003 8891
rect 16945 8851 17003 8857
rect 17037 8891 17095 8897
rect 17037 8857 17049 8891
rect 17083 8888 17095 8891
rect 17586 8888 17592 8900
rect 17083 8860 17592 8888
rect 17083 8857 17095 8860
rect 17037 8851 17095 8857
rect 9858 8820 9864 8832
rect 6288 8792 9864 8820
rect 5445 8783 5503 8789
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12032 8792 12541 8820
rect 12032 8780 12038 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 12529 8783 12587 8789
rect 12894 8780 12900 8832
rect 12952 8780 12958 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 14553 8823 14611 8829
rect 14553 8789 14565 8823
rect 14599 8820 14611 8823
rect 15378 8820 15384 8832
rect 14599 8792 15384 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15764 8820 15792 8851
rect 16482 8820 16488 8832
rect 15764 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16960 8820 16988 8851
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 17494 8820 17500 8832
rect 16960 8792 17500 8820
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 18248 8820 18276 8919
rect 18322 8916 18328 8968
rect 18380 8916 18386 8968
rect 18414 8916 18420 8968
rect 18472 8916 18478 8968
rect 18506 8916 18512 8968
rect 18564 8916 18570 8968
rect 18598 8916 18604 8968
rect 18656 8916 18662 8968
rect 18698 8959 18756 8965
rect 18698 8925 18710 8959
rect 18744 8956 18756 8959
rect 18874 8956 18880 8968
rect 18744 8928 18880 8956
rect 18744 8925 18756 8928
rect 18698 8919 18756 8925
rect 18432 8888 18460 8916
rect 18708 8888 18736 8919
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19628 8956 19656 8996
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 19300 8928 19656 8956
rect 19300 8916 19306 8928
rect 19702 8916 19708 8968
rect 19760 8916 19766 8968
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 20128 8928 20821 8956
rect 20128 8916 20134 8928
rect 20809 8925 20821 8928
rect 20855 8956 20867 8959
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 20855 8928 22661 8956
rect 20855 8925 20867 8928
rect 20809 8919 20867 8925
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 25041 8959 25099 8965
rect 25041 8956 25053 8959
rect 23440 8928 25053 8956
rect 23440 8916 23446 8928
rect 25041 8925 25053 8928
rect 25087 8956 25099 8959
rect 25130 8956 25136 8968
rect 25087 8928 25136 8956
rect 25087 8925 25099 8928
rect 25041 8919 25099 8925
rect 25130 8916 25136 8928
rect 25188 8956 25194 8968
rect 26694 8956 26700 8968
rect 25188 8928 26700 8956
rect 25188 8916 25194 8928
rect 26694 8916 26700 8928
rect 26752 8956 26758 8968
rect 26881 8959 26939 8965
rect 26881 8956 26893 8959
rect 26752 8928 26893 8956
rect 26752 8916 26758 8928
rect 26881 8925 26893 8928
rect 26927 8956 26939 8959
rect 26970 8956 26976 8968
rect 26927 8928 26976 8956
rect 26927 8925 26939 8928
rect 26881 8919 26939 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 18432 8860 18736 8888
rect 19426 8848 19432 8900
rect 19484 8848 19490 8900
rect 20622 8888 20628 8900
rect 19813 8860 20628 8888
rect 19813 8820 19841 8860
rect 20622 8848 20628 8860
rect 20680 8848 20686 8900
rect 21082 8897 21088 8900
rect 21076 8888 21088 8897
rect 21043 8860 21088 8888
rect 21076 8851 21088 8860
rect 21082 8848 21088 8851
rect 21140 8848 21146 8900
rect 22916 8891 22974 8897
rect 22066 8860 22324 8888
rect 18248 8792 19841 8820
rect 19886 8780 19892 8832
rect 19944 8780 19950 8832
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20254 8820 20260 8832
rect 20128 8792 20260 8820
rect 20128 8780 20134 8792
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20990 8780 20996 8832
rect 21048 8820 21054 8832
rect 22066 8820 22094 8860
rect 21048 8792 22094 8820
rect 21048 8780 21054 8792
rect 22186 8780 22192 8832
rect 22244 8780 22250 8832
rect 22296 8820 22324 8860
rect 22916 8857 22928 8891
rect 22962 8888 22974 8891
rect 23106 8888 23112 8900
rect 22962 8860 23112 8888
rect 22962 8857 22974 8860
rect 22916 8851 22974 8857
rect 23106 8848 23112 8860
rect 23164 8848 23170 8900
rect 24394 8888 24400 8900
rect 23216 8860 24400 8888
rect 22830 8820 22836 8832
rect 22296 8792 22836 8820
rect 22830 8780 22836 8792
rect 22888 8820 22894 8832
rect 23216 8820 23244 8860
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 25314 8897 25320 8900
rect 25308 8888 25320 8897
rect 25275 8860 25320 8888
rect 25308 8851 25320 8860
rect 25314 8848 25320 8851
rect 25372 8848 25378 8900
rect 26602 8848 26608 8900
rect 26660 8888 26666 8900
rect 27154 8897 27160 8900
rect 27126 8891 27160 8897
rect 27126 8888 27138 8891
rect 26660 8860 27138 8888
rect 26660 8848 26666 8860
rect 27126 8857 27138 8860
rect 27126 8851 27160 8857
rect 27154 8848 27160 8851
rect 27212 8848 27218 8900
rect 22888 8792 23244 8820
rect 22888 8780 22894 8792
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 6822 8576 6828 8628
rect 6880 8576 6886 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7282 8616 7288 8628
rect 7064 8588 7288 8616
rect 7064 8576 7070 8588
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7800 8588 7941 8616
rect 7800 8576 7806 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12492 8588 13093 8616
rect 12492 8576 12498 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 15841 8619 15899 8625
rect 13780 8588 15516 8616
rect 13780 8576 13786 8588
rect 5460 8548 5488 8576
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 5276 8520 5488 8548
rect 5736 8520 6561 8548
rect 5276 8492 5304 8520
rect 5258 8440 5264 8492
rect 5316 8440 5322 8492
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5736 8489 5764 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6840 8548 6868 8576
rect 6840 8520 7144 8548
rect 6549 8511 6607 8517
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5684 8452 5733 8480
rect 5684 8440 5690 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6512 8452 6745 8480
rect 6512 8440 6518 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6638 8412 6644 8424
rect 6052 8384 6644 8412
rect 6052 8372 6058 8384
rect 6638 8372 6644 8384
rect 6696 8412 6702 8424
rect 6840 8412 6868 8443
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7116 8489 7144 8520
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 11946 8551 12004 8557
rect 11946 8548 11958 8551
rect 10560 8520 11958 8548
rect 10560 8508 10566 8520
rect 11946 8517 11958 8520
rect 11992 8517 12004 8551
rect 11946 8511 12004 8517
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 12216 8520 15393 8548
rect 12216 8508 12222 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15488 8548 15516 8588
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 16114 8616 16120 8628
rect 15887 8588 16120 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 16908 8588 17877 8616
rect 16908 8576 16914 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 19334 8616 19340 8628
rect 18012 8588 19340 8616
rect 18012 8576 18018 8588
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19886 8616 19892 8628
rect 19444 8588 19892 8616
rect 19444 8548 19472 8588
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20990 8616 20996 8628
rect 20272 8588 20996 8616
rect 15488 8520 19472 8548
rect 19521 8551 19579 8557
rect 15381 8511 15439 8517
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 20272 8548 20300 8588
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 23566 8616 23572 8628
rect 22060 8588 23572 8616
rect 22060 8576 22066 8588
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 25130 8616 25136 8628
rect 24912 8588 25136 8616
rect 24912 8576 24918 8588
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25590 8576 25596 8628
rect 25648 8616 25654 8628
rect 25866 8616 25872 8628
rect 25648 8588 25872 8616
rect 25648 8576 25654 8588
rect 25866 8576 25872 8588
rect 25924 8616 25930 8628
rect 26145 8619 26203 8625
rect 26145 8616 26157 8619
rect 25924 8588 26157 8616
rect 25924 8576 25930 8588
rect 26145 8585 26157 8588
rect 26191 8585 26203 8619
rect 26145 8579 26203 8585
rect 19567 8520 20300 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 20404 8520 20729 8548
rect 20404 8508 20410 8520
rect 20717 8517 20729 8520
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 22986 8551 23044 8557
rect 22986 8548 22998 8551
rect 20864 8520 22998 8548
rect 20864 8508 20870 8520
rect 22986 8517 22998 8520
rect 23032 8517 23044 8551
rect 22986 8511 23044 8517
rect 24946 8508 24952 8560
rect 25004 8548 25010 8560
rect 25004 8520 25075 8548
rect 25004 8508 25010 8520
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6972 8452 7021 8480
rect 6972 8440 6978 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 6696 8384 6868 8412
rect 6696 8372 6702 8384
rect 5534 8304 5540 8356
rect 5592 8304 5598 8356
rect 5629 8347 5687 8353
rect 5629 8313 5641 8347
rect 5675 8344 5687 8347
rect 5718 8344 5724 8356
rect 5675 8316 5724 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 5718 8304 5724 8316
rect 5776 8344 5782 8356
rect 6546 8344 6552 8356
rect 5776 8316 6552 8344
rect 5776 8304 5782 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7668 8344 7696 8443
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11204 8452 11713 8480
rect 11204 8440 11210 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12986 8480 12992 8492
rect 12584 8452 12992 8480
rect 12584 8440 12590 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13998 8480 14004 8492
rect 13587 8452 14004 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 15654 8440 15660 8492
rect 15712 8440 15718 8492
rect 18046 8440 18052 8492
rect 18104 8440 18110 8492
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18322 8489 18328 8492
rect 18310 8483 18328 8489
rect 18310 8449 18322 8483
rect 18310 8443 18328 8449
rect 18322 8440 18328 8443
rect 18380 8440 18386 8492
rect 18782 8480 18788 8492
rect 18427 8473 18485 8479
rect 7760 8412 7788 8440
rect 18427 8439 18439 8473
rect 18473 8470 18485 8473
rect 18524 8470 18788 8480
rect 18473 8452 18788 8470
rect 18473 8442 18552 8452
rect 18473 8439 18485 8442
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 19705 8486 19763 8489
rect 19794 8486 19800 8492
rect 19705 8483 19800 8486
rect 19705 8449 19717 8483
rect 19751 8458 19800 8483
rect 19751 8449 19763 8458
rect 19705 8443 19763 8449
rect 19794 8440 19800 8458
rect 19852 8440 19858 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 20622 8480 20628 8492
rect 20579 8452 20628 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 25047 8489 25075 8520
rect 22741 8483 22799 8489
rect 22741 8480 22753 8483
rect 22612 8452 22753 8480
rect 22612 8440 22618 8452
rect 22741 8449 22753 8452
rect 22787 8480 22799 8483
rect 25032 8483 25090 8489
rect 22787 8452 24808 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 18427 8433 18485 8439
rect 24780 8424 24808 8452
rect 25032 8449 25044 8483
rect 25078 8480 25090 8483
rect 25590 8480 25596 8492
rect 25078 8452 25596 8480
rect 25078 8449 25090 8452
rect 25032 8443 25090 8449
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7760 8384 7941 8412
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9582 8412 9588 8424
rect 9272 8384 9588 8412
rect 9272 8372 9278 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 17494 8412 17500 8424
rect 15611 8384 17500 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 6932 8316 7696 8344
rect 7745 8347 7803 8353
rect 6932 8288 6960 8316
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 7791 8316 9628 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 9600 8276 9628 8316
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 13504 8316 15848 8344
rect 13504 8304 13510 8316
rect 10318 8276 10324 8288
rect 9600 8248 10324 8276
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 13630 8276 13636 8288
rect 10468 8248 13636 8276
rect 10468 8236 10474 8248
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13740 8285 13768 8316
rect 13725 8279 13783 8285
rect 13725 8245 13737 8279
rect 13771 8245 13783 8279
rect 13725 8239 13783 8245
rect 15654 8236 15660 8288
rect 15712 8236 15718 8288
rect 15820 8276 15848 8316
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 17126 8344 17132 8356
rect 16264 8316 17132 8344
rect 16264 8304 16270 8316
rect 17126 8304 17132 8316
rect 17184 8344 17190 8356
rect 17954 8344 17960 8356
rect 17184 8316 17960 8344
rect 17184 8304 17190 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 20162 8344 20168 8356
rect 18932 8316 19472 8344
rect 18932 8304 18938 8316
rect 19242 8276 19248 8288
rect 15820 8248 19248 8276
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 19444 8276 19472 8316
rect 19781 8316 20168 8344
rect 19781 8276 19809 8316
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 24118 8304 24124 8356
rect 24176 8304 24182 8356
rect 19444 8248 19809 8276
rect 19886 8236 19892 8288
rect 19944 8236 19950 8288
rect 22189 8279 22247 8285
rect 22189 8245 22201 8279
rect 22235 8276 22247 8279
rect 22554 8276 22560 8288
rect 22235 8248 22560 8276
rect 22235 8245 22247 8248
rect 22189 8239 22247 8245
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 27062 8276 27068 8288
rect 23440 8248 27068 8276
rect 23440 8236 23446 8248
rect 27062 8236 27068 8248
rect 27120 8236 27126 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8041 4583 8075
rect 4525 8035 4583 8041
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 4982 8072 4988 8084
rect 4755 8044 4988 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 4540 8004 4568 8035
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 18233 8075 18291 8081
rect 9548 8044 16252 8072
rect 9548 8032 9554 8044
rect 5350 8004 5356 8016
rect 4540 7976 5356 8004
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 11848 7976 12655 8004
rect 11848 7964 11854 7976
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6788 7908 7113 7936
rect 6788 7896 6794 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 12526 7936 12532 7948
rect 7101 7899 7159 7905
rect 10796 7908 12532 7936
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 992 7840 1777 7868
rect 992 7828 998 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4338 7868 4344 7880
rect 4295 7840 4344 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4338 7828 4344 7840
rect 4396 7868 4402 7880
rect 5074 7868 5080 7880
rect 4396 7840 5080 7868
rect 4396 7828 4402 7840
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6052 7840 6377 7868
rect 6052 7828 6058 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6512 7840 6561 7868
rect 6512 7828 6518 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9484 7871 9542 7877
rect 9484 7837 9496 7871
rect 9530 7868 9542 7871
rect 10686 7868 10692 7880
rect 9530 7840 10692 7868
rect 9530 7837 9542 7840
rect 9484 7831 9542 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 10796 7800 10824 7908
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12627 7936 12655 7976
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 13265 8007 13323 8013
rect 12952 7976 13125 8004
rect 12952 7964 12958 7976
rect 12627 7908 12940 7936
rect 12802 7877 12808 7880
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12769 7871 12808 7877
rect 12769 7837 12781 7871
rect 12769 7831 12808 7837
rect 6564 7772 10824 7800
rect 6564 7744 6592 7772
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 4246 7732 4252 7744
rect 1627 7704 4252 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6365 7735 6423 7741
rect 6365 7732 6377 7735
rect 5592 7704 6377 7732
rect 5592 7692 5598 7704
rect 6365 7701 6377 7704
rect 6411 7701 6423 7735
rect 6365 7695 6423 7701
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 10594 7692 10600 7744
rect 10652 7692 10658 7744
rect 12636 7732 12664 7831
rect 12802 7828 12808 7831
rect 12860 7828 12866 7880
rect 12912 7809 12940 7908
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13097 7877 13125 7976
rect 13265 7973 13277 8007
rect 13311 8004 13323 8007
rect 13354 8004 13360 8016
rect 13311 7976 13360 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 13086 7871 13144 7877
rect 13086 7837 13098 7871
rect 13132 7837 13144 7871
rect 13086 7831 13144 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13964 7840 14289 7868
rect 13964 7828 13970 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14533 7871 14591 7877
rect 14533 7868 14545 7871
rect 14424 7840 14545 7868
rect 14424 7828 14430 7840
rect 14533 7837 14545 7840
rect 14579 7837 14591 7871
rect 14533 7831 14591 7837
rect 15562 7828 15568 7880
rect 15620 7828 15626 7880
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 16224 7877 16252 8044
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18279 8044 20760 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 16574 8004 16580 8016
rect 16500 7976 16580 8004
rect 16210 7871 16268 7877
rect 16210 7837 16222 7871
rect 16256 7837 16268 7871
rect 16210 7831 16268 7837
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 16500 7877 16528 7976
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 19058 8004 19064 8016
rect 18248 7976 19064 8004
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16623 7871 16681 7877
rect 16623 7837 16635 7871
rect 16669 7868 16681 7871
rect 18248 7868 18276 7976
rect 19058 7964 19064 7976
rect 19116 7964 19122 8016
rect 20732 8004 20760 8044
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21177 8075 21235 8081
rect 21177 8072 21189 8075
rect 20864 8044 21189 8072
rect 20864 8032 20870 8044
rect 21177 8041 21189 8044
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 22278 8032 22284 8084
rect 22336 8032 22342 8084
rect 23198 8032 23204 8084
rect 23256 8072 23262 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 23256 8044 23397 8072
rect 23256 8032 23262 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 23385 8035 23443 8041
rect 27890 8032 27896 8084
rect 27948 8072 27954 8084
rect 28353 8075 28411 8081
rect 28353 8072 28365 8075
rect 27948 8044 28365 8072
rect 27948 8032 27954 8044
rect 28353 8041 28365 8044
rect 28399 8041 28411 8075
rect 28353 8035 28411 8041
rect 20898 8004 20904 8016
rect 20732 7976 20904 8004
rect 20898 7964 20904 7976
rect 20956 7964 20962 8016
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 23290 8004 23296 8016
rect 22152 7976 23296 8004
rect 22152 7964 22158 7976
rect 23290 7964 23296 7976
rect 23348 8004 23354 8016
rect 24302 8004 24308 8016
rect 23348 7976 24308 8004
rect 23348 7964 23354 7976
rect 24302 7964 24308 7976
rect 24360 7964 24366 8016
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7936 18475 7939
rect 18874 7936 18880 7948
rect 18463 7908 18880 7936
rect 18463 7905 18475 7908
rect 18417 7899 18475 7905
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 21600 7908 23060 7936
rect 21600 7896 21606 7908
rect 16669 7840 18276 7868
rect 18325 7871 18383 7877
rect 16669 7837 16681 7840
rect 16623 7831 16681 7837
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 12897 7803 12955 7809
rect 12897 7769 12909 7803
rect 12943 7800 12955 7803
rect 15580 7800 15608 7828
rect 12943 7772 15608 7800
rect 15672 7772 17080 7800
rect 12943 7769 12955 7772
rect 12897 7763 12955 7769
rect 15562 7732 15568 7744
rect 12636 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 15672 7741 15700 7772
rect 15657 7735 15715 7741
rect 15657 7701 15669 7735
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 15804 7704 16773 7732
rect 15804 7692 15810 7704
rect 16761 7701 16773 7704
rect 16807 7701 16819 7735
rect 17052 7732 17080 7772
rect 17126 7760 17132 7812
rect 17184 7800 17190 7812
rect 18230 7800 18236 7812
rect 17184 7772 18236 7800
rect 17184 7760 17190 7772
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 18340 7800 18368 7831
rect 18506 7828 18512 7880
rect 18564 7868 18570 7880
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18564 7840 18705 7868
rect 18564 7828 18570 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19760 7840 19809 7868
rect 19760 7828 19766 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 21818 7877 21824 7880
rect 21637 7871 21695 7877
rect 21637 7868 21649 7871
rect 19944 7840 21649 7868
rect 19944 7828 19950 7840
rect 21637 7837 21649 7840
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 21785 7871 21824 7877
rect 21785 7837 21797 7871
rect 21785 7831 21824 7837
rect 21818 7828 21824 7831
rect 21876 7828 21882 7880
rect 22094 7828 22100 7880
rect 22152 7877 22158 7880
rect 22152 7868 22160 7877
rect 22152 7840 22197 7868
rect 22152 7831 22160 7840
rect 22152 7828 22158 7831
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 22922 7877 22928 7880
rect 22889 7871 22928 7877
rect 22889 7837 22901 7871
rect 22889 7831 22928 7837
rect 22922 7828 22928 7831
rect 22980 7828 22986 7880
rect 23032 7868 23060 7908
rect 23206 7871 23264 7877
rect 23206 7868 23218 7871
rect 23032 7840 23218 7868
rect 23206 7837 23218 7840
rect 23252 7837 23264 7871
rect 23206 7831 23264 7837
rect 24854 7828 24860 7880
rect 24912 7868 24918 7880
rect 25041 7871 25099 7877
rect 25041 7868 25053 7871
rect 24912 7840 25053 7868
rect 24912 7828 24918 7840
rect 25041 7837 25053 7840
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 25308 7871 25366 7877
rect 25308 7837 25320 7871
rect 25354 7868 25366 7871
rect 25774 7868 25780 7880
rect 25354 7840 25780 7868
rect 25354 7837 25366 7840
rect 25308 7831 25366 7837
rect 25774 7828 25780 7840
rect 25832 7828 25838 7880
rect 26694 7828 26700 7880
rect 26752 7868 26758 7880
rect 26973 7871 27031 7877
rect 26973 7868 26985 7871
rect 26752 7840 26985 7868
rect 26752 7828 26758 7840
rect 26973 7837 26985 7840
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 20070 7809 20076 7812
rect 18340 7772 20024 7800
rect 17402 7732 17408 7744
rect 17052 7704 17408 7732
rect 16761 7695 16819 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 19058 7732 19064 7744
rect 18647 7704 19064 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 19996 7732 20024 7772
rect 20064 7763 20076 7809
rect 20128 7800 20134 7812
rect 20128 7772 20164 7800
rect 20070 7760 20076 7763
rect 20128 7760 20134 7772
rect 20622 7760 20628 7812
rect 20680 7800 20686 7812
rect 21913 7803 21971 7809
rect 21913 7800 21925 7803
rect 20680 7772 21925 7800
rect 20680 7760 20686 7772
rect 21913 7769 21925 7772
rect 21959 7769 21971 7803
rect 21913 7763 21971 7769
rect 22005 7803 22063 7809
rect 22005 7769 22017 7803
rect 22051 7769 22063 7803
rect 22005 7763 22063 7769
rect 20346 7732 20352 7744
rect 19996 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 22020 7732 22048 7763
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 23017 7803 23075 7809
rect 23017 7800 23029 7803
rect 22704 7772 23029 7800
rect 22704 7760 22710 7772
rect 23017 7769 23029 7772
rect 23063 7769 23075 7803
rect 23017 7763 23075 7769
rect 23109 7803 23167 7809
rect 23109 7769 23121 7803
rect 23155 7800 23167 7803
rect 23750 7800 23756 7812
rect 23155 7772 23756 7800
rect 23155 7769 23167 7772
rect 23109 7763 23167 7769
rect 23750 7760 23756 7772
rect 23808 7760 23814 7812
rect 26510 7760 26516 7812
rect 26568 7800 26574 7812
rect 27218 7803 27276 7809
rect 27218 7800 27230 7803
rect 26568 7772 27230 7800
rect 26568 7760 26574 7772
rect 27218 7769 27230 7772
rect 27264 7800 27276 7803
rect 27338 7800 27344 7812
rect 27264 7772 27344 7800
rect 27264 7769 27276 7772
rect 27218 7763 27276 7769
rect 27338 7760 27344 7772
rect 27396 7760 27402 7812
rect 26326 7732 26332 7744
rect 22020 7704 26332 7732
rect 26326 7692 26332 7704
rect 26384 7732 26390 7744
rect 26421 7735 26479 7741
rect 26421 7732 26433 7735
rect 26384 7704 26433 7732
rect 26384 7692 26390 7704
rect 26421 7701 26433 7704
rect 26467 7701 26479 7735
rect 26421 7695 26479 7701
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 8904 7500 10824 7528
rect 8904 7488 8910 7500
rect 5718 7460 5724 7472
rect 5644 7432 5724 7460
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3878 7392 3884 7404
rect 2915 7364 3884 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 5644 7401 5672 7432
rect 5718 7420 5724 7432
rect 5776 7460 5782 7472
rect 7190 7460 7196 7472
rect 5776 7432 7196 7460
rect 5776 7420 5782 7432
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 8564 7463 8622 7469
rect 8564 7460 8576 7463
rect 8352 7432 8576 7460
rect 8352 7420 8358 7432
rect 8564 7429 8576 7432
rect 8610 7460 8622 7463
rect 9122 7460 9128 7472
rect 8610 7432 9128 7460
rect 8610 7429 8622 7432
rect 8564 7423 8622 7429
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 9398 7420 9404 7472
rect 9456 7460 9462 7472
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9456 7432 10149 7460
rect 9456 7420 9462 7432
rect 10137 7429 10149 7432
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 10244 7432 10732 7460
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6086 7392 6092 7404
rect 5951 7364 6092 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 10244 7392 10272 7432
rect 8444 7364 10272 7392
rect 10321 7395 10379 7401
rect 8444 7352 8450 7364
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 7064 7296 8309 7324
rect 7064 7284 7070 7296
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 9674 7216 9680 7268
rect 9732 7216 9738 7268
rect 10336 7256 10364 7355
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10704 7401 10732 7432
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7361 10747 7395
rect 10796 7392 10824 7500
rect 12250 7488 12256 7540
rect 12308 7488 12314 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12759 7500 15792 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12268 7401 12296 7488
rect 12345 7463 12403 7469
rect 12345 7429 12357 7463
rect 12391 7460 12403 7463
rect 13078 7460 13084 7472
rect 12391 7432 13084 7460
rect 12391 7429 12403 7432
rect 12345 7423 12403 7429
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 13173 7463 13231 7469
rect 13173 7429 13185 7463
rect 13219 7429 13231 7463
rect 13173 7423 13231 7429
rect 12618 7401 12624 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 10796 7364 12081 7392
rect 10689 7355 10747 7361
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12217 7395 12296 7401
rect 12217 7361 12229 7395
rect 12263 7364 12296 7395
rect 12437 7395 12495 7401
rect 12263 7361 12275 7364
rect 12217 7355 12275 7361
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 12575 7395 12624 7401
rect 12575 7361 12587 7395
rect 12621 7361 12624 7395
rect 12575 7355 12624 7361
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 12452 7324 12480 7355
rect 12618 7352 12624 7355
rect 12676 7352 12682 7404
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 13188 7392 13216 7423
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 13373 7463 13431 7469
rect 13373 7460 13385 7463
rect 13320 7432 13385 7460
rect 13320 7420 13326 7432
rect 13373 7429 13385 7432
rect 13419 7429 13431 7463
rect 13373 7423 13431 7429
rect 14001 7463 14059 7469
rect 14001 7429 14013 7463
rect 14047 7460 14059 7463
rect 15378 7460 15384 7472
rect 14047 7432 15384 7460
rect 14047 7429 14059 7432
rect 14001 7423 14059 7429
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 13538 7392 13544 7404
rect 12860 7364 13544 7392
rect 12860 7352 12866 7364
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 15764 7401 15792 7500
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 20622 7528 20628 7540
rect 20088 7500 20628 7528
rect 17052 7460 17080 7488
rect 15948 7432 17080 7460
rect 15948 7401 15976 7432
rect 17126 7420 17132 7472
rect 17184 7420 17190 7472
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7460 17279 7463
rect 18966 7460 18972 7472
rect 17267 7432 18972 7460
rect 17267 7429 17279 7432
rect 17221 7423 17279 7429
rect 18966 7420 18972 7432
rect 19024 7460 19030 7472
rect 19886 7460 19892 7472
rect 19024 7432 19892 7460
rect 19024 7420 19030 7432
rect 19886 7420 19892 7432
rect 19944 7420 19950 7472
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17001 7395 17059 7401
rect 17001 7361 17013 7395
rect 17047 7392 17059 7395
rect 17047 7361 17080 7392
rect 17001 7355 17080 7361
rect 10836 7296 12480 7324
rect 12544 7296 13492 7324
rect 10836 7284 10842 7296
rect 12544 7256 12572 7296
rect 10336 7228 12572 7256
rect 12636 7228 13400 7256
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 2774 7188 2780 7200
rect 1627 7160 2780 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 2958 7148 2964 7200
rect 3016 7148 3022 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4798 7188 4804 7200
rect 4212 7160 4804 7188
rect 4212 7148 4218 7160
rect 4798 7148 4804 7160
rect 4856 7188 4862 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 4856 7160 5457 7188
rect 4856 7148 4862 7160
rect 5445 7157 5457 7160
rect 5491 7157 5503 7191
rect 5445 7151 5503 7157
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10376 7160 10609 7188
rect 10376 7148 10382 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10597 7151 10655 7157
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 12636 7188 12664 7228
rect 13372 7197 13400 7228
rect 10928 7160 12664 7188
rect 13357 7191 13415 7197
rect 10928 7148 10934 7160
rect 13357 7157 13369 7191
rect 13403 7157 13415 7191
rect 13464 7188 13492 7296
rect 14182 7284 14188 7336
rect 14240 7284 14246 7336
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16868 7324 16896 7355
rect 15344 7296 16896 7324
rect 17052 7324 17080 7355
rect 17310 7352 17316 7404
rect 17368 7401 17374 7404
rect 17368 7392 17376 7401
rect 17678 7392 17684 7404
rect 17368 7364 17684 7392
rect 17368 7355 17376 7364
rect 17368 7352 17374 7355
rect 17678 7352 17684 7364
rect 17736 7392 17742 7404
rect 18506 7392 18512 7404
rect 17736 7364 18512 7392
rect 17736 7352 17742 7364
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 19978 7392 19984 7404
rect 18831 7364 19984 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 17862 7324 17868 7336
rect 17052 7296 17868 7324
rect 15344 7284 15350 7296
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18601 7327 18659 7333
rect 18601 7293 18613 7327
rect 18647 7324 18659 7327
rect 18966 7324 18972 7336
rect 18647 7296 18972 7324
rect 18647 7293 18659 7296
rect 18601 7287 18659 7293
rect 18966 7284 18972 7296
rect 19024 7324 19030 7336
rect 19242 7324 19248 7336
rect 19024 7296 19248 7324
rect 19024 7284 19030 7296
rect 19242 7284 19248 7296
rect 19300 7284 19306 7336
rect 13541 7259 13599 7265
rect 13541 7225 13553 7259
rect 13587 7256 13599 7259
rect 14090 7256 14096 7268
rect 13587 7228 14096 7256
rect 13587 7225 13599 7228
rect 13541 7219 13599 7225
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 15194 7256 15200 7268
rect 14200 7228 15200 7256
rect 14200 7188 14228 7228
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 17954 7256 17960 7268
rect 15948 7228 17960 7256
rect 13464 7160 14228 7188
rect 13357 7151 13415 7157
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 15948 7197 15976 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 20088 7256 20116 7500
rect 20364 7469 20392 7500
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 22370 7528 22376 7540
rect 20763 7500 22376 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 23937 7531 23995 7537
rect 23937 7497 23949 7531
rect 23983 7528 23995 7531
rect 24210 7528 24216 7540
rect 23983 7500 24216 7528
rect 23983 7497 23995 7500
rect 23937 7491 23995 7497
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 26602 7488 26608 7540
rect 26660 7488 26666 7540
rect 20349 7463 20407 7469
rect 20349 7429 20361 7463
rect 20395 7429 20407 7463
rect 20349 7423 20407 7429
rect 20438 7420 20444 7472
rect 20496 7460 20502 7472
rect 22186 7460 22192 7472
rect 20496 7432 22192 7460
rect 20496 7420 20502 7432
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20180 7324 20208 7355
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20312 7364 20545 7392
rect 20312 7352 20318 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 22813 7395 22871 7401
rect 22813 7392 22825 7395
rect 21692 7364 22825 7392
rect 21692 7352 21698 7364
rect 22813 7361 22825 7364
rect 22859 7361 22871 7395
rect 22813 7355 22871 7361
rect 25038 7352 25044 7404
rect 25096 7392 25102 7404
rect 25492 7395 25550 7401
rect 25492 7392 25504 7395
rect 25096 7364 25504 7392
rect 25096 7352 25102 7364
rect 25492 7361 25504 7364
rect 25538 7392 25550 7395
rect 25866 7392 25872 7404
rect 25538 7364 25872 7392
rect 25538 7361 25550 7364
rect 25492 7355 25550 7361
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 20714 7324 20720 7336
rect 20180 7296 20720 7324
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 23566 7284 23572 7336
rect 23624 7324 23630 7336
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 23624 7296 25237 7324
rect 23624 7284 23630 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 24118 7256 24124 7268
rect 18984 7228 20116 7256
rect 23676 7228 24124 7256
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14424 7160 14473 7188
rect 14424 7148 14430 7160
rect 14461 7157 14473 7160
rect 14507 7157 14519 7191
rect 14461 7151 14519 7157
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 17402 7148 17408 7200
rect 17460 7188 17466 7200
rect 18984 7197 19012 7228
rect 18969 7191 19027 7197
rect 18969 7188 18981 7191
rect 17460 7160 18981 7188
rect 17460 7148 17466 7160
rect 18969 7157 18981 7160
rect 19015 7157 19027 7191
rect 18969 7151 19027 7157
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 23676 7188 23704 7228
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 19116 7160 23704 7188
rect 25240 7188 25268 7287
rect 27154 7188 27160 7200
rect 25240 7160 27160 7188
rect 19116 7148 19122 7160
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 9272 6956 9321 6984
rect 9272 6944 9278 6956
rect 9309 6953 9321 6956
rect 9355 6953 9367 6987
rect 9309 6947 9367 6953
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 10192 6956 12434 6984
rect 10192 6944 10198 6956
rect 5368 6888 6215 6916
rect 1578 6808 1584 6860
rect 1636 6808 1642 6860
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 5368 6848 5396 6888
rect 6086 6848 6092 6860
rect 3016 6820 5396 6848
rect 5460 6820 6092 6848
rect 3016 6808 3022 6820
rect 1848 6783 1906 6789
rect 1848 6749 1860 6783
rect 1894 6780 1906 6783
rect 2682 6780 2688 6792
rect 1894 6752 2688 6780
rect 1894 6749 1906 6752
rect 1848 6743 1906 6749
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 5460 6789 5488 6820
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6187 6848 6215 6888
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 10870 6916 10876 6928
rect 7708 6888 10876 6916
rect 7708 6876 7714 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 12066 6876 12072 6928
rect 12124 6876 12130 6928
rect 12406 6916 12434 6956
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13504 6956 13553 6984
rect 13504 6944 13510 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 14274 6944 14280 6996
rect 14332 6984 14338 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14332 6956 14473 6984
rect 14332 6944 14338 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 14461 6947 14519 6953
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 15620 6956 16681 6984
rect 15620 6944 15626 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 16669 6947 16727 6953
rect 20809 6987 20867 6993
rect 20809 6953 20821 6987
rect 20855 6953 20867 6987
rect 20809 6947 20867 6953
rect 14366 6916 14372 6928
rect 12406 6888 14372 6916
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 20824 6916 20852 6947
rect 21726 6944 21732 6996
rect 21784 6984 21790 6996
rect 21784 6956 23428 6984
rect 21784 6944 21790 6956
rect 16172 6888 20852 6916
rect 16172 6876 16178 6888
rect 21910 6876 21916 6928
rect 21968 6916 21974 6928
rect 22370 6916 22376 6928
rect 21968 6888 22376 6916
rect 21968 6876 21974 6888
rect 22370 6876 22376 6888
rect 22428 6916 22434 6928
rect 23290 6916 23296 6928
rect 22428 6888 23296 6916
rect 22428 6876 22434 6888
rect 23290 6876 23296 6888
rect 23348 6876 23354 6928
rect 23400 6916 23428 6956
rect 23934 6944 23940 6996
rect 23992 6984 23998 6996
rect 24029 6987 24087 6993
rect 24029 6984 24041 6987
rect 23992 6956 24041 6984
rect 23992 6944 23998 6956
rect 24029 6953 24041 6956
rect 24075 6953 24087 6987
rect 25130 6984 25136 6996
rect 24029 6947 24087 6953
rect 24136 6956 25136 6984
rect 24136 6916 24164 6956
rect 25130 6944 25136 6956
rect 25188 6984 25194 6996
rect 25188 6956 25820 6984
rect 25188 6944 25194 6956
rect 23400 6888 24164 6916
rect 25792 6916 25820 6956
rect 26234 6944 26240 6996
rect 26292 6944 26298 6996
rect 28077 6987 28135 6993
rect 28077 6984 28089 6987
rect 26344 6956 28089 6984
rect 26344 6916 26372 6956
rect 28077 6953 28089 6956
rect 28123 6953 28135 6987
rect 28077 6947 28135 6953
rect 25792 6888 26372 6916
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6187 6820 6469 6848
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 12084 6848 12112 6876
rect 6457 6811 6515 6817
rect 11716 6820 12112 6848
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 6472 6780 6500 6811
rect 7006 6780 7012 6792
rect 6472 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8996 6752 9137 6780
rect 8996 6740 9002 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 11716 6789 11744 6820
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 16206 6848 16212 6860
rect 12308 6820 14780 6848
rect 12308 6808 12314 6820
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11665 6783 11744 6789
rect 11665 6749 11677 6783
rect 11711 6752 11744 6783
rect 11711 6749 11723 6752
rect 11665 6743 11723 6749
rect 5629 6715 5687 6721
rect 5629 6681 5641 6715
rect 5675 6712 5687 6715
rect 5810 6712 5816 6724
rect 5675 6684 5816 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 6270 6672 6276 6724
rect 6328 6712 6334 6724
rect 6724 6715 6782 6721
rect 6724 6712 6736 6715
rect 6328 6684 6736 6712
rect 6328 6672 6334 6684
rect 6724 6681 6736 6684
rect 6770 6712 6782 6715
rect 7466 6712 7472 6724
rect 6770 6684 7472 6712
rect 6770 6681 6782 6684
rect 6724 6675 6782 6681
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3142 6644 3148 6656
rect 3007 6616 3148 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5350 6644 5356 6656
rect 4948 6616 5356 6644
rect 4948 6604 4954 6616
rect 5350 6604 5356 6616
rect 5408 6644 5414 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5408 6616 5549 6644
rect 5408 6604 5414 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5537 6607 5595 6613
rect 7837 6647 7895 6653
rect 7837 6613 7849 6647
rect 7883 6644 7895 6647
rect 8294 6644 8300 6656
rect 7883 6616 8300 6644
rect 7883 6613 7895 6616
rect 7837 6607 7895 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9858 6604 9864 6656
rect 9916 6604 9922 6656
rect 11532 6644 11560 6743
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 12023 6783 12081 6789
rect 12023 6749 12035 6783
rect 12069 6780 12081 6783
rect 12802 6780 12808 6792
rect 12069 6752 12808 6780
rect 12069 6749 12081 6752
rect 12023 6743 12081 6749
rect 12802 6740 12808 6752
rect 12860 6780 12866 6792
rect 14752 6789 14780 6820
rect 14936 6820 16212 6848
rect 14936 6789 14964 6820
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 16724 6820 17080 6848
rect 16724 6808 16730 6820
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 12860 6752 14657 6780
rect 12860 6740 12866 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15010 6740 15016 6792
rect 15068 6740 15074 6792
rect 15838 6740 15844 6792
rect 15896 6740 15902 6792
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 11882 6672 11888 6724
rect 11940 6672 11946 6724
rect 12526 6712 12532 6724
rect 11992 6684 12532 6712
rect 11992 6644 12020 6684
rect 12526 6672 12532 6684
rect 12584 6672 12590 6724
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 12768 6684 13369 6712
rect 12768 6672 12774 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 15948 6712 15976 6743
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16816 6752 16865 6780
rect 16816 6740 16822 6752
rect 16853 6749 16865 6752
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16942 6740 16948 6792
rect 17000 6740 17006 6792
rect 17052 6789 17080 6820
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 17276 6820 17325 6848
rect 17276 6808 17282 6820
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 17313 6811 17371 6817
rect 19306 6820 19441 6848
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 19306 6780 19334 6820
rect 19429 6817 19441 6820
rect 19475 6848 19487 6851
rect 20162 6848 20168 6860
rect 19475 6820 20168 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 21726 6848 21732 6860
rect 21560 6820 21732 6848
rect 17083 6752 19334 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 20254 6740 20260 6792
rect 20312 6740 20318 6792
rect 20622 6740 20628 6792
rect 20680 6789 20686 6792
rect 20680 6783 20707 6789
rect 20695 6749 20707 6783
rect 20680 6743 20707 6749
rect 20680 6740 20686 6743
rect 21174 6740 21180 6792
rect 21232 6774 21238 6792
rect 21560 6789 21588 6820
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 26326 6848 26332 6860
rect 25884 6820 26332 6848
rect 21269 6783 21327 6789
rect 21269 6774 21281 6783
rect 21232 6749 21281 6774
rect 21315 6749 21327 6783
rect 21232 6746 21327 6749
rect 21232 6740 21238 6746
rect 21269 6743 21327 6746
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21637 6783 21695 6789
rect 21637 6749 21649 6783
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 17155 6715 17213 6721
rect 17155 6712 17167 6715
rect 13357 6675 13415 6681
rect 13577 6684 15976 6712
rect 16132 6684 17167 6712
rect 13577 6656 13605 6684
rect 11532 6616 12020 6644
rect 12158 6604 12164 6656
rect 12216 6604 12222 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13538 6644 13544 6656
rect 13596 6653 13605 6656
rect 13596 6647 13620 6653
rect 12400 6616 13544 6644
rect 12400 6604 12406 6616
rect 13538 6604 13544 6616
rect 13608 6613 13620 6647
rect 13596 6607 13620 6613
rect 13596 6604 13602 6607
rect 13722 6604 13728 6656
rect 13780 6604 13786 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16132 6653 16160 6684
rect 17155 6681 17167 6684
rect 17201 6681 17213 6715
rect 17155 6675 17213 6681
rect 18690 6672 18696 6724
rect 18748 6712 18754 6724
rect 18966 6712 18972 6724
rect 18748 6684 18972 6712
rect 18748 6672 18754 6684
rect 18966 6672 18972 6684
rect 19024 6712 19030 6724
rect 20070 6712 20076 6724
rect 19024 6684 20076 6712
rect 19024 6672 19030 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20441 6715 20499 6721
rect 20441 6681 20453 6715
rect 20487 6681 20499 6715
rect 20441 6675 20499 6681
rect 16117 6647 16175 6653
rect 16117 6644 16129 6647
rect 15988 6616 16129 6644
rect 15988 6604 15994 6616
rect 16117 6613 16129 6616
rect 16163 6613 16175 6647
rect 16117 6607 16175 6613
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 19886 6604 19892 6656
rect 19944 6644 19950 6656
rect 20456 6644 20484 6675
rect 20530 6672 20536 6724
rect 20588 6672 20594 6724
rect 21453 6715 21511 6721
rect 21453 6712 21465 6715
rect 20640 6684 21465 6712
rect 20640 6644 20668 6684
rect 21453 6681 21465 6684
rect 21499 6681 21511 6715
rect 21652 6712 21680 6743
rect 21818 6740 21824 6792
rect 21876 6780 21882 6792
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 21876 6752 22293 6780
rect 21876 6740 21882 6752
rect 22281 6749 22293 6752
rect 22327 6749 22339 6783
rect 22281 6743 22339 6749
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6780 22523 6783
rect 22830 6780 22836 6792
rect 22511 6752 22836 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 22830 6740 22836 6752
rect 22888 6740 22894 6792
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6780 23535 6783
rect 23845 6783 23903 6789
rect 23523 6752 23612 6780
rect 23523 6749 23535 6752
rect 23477 6743 23535 6749
rect 21910 6712 21916 6724
rect 21652 6684 21916 6712
rect 21453 6675 21511 6681
rect 21910 6672 21916 6684
rect 21968 6672 21974 6724
rect 22649 6715 22707 6721
rect 22649 6681 22661 6715
rect 22695 6681 22707 6715
rect 22649 6675 22707 6681
rect 19944 6616 20668 6644
rect 19944 6604 19950 6616
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 21821 6647 21879 6653
rect 21821 6644 21833 6647
rect 20956 6616 21833 6644
rect 20956 6604 20962 6616
rect 21821 6613 21833 6616
rect 21867 6613 21879 6647
rect 22664 6644 22692 6675
rect 23474 6644 23480 6656
rect 22664 6616 23480 6644
rect 21821 6607 21879 6613
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 23584 6644 23612 6752
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24762 6780 24768 6792
rect 23891 6752 24768 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 24854 6740 24860 6792
rect 24912 6740 24918 6792
rect 25124 6783 25182 6789
rect 25124 6749 25136 6783
rect 25170 6780 25182 6783
rect 25884 6780 25912 6820
rect 26326 6808 26332 6820
rect 26384 6808 26390 6860
rect 26694 6808 26700 6860
rect 26752 6808 26758 6860
rect 26510 6780 26516 6792
rect 25170 6752 25912 6780
rect 26160 6752 26516 6780
rect 25170 6749 25182 6752
rect 25124 6743 25182 6749
rect 23658 6672 23664 6724
rect 23716 6672 23722 6724
rect 23753 6715 23811 6721
rect 23753 6681 23765 6715
rect 23799 6712 23811 6715
rect 26160 6712 26188 6752
rect 26510 6740 26516 6752
rect 26568 6740 26574 6792
rect 23799 6684 26188 6712
rect 23799 6681 23811 6684
rect 23753 6675 23811 6681
rect 26234 6672 26240 6724
rect 26292 6712 26298 6724
rect 26942 6715 27000 6721
rect 26942 6712 26954 6715
rect 26292 6684 26954 6712
rect 26292 6672 26298 6684
rect 26942 6681 26954 6684
rect 26988 6681 27000 6715
rect 26942 6675 27000 6681
rect 25038 6644 25044 6656
rect 23584 6616 25044 6644
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 4798 6440 4804 6452
rect 3007 6412 4804 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 5500 6412 5549 6440
rect 5500 6400 5506 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6641 6443 6699 6449
rect 6641 6440 6653 6443
rect 5960 6412 6653 6440
rect 5960 6400 5966 6412
rect 6641 6409 6653 6412
rect 6687 6409 6699 6443
rect 6641 6403 6699 6409
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8260 6412 13676 6440
rect 8260 6400 8266 6412
rect 1848 6375 1906 6381
rect 1848 6341 1860 6375
rect 1894 6372 1906 6375
rect 3694 6372 3700 6384
rect 1894 6344 3700 6372
rect 1894 6341 1906 6344
rect 1848 6335 1906 6341
rect 3694 6332 3700 6344
rect 3752 6332 3758 6384
rect 3878 6332 3884 6384
rect 3936 6372 3942 6384
rect 3936 6344 4568 6372
rect 3936 6332 3942 6344
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 2832 6276 3525 6304
rect 2832 6264 2838 6276
rect 3513 6273 3525 6276
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 4356 6100 4384 6267
rect 4540 6177 4568 6344
rect 5736 6344 6500 6372
rect 5736 6313 5764 6344
rect 6472 6316 6500 6344
rect 7374 6332 7380 6384
rect 7432 6372 7438 6384
rect 7552 6375 7610 6381
rect 7552 6372 7564 6375
rect 7432 6344 7564 6372
rect 7432 6332 7438 6344
rect 7552 6341 7564 6344
rect 7598 6372 7610 6375
rect 7650 6372 7656 6384
rect 7598 6344 7656 6372
rect 7598 6341 7610 6344
rect 7552 6335 7610 6341
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 9944 6375 10002 6381
rect 9944 6341 9956 6375
rect 9990 6372 10002 6375
rect 10594 6372 10600 6384
rect 9990 6344 10600 6372
rect 9990 6341 10002 6344
rect 9944 6335 10002 6341
rect 10594 6332 10600 6344
rect 10652 6372 10658 6384
rect 12250 6372 12256 6384
rect 10652 6344 12256 6372
rect 10652 6332 10658 6344
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6512 6276 6561 6304
rect 6512 6264 6518 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 6822 6304 6828 6316
rect 6779 6276 6828 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 6748 6236 6776 6267
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 8938 6304 8944 6316
rect 6932 6276 8944 6304
rect 5951 6208 6776 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 4525 6171 4583 6177
rect 4525 6137 4537 6171
rect 4571 6168 4583 6171
rect 6932 6168 6960 6276
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9272 6276 9689 6304
rect 9272 6264 9278 6276
rect 9677 6273 9689 6276
rect 9723 6304 9735 6307
rect 10410 6304 10416 6316
rect 9723 6276 10416 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 10410 6264 10416 6276
rect 10468 6304 10474 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 10468 6276 11713 6304
rect 10468 6264 10474 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11968 6307 12026 6313
rect 11968 6273 11980 6307
rect 12014 6304 12026 6307
rect 12342 6304 12348 6316
rect 12014 6276 12348 6304
rect 12014 6273 12026 6276
rect 11968 6267 12026 6273
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 13538 6264 13544 6316
rect 13596 6264 13602 6316
rect 13648 6313 13676 6412
rect 13832 6412 15148 6440
rect 13832 6381 13860 6412
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6341 13875 6375
rect 13817 6335 13875 6341
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 14458 6372 14464 6384
rect 13955 6344 14464 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 15120 6372 15148 6412
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 15712 6412 15761 6440
rect 15712 6400 15718 6412
rect 15749 6409 15761 6412
rect 15795 6409 15807 6443
rect 16390 6440 16396 6452
rect 15749 6403 15807 6409
rect 15847 6412 16396 6440
rect 15847 6372 15875 6412
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 17644 6412 20545 6440
rect 17644 6400 17650 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 22373 6443 22431 6449
rect 20533 6403 20591 6409
rect 21928 6412 22324 6440
rect 20898 6372 20904 6384
rect 15120 6344 15875 6372
rect 16316 6344 20904 6372
rect 13634 6307 13692 6313
rect 13634 6273 13646 6307
rect 13680 6273 13692 6307
rect 13634 6267 13692 6273
rect 14047 6307 14105 6313
rect 14047 6273 14059 6307
rect 14093 6304 14105 6307
rect 14550 6304 14556 6316
rect 14093 6276 14556 6304
rect 14093 6273 14105 6276
rect 14047 6267 14105 6273
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7064 6208 7297 6236
rect 7064 6196 7070 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 14752 6236 14780 6267
rect 14918 6264 14924 6316
rect 14976 6264 14982 6316
rect 15010 6264 15016 6316
rect 15068 6264 15074 6316
rect 15120 6313 15148 6344
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15344 6276 15945 6304
rect 15344 6264 15350 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 15654 6236 15660 6248
rect 14752 6208 15660 6236
rect 7285 6199 7343 6205
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 4571 6140 6960 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 15102 6128 15108 6180
rect 15160 6168 15166 6180
rect 16040 6168 16068 6267
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16316 6313 16344 6344
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 21928 6372 21956 6412
rect 22031 6375 22089 6381
rect 22031 6372 22043 6375
rect 21928 6344 22043 6372
rect 22031 6341 22043 6344
rect 22077 6341 22089 6375
rect 22205 6375 22263 6381
rect 22205 6372 22217 6375
rect 22031 6335 22089 6341
rect 22204 6341 22217 6372
rect 22251 6341 22263 6375
rect 22296 6372 22324 6412
rect 22373 6409 22385 6443
rect 22419 6440 22431 6443
rect 24578 6440 24584 6452
rect 22419 6412 24584 6440
rect 22419 6409 22431 6412
rect 22373 6403 22431 6409
rect 24578 6400 24584 6412
rect 24636 6400 24642 6452
rect 24670 6400 24676 6452
rect 24728 6400 24734 6452
rect 24762 6400 24768 6452
rect 24820 6440 24826 6452
rect 26050 6440 26056 6452
rect 24820 6412 26056 6440
rect 24820 6400 24826 6412
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 26418 6400 26424 6452
rect 26476 6440 26482 6452
rect 26513 6443 26571 6449
rect 26513 6440 26525 6443
rect 26476 6412 26525 6440
rect 26476 6400 26482 6412
rect 26513 6409 26525 6412
rect 26559 6409 26571 6443
rect 26513 6403 26571 6409
rect 23106 6372 23112 6384
rect 22296 6344 23112 6372
rect 22204 6335 22263 6341
rect 17586 6313 17592 6316
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 17580 6304 17592 6313
rect 17547 6276 17592 6304
rect 16301 6267 16359 6273
rect 17580 6267 17592 6276
rect 17586 6264 17592 6267
rect 17644 6264 17650 6316
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 19153 6307 19211 6313
rect 19153 6304 19165 6307
rect 18196 6276 19165 6304
rect 18196 6264 18202 6276
rect 19153 6273 19165 6276
rect 19199 6304 19211 6307
rect 19242 6304 19248 6316
rect 19199 6276 19248 6304
rect 19199 6273 19211 6276
rect 19153 6267 19211 6273
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 19420 6307 19478 6313
rect 19420 6273 19432 6307
rect 19466 6304 19478 6307
rect 20438 6304 20444 6316
rect 19466 6276 20444 6304
rect 19466 6273 19478 6276
rect 19420 6267 19478 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 22204 6304 22232 6335
rect 23106 6332 23112 6344
rect 23164 6332 23170 6384
rect 24688 6372 24716 6400
rect 25378 6375 25436 6381
rect 25378 6372 25390 6375
rect 24688 6344 25390 6372
rect 25378 6341 25390 6344
rect 25424 6341 25436 6375
rect 25378 6335 25436 6341
rect 23549 6307 23607 6313
rect 23549 6304 23561 6307
rect 20588 6276 22232 6304
rect 22756 6276 23561 6304
rect 20588 6264 20594 6276
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 15160 6140 16068 6168
rect 15160 6128 15166 6140
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 17328 6168 17356 6199
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 22756 6236 22784 6276
rect 23549 6273 23561 6276
rect 23595 6273 23607 6307
rect 23549 6267 23607 6273
rect 21600 6208 22784 6236
rect 23293 6239 23351 6245
rect 21600 6196 21606 6208
rect 23293 6205 23305 6239
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 16264 6140 17356 6168
rect 16264 6128 16270 6140
rect 20254 6128 20260 6180
rect 20312 6168 20318 6180
rect 22922 6168 22928 6180
rect 20312 6140 22928 6168
rect 20312 6128 20318 6140
rect 22922 6128 22928 6140
rect 22980 6128 22986 6180
rect 8294 6100 8300 6112
rect 3743 6072 8300 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9306 6100 9312 6112
rect 8720 6072 9312 6100
rect 8720 6060 8726 6072
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 13998 6100 14004 6112
rect 13127 6072 14004 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14182 6060 14188 6112
rect 14240 6060 14246 6112
rect 17494 6060 17500 6112
rect 17552 6100 17558 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 17552 6072 18705 6100
rect 17552 6060 17558 6072
rect 18693 6069 18705 6072
rect 18739 6100 18751 6103
rect 19334 6100 19340 6112
rect 18739 6072 19340 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 22189 6103 22247 6109
rect 22189 6069 22201 6103
rect 22235 6100 22247 6103
rect 22278 6100 22284 6112
rect 22235 6072 22284 6100
rect 22235 6069 22247 6072
rect 22189 6063 22247 6069
rect 22278 6060 22284 6072
rect 22336 6060 22342 6112
rect 23308 6100 23336 6199
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 24854 6236 24860 6248
rect 24636 6208 24860 6236
rect 24636 6196 24642 6208
rect 24854 6196 24860 6208
rect 24912 6236 24918 6248
rect 25130 6236 25136 6248
rect 24912 6208 25136 6236
rect 24912 6196 24918 6208
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 24578 6100 24584 6112
rect 23308 6072 24584 6100
rect 24578 6060 24584 6072
rect 24636 6060 24642 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3050 5896 3056 5908
rect 3007 5868 3056 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 3786 5896 3792 5908
rect 3375 5868 3792 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 1578 5720 1584 5772
rect 1636 5720 1642 5772
rect 1848 5695 1906 5701
rect 1848 5661 1860 5695
rect 1894 5692 1906 5695
rect 3344 5692 3372 5859
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 5166 5856 5172 5908
rect 5224 5856 5230 5908
rect 7006 5896 7012 5908
rect 6656 5868 7012 5896
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5760 4031 5763
rect 5350 5760 5356 5772
rect 4019 5732 5356 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 6656 5769 6684 5868
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8386 5896 8392 5908
rect 8067 5868 8392 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 1894 5664 3372 5692
rect 1894 5661 1906 5664
rect 1848 5655 1906 5661
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5442 5692 5448 5704
rect 5031 5664 5448 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 8036 5692 8064 5859
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 10502 5856 10508 5908
rect 10560 5856 10566 5908
rect 11793 5899 11851 5905
rect 11793 5865 11805 5899
rect 11839 5896 11851 5899
rect 13538 5896 13544 5908
rect 11839 5868 13544 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 15102 5896 15108 5908
rect 14332 5868 15108 5896
rect 14332 5856 14338 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15436 5868 15485 5896
rect 15436 5856 15442 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 18690 5856 18696 5908
rect 18748 5856 18754 5908
rect 18874 5856 18880 5908
rect 18932 5856 18938 5908
rect 20180 5868 21220 5896
rect 12802 5788 12808 5840
rect 12860 5788 12866 5840
rect 13262 5788 13268 5840
rect 13320 5828 13326 5840
rect 13906 5828 13912 5840
rect 13320 5800 13912 5828
rect 13320 5788 13326 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 14642 5828 14648 5840
rect 14056 5800 14648 5828
rect 14056 5788 14062 5800
rect 14642 5788 14648 5800
rect 14700 5788 14706 5840
rect 15930 5828 15936 5840
rect 15120 5800 15936 5828
rect 9122 5720 9128 5772
rect 9180 5720 9186 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13722 5760 13728 5772
rect 12492 5732 13728 5760
rect 12492 5720 12498 5732
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 5776 5664 8064 5692
rect 5776 5652 5782 5664
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9381 5695 9439 5701
rect 9381 5692 9393 5695
rect 9088 5686 9168 5692
rect 9324 5686 9393 5692
rect 9088 5664 9393 5686
rect 9088 5652 9094 5664
rect 9140 5658 9352 5664
rect 9381 5661 9393 5664
rect 9427 5661 9439 5695
rect 9381 5655 9439 5661
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11348 5664 11529 5692
rect 4801 5627 4859 5633
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 5534 5624 5540 5636
rect 4847 5596 5540 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 5534 5584 5540 5596
rect 5592 5584 5598 5636
rect 6908 5627 6966 5633
rect 6908 5593 6920 5627
rect 6954 5624 6966 5627
rect 7098 5624 7104 5636
rect 6954 5596 7104 5624
rect 6954 5593 6966 5596
rect 6908 5587 6966 5593
rect 7098 5584 7104 5596
rect 7156 5624 7162 5636
rect 7558 5624 7564 5636
rect 7156 5596 7564 5624
rect 7156 5584 7162 5596
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 11348 5624 11376 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 12066 5692 12072 5704
rect 11655 5664 12072 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 13170 5692 13176 5704
rect 12667 5664 13176 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 9646 5596 11376 5624
rect 11425 5627 11483 5633
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3878 5556 3884 5568
rect 2832 5528 3884 5556
rect 2832 5516 2838 5528
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9646 5556 9674 5596
rect 11425 5593 11437 5627
rect 11471 5624 11483 5627
rect 11698 5624 11704 5636
rect 11471 5596 11704 5624
rect 11471 5593 11483 5596
rect 11425 5587 11483 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 12636 5624 12664 5655
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13354 5652 13360 5704
rect 13412 5652 13418 5704
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 13630 5692 13636 5704
rect 13495 5664 13636 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 13630 5652 13636 5664
rect 13688 5692 13694 5704
rect 13906 5692 13912 5704
rect 13688 5664 13912 5692
rect 13688 5652 13694 5664
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 15010 5701 15016 5704
rect 14977 5695 15016 5701
rect 14977 5661 14989 5695
rect 14977 5655 15016 5661
rect 15010 5652 15016 5655
rect 15068 5652 15074 5704
rect 15120 5701 15148 5800
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 17957 5831 18015 5837
rect 17957 5797 17969 5831
rect 18003 5828 18015 5831
rect 20180 5828 20208 5868
rect 18003 5800 20208 5828
rect 18003 5797 18015 5800
rect 17957 5791 18015 5797
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 18782 5760 18788 5772
rect 15436 5732 18788 5760
rect 15436 5720 15442 5732
rect 18782 5720 18788 5732
rect 18840 5720 18846 5772
rect 19242 5720 19248 5772
rect 19300 5760 19306 5772
rect 19702 5760 19708 5772
rect 19300 5732 19708 5760
rect 19300 5720 19306 5732
rect 19702 5720 19708 5732
rect 19760 5760 19766 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19760 5732 20177 5760
rect 19760 5720 19766 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 21192 5760 21220 5868
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 21545 5899 21603 5905
rect 21545 5896 21557 5899
rect 21508 5868 21557 5896
rect 21508 5856 21514 5868
rect 21545 5865 21557 5868
rect 21591 5865 21603 5899
rect 21545 5859 21603 5865
rect 22557 5899 22615 5905
rect 22557 5865 22569 5899
rect 22603 5896 22615 5899
rect 22738 5896 22744 5908
rect 22603 5868 22744 5896
rect 22603 5865 22615 5868
rect 22557 5859 22615 5865
rect 22738 5856 22744 5868
rect 22796 5856 22802 5908
rect 25590 5856 25596 5908
rect 25648 5896 25654 5908
rect 25961 5899 26019 5905
rect 25961 5896 25973 5899
rect 25648 5868 25973 5896
rect 25648 5856 25654 5868
rect 25961 5865 25973 5868
rect 26007 5865 26019 5899
rect 25961 5859 26019 5865
rect 22462 5760 22468 5772
rect 21192 5732 22468 5760
rect 20165 5723 20223 5729
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 24578 5720 24584 5772
rect 24636 5720 24642 5772
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 15286 5652 15292 5704
rect 15344 5701 15350 5704
rect 15344 5692 15352 5701
rect 15344 5664 15389 5692
rect 15344 5655 15352 5664
rect 15344 5652 15350 5655
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 17770 5652 17776 5704
rect 17828 5652 17834 5704
rect 21358 5692 21364 5704
rect 18432 5664 21364 5692
rect 12216 5596 12664 5624
rect 12216 5584 12222 5596
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 15197 5627 15255 5633
rect 15197 5624 15209 5627
rect 14056 5596 15209 5624
rect 14056 5584 14062 5596
rect 15197 5593 15209 5596
rect 15243 5593 15255 5627
rect 15197 5587 15255 5593
rect 16574 5584 16580 5636
rect 16632 5584 16638 5636
rect 17586 5584 17592 5636
rect 17644 5584 17650 5636
rect 17678 5584 17684 5636
rect 17736 5584 17742 5636
rect 9364 5528 9674 5556
rect 9364 5516 9370 5528
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 13633 5559 13691 5565
rect 13633 5556 13645 5559
rect 12768 5528 13645 5556
rect 12768 5516 12774 5528
rect 13633 5525 13645 5528
rect 13679 5525 13691 5559
rect 13633 5519 13691 5525
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 18432 5556 18460 5664
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 22005 5695 22063 5701
rect 22005 5692 22017 5695
rect 21692 5664 22017 5692
rect 21692 5652 21698 5664
rect 22005 5661 22017 5664
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 26510 5692 26516 5704
rect 24780 5664 26516 5692
rect 18509 5627 18567 5633
rect 18509 5593 18521 5627
rect 18555 5624 18567 5627
rect 18966 5624 18972 5636
rect 18555 5596 18972 5624
rect 18555 5593 18567 5596
rect 18509 5587 18567 5593
rect 18966 5584 18972 5596
rect 19024 5584 19030 5636
rect 20432 5627 20490 5633
rect 20432 5593 20444 5627
rect 20478 5624 20490 5627
rect 21174 5624 21180 5636
rect 20478 5596 21180 5624
rect 20478 5593 20490 5596
rect 20432 5587 20490 5593
rect 21174 5584 21180 5596
rect 21232 5624 21238 5636
rect 21232 5596 21404 5624
rect 21232 5584 21238 5596
rect 16724 5528 18460 5556
rect 18719 5559 18777 5565
rect 16724 5516 16730 5528
rect 18719 5525 18731 5559
rect 18765 5556 18777 5559
rect 19610 5556 19616 5568
rect 18765 5528 19616 5556
rect 18765 5525 18777 5528
rect 18719 5519 18777 5525
rect 19610 5516 19616 5528
rect 19668 5556 19674 5568
rect 20530 5556 20536 5568
rect 19668 5528 20536 5556
rect 19668 5516 19674 5528
rect 20530 5516 20536 5528
rect 20588 5516 20594 5568
rect 21376 5556 21404 5596
rect 21450 5584 21456 5636
rect 21508 5624 21514 5636
rect 22189 5627 22247 5633
rect 22189 5624 22201 5627
rect 21508 5596 22201 5624
rect 21508 5584 21514 5596
rect 22189 5593 22201 5596
rect 22235 5593 22247 5627
rect 22189 5587 22247 5593
rect 22281 5627 22339 5633
rect 22281 5593 22293 5627
rect 22327 5624 22339 5627
rect 24780 5624 24808 5664
rect 26510 5652 26516 5664
rect 26568 5652 26574 5704
rect 26973 5695 27031 5701
rect 26973 5692 26985 5695
rect 26620 5664 26985 5692
rect 22327 5596 24808 5624
rect 24848 5627 24906 5633
rect 22327 5593 22339 5596
rect 22281 5587 22339 5593
rect 24848 5593 24860 5627
rect 24894 5593 24906 5627
rect 24848 5587 24906 5593
rect 24026 5556 24032 5568
rect 21376 5528 24032 5556
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 24118 5516 24124 5568
rect 24176 5556 24182 5568
rect 24863 5556 24891 5587
rect 25222 5584 25228 5636
rect 25280 5624 25286 5636
rect 26620 5624 26648 5664
rect 26973 5661 26985 5664
rect 27019 5661 27031 5695
rect 26973 5655 27031 5661
rect 25280 5596 26648 5624
rect 25280 5584 25286 5596
rect 26786 5584 26792 5636
rect 26844 5624 26850 5636
rect 27218 5627 27276 5633
rect 27218 5624 27230 5627
rect 26844 5596 27230 5624
rect 26844 5584 26850 5596
rect 27218 5593 27230 5596
rect 27264 5593 27276 5627
rect 27218 5587 27276 5593
rect 24176 5528 24891 5556
rect 24176 5516 24182 5528
rect 26510 5516 26516 5568
rect 26568 5556 26574 5568
rect 28353 5559 28411 5565
rect 28353 5556 28365 5559
rect 26568 5528 28365 5556
rect 26568 5516 26574 5528
rect 28353 5525 28365 5528
rect 28399 5525 28411 5559
rect 28353 5519 28411 5525
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 2774 5352 2780 5364
rect 1964 5324 2780 5352
rect 1964 5225 1992 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3050 5352 3056 5364
rect 2884 5324 3056 5352
rect 2884 5284 2912 5324
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6270 5352 6276 5364
rect 6043 5324 6276 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 9088 5324 9321 5352
rect 9088 5312 9094 5324
rect 9309 5321 9321 5324
rect 9355 5352 9367 5355
rect 9490 5352 9496 5364
rect 9355 5324 9496 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 12342 5352 12348 5364
rect 11195 5324 12348 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12526 5312 12532 5364
rect 12584 5312 12590 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15252 5324 15577 5352
rect 15252 5312 15258 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 15565 5315 15623 5321
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 20806 5352 20812 5364
rect 19567 5324 20812 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 26234 5312 26240 5364
rect 26292 5352 26298 5364
rect 26605 5355 26663 5361
rect 26605 5352 26617 5355
rect 26292 5324 26617 5352
rect 26292 5312 26298 5324
rect 26605 5321 26617 5324
rect 26651 5321 26663 5355
rect 26605 5315 26663 5321
rect 2700 5256 2912 5284
rect 2700 5225 2728 5256
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2884 5216 2912 5256
rect 2952 5287 3010 5293
rect 2952 5253 2964 5287
rect 2998 5284 3010 5287
rect 5166 5284 5172 5296
rect 2998 5256 5172 5284
rect 2998 5253 3010 5256
rect 2952 5247 3010 5253
rect 5166 5244 5172 5256
rect 5224 5284 5230 5296
rect 5224 5256 12020 5284
rect 5224 5244 5230 5256
rect 4062 5216 4068 5228
rect 2884 5188 4068 5216
rect 2685 5179 2743 5185
rect 4062 5176 4068 5188
rect 4120 5216 4126 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4120 5188 4629 5216
rect 4120 5176 4126 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4884 5219 4942 5225
rect 4884 5185 4896 5219
rect 4930 5216 4942 5219
rect 6822 5216 6828 5228
rect 4930 5188 6828 5216
rect 4930 5185 4942 5188
rect 4884 5179 4942 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8202 5225 8208 5228
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7064 5188 7941 5216
rect 7064 5176 7070 5188
rect 7929 5185 7941 5188
rect 7975 5185 7987 5219
rect 8196 5216 8208 5225
rect 8163 5188 8208 5216
rect 7929 5179 7987 5185
rect 8196 5179 8208 5188
rect 8202 5176 8208 5179
rect 8260 5176 8266 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 9858 5216 9864 5228
rect 9815 5188 9864 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 11992 5225 12020 5256
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 12124 5256 12173 5284
rect 12124 5244 12130 5256
rect 12161 5253 12173 5256
rect 12207 5284 12219 5287
rect 12434 5284 12440 5296
rect 12207 5256 12440 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 13532 5287 13590 5293
rect 13532 5253 13544 5287
rect 13578 5284 13590 5287
rect 14274 5284 14280 5296
rect 13578 5256 14280 5284
rect 13578 5253 13590 5256
rect 13532 5247 13590 5253
rect 14274 5244 14280 5256
rect 14332 5244 14338 5296
rect 15286 5244 15292 5296
rect 15344 5284 15350 5296
rect 17221 5287 17279 5293
rect 17221 5284 17233 5287
rect 15344 5256 17233 5284
rect 15344 5244 15350 5256
rect 17221 5253 17233 5256
rect 17267 5253 17279 5287
rect 17221 5247 17279 5253
rect 18230 5244 18236 5296
rect 18288 5284 18294 5296
rect 18414 5293 18420 5296
rect 18408 5284 18420 5293
rect 18288 5256 18420 5284
rect 18288 5244 18294 5256
rect 18408 5247 18420 5256
rect 18414 5244 18420 5247
rect 18472 5244 18478 5296
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 19981 5287 20039 5293
rect 19981 5284 19993 5287
rect 19116 5256 19993 5284
rect 19116 5244 19122 5256
rect 19981 5253 19993 5256
rect 20027 5253 20039 5287
rect 19981 5247 20039 5253
rect 20197 5287 20255 5293
rect 20197 5253 20209 5287
rect 20243 5284 20255 5287
rect 22830 5284 22836 5296
rect 20243 5256 22836 5284
rect 20243 5253 20255 5256
rect 20197 5247 20255 5253
rect 22830 5244 22836 5256
rect 22888 5244 22894 5296
rect 24486 5244 24492 5296
rect 24544 5284 24550 5296
rect 25470 5287 25528 5293
rect 25470 5284 25482 5287
rect 24544 5256 25482 5284
rect 24544 5244 24550 5256
rect 25470 5253 25482 5256
rect 25516 5284 25528 5287
rect 27798 5284 27804 5296
rect 25516 5256 27804 5284
rect 25516 5253 25528 5256
rect 25470 5247 25528 5253
rect 27798 5244 27804 5256
rect 27856 5244 27862 5296
rect 10036 5219 10094 5225
rect 10036 5185 10048 5219
rect 10082 5216 10094 5219
rect 11977 5219 12035 5225
rect 10082 5188 11284 5216
rect 10082 5185 10094 5188
rect 10036 5179 10094 5185
rect 6178 5080 6184 5092
rect 5920 5052 6184 5080
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 3786 5012 3792 5024
rect 2179 4984 3792 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 5920 5012 5948 5052
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 4111 4984 5948 5012
rect 11256 5012 11284 5188
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12618 5216 12624 5228
rect 12391 5188 12624 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12618 5176 12624 5188
rect 12676 5216 12682 5228
rect 12986 5216 12992 5228
rect 12676 5188 12992 5216
rect 12676 5176 12682 5188
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13262 5176 13268 5228
rect 13320 5176 13326 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 13872 5188 15117 5216
rect 13872 5176 13878 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15746 5216 15752 5228
rect 15427 5188 15752 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16666 5216 16672 5228
rect 16163 5188 16672 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16816 5188 17049 5216
rect 16816 5176 16822 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 19076 5216 19104 5244
rect 17037 5179 17095 5185
rect 17512 5188 19104 5216
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5148 15347 5151
rect 16298 5148 16304 5160
rect 15335 5120 16304 5148
rect 15335 5117 15347 5120
rect 15289 5111 15347 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17512 5148 17540 5188
rect 25222 5176 25228 5228
rect 25280 5176 25286 5228
rect 26418 5176 26424 5228
rect 26476 5216 26482 5228
rect 27433 5219 27491 5225
rect 27433 5216 27445 5219
rect 26476 5188 27445 5216
rect 26476 5176 26482 5188
rect 27433 5185 27445 5188
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 16899 5120 17540 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 20162 5108 20168 5160
rect 20220 5148 20226 5160
rect 24394 5148 24400 5160
rect 20220 5120 24400 5148
rect 20220 5108 20226 5120
rect 24394 5108 24400 5120
rect 24452 5108 24458 5160
rect 27154 5108 27160 5160
rect 27212 5108 27218 5160
rect 17954 5080 17960 5092
rect 15396 5052 17960 5080
rect 14550 5012 14556 5024
rect 11256 4984 14556 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 14550 4972 14556 4984
rect 14608 5012 14614 5024
rect 15396 5021 15424 5052
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 14608 4984 14657 5012
rect 14608 4972 14614 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 14645 4975 14703 4981
rect 15381 5015 15439 5021
rect 15381 4981 15393 5015
rect 15427 4981 15439 5015
rect 15381 4975 15439 4981
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16390 5012 16396 5024
rect 16264 4984 16396 5012
rect 16264 4972 16270 4984
rect 16390 4972 16396 4984
rect 16448 5012 16454 5024
rect 18156 5012 18184 5108
rect 22462 5080 22468 5092
rect 20180 5052 22468 5080
rect 20180 5021 20208 5052
rect 22462 5040 22468 5052
rect 22520 5040 22526 5092
rect 16448 4984 18184 5012
rect 20165 5015 20223 5021
rect 16448 4972 16454 4984
rect 20165 4981 20177 5015
rect 20211 4981 20223 5015
rect 20165 4975 20223 4981
rect 20346 4972 20352 5024
rect 20404 4972 20410 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4808 5963 4811
rect 7098 4808 7104 4820
rect 5951 4780 7104 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 10778 4768 10784 4820
rect 10836 4768 10842 4820
rect 12526 4808 12532 4820
rect 12360 4780 12532 4808
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1636 4644 1777 4672
rect 1636 4632 1642 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 1765 4635 1823 4641
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4120 4644 4537 4672
rect 4120 4632 4126 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 12360 4681 12388 4780
rect 12526 4768 12532 4780
rect 12584 4808 12590 4820
rect 13262 4808 13268 4820
rect 12584 4780 13268 4808
rect 12584 4768 12590 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13725 4811 13783 4817
rect 13725 4777 13737 4811
rect 13771 4808 13783 4811
rect 14274 4808 14280 4820
rect 13771 4780 14280 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14700 4780 14841 4808
rect 14700 4768 14706 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 16758 4808 16764 4820
rect 14829 4771 14887 4777
rect 15111 4780 16764 4808
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 15013 4743 15071 4749
rect 15013 4740 15025 4743
rect 14792 4712 15025 4740
rect 14792 4700 14798 4712
rect 15013 4709 15025 4712
rect 15059 4709 15071 4743
rect 15013 4703 15071 4709
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 10468 4644 12357 4672
rect 10468 4632 10474 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 2021 4607 2079 4613
rect 2021 4604 2033 4607
rect 1544 4576 2033 4604
rect 1544 4564 1550 4576
rect 2021 4573 2033 4576
rect 2067 4573 2079 4607
rect 2021 4567 2079 4573
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 7156 4576 7205 4604
rect 7156 4564 7162 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7460 4607 7518 4613
rect 7460 4573 7472 4607
rect 7506 4604 7518 4607
rect 8662 4604 8668 4616
rect 7506 4576 8668 4604
rect 7506 4573 7518 4576
rect 7460 4567 7518 4573
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9950 4604 9956 4616
rect 9447 4576 9956 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9950 4564 9956 4576
rect 10008 4604 10014 4616
rect 10870 4604 10876 4616
rect 10008 4576 10876 4604
rect 10008 4564 10014 4576
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 15111 4604 15139 4780
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 20162 4808 20168 4820
rect 18279 4780 20168 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21542 4768 21548 4820
rect 21600 4808 21606 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21600 4780 21925 4808
rect 21600 4768 21606 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 21913 4771 21971 4777
rect 24026 4768 24032 4820
rect 24084 4768 24090 4820
rect 25958 4768 25964 4820
rect 26016 4768 26022 4820
rect 27798 4768 27804 4820
rect 27856 4768 27862 4820
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 16724 4712 18429 4740
rect 16724 4700 16730 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 19518 4700 19524 4752
rect 19576 4740 19582 4752
rect 20073 4743 20131 4749
rect 20073 4740 20085 4743
rect 19576 4712 20085 4740
rect 19576 4700 19582 4712
rect 20073 4709 20085 4712
rect 20119 4709 20131 4743
rect 20073 4703 20131 4709
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 18966 4672 18972 4684
rect 18104 4644 18972 4672
rect 18104 4632 18110 4644
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19812 4644 20484 4672
rect 14844 4576 15139 4604
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 4770 4539 4828 4545
rect 4770 4536 4782 4539
rect 4304 4508 4782 4536
rect 4304 4496 4310 4508
rect 4770 4505 4782 4508
rect 4816 4505 4828 4539
rect 4770 4499 4828 4505
rect 9668 4539 9726 4545
rect 9668 4505 9680 4539
rect 9714 4536 9726 4539
rect 11054 4536 11060 4548
rect 9714 4508 11060 4536
rect 9714 4505 9726 4508
rect 9668 4499 9726 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 12618 4545 12624 4548
rect 12612 4536 12624 4545
rect 12579 4508 12624 4536
rect 12612 4499 12624 4508
rect 12618 4496 12624 4499
rect 12676 4496 12682 4548
rect 14090 4496 14096 4548
rect 14148 4536 14154 4548
rect 14844 4545 14872 4576
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 15838 4613 15844 4616
rect 15832 4567 15844 4613
rect 15896 4604 15902 4616
rect 15896 4576 18552 4604
rect 15838 4564 15844 4567
rect 15896 4564 15902 4576
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 14148 4508 14657 4536
rect 14148 4496 14154 4508
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 14844 4539 14903 4545
rect 14844 4508 14857 4539
rect 14645 4499 14703 4505
rect 14845 4505 14857 4508
rect 14891 4505 14903 4539
rect 17402 4536 17408 4548
rect 14845 4499 14903 4505
rect 14936 4508 17408 4536
rect 8570 4428 8576 4480
rect 8628 4428 8634 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 14936 4468 14964 4508
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 18046 4496 18052 4548
rect 18104 4496 18110 4548
rect 18138 4496 18144 4548
rect 18196 4536 18202 4548
rect 18249 4539 18307 4545
rect 18249 4536 18261 4539
rect 18196 4508 18261 4536
rect 18196 4496 18202 4508
rect 18249 4505 18261 4508
rect 18295 4505 18307 4539
rect 18249 4499 18307 4505
rect 10560 4440 14964 4468
rect 10560 4428 10566 4440
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16816 4440 16957 4468
rect 16816 4428 16822 4440
rect 16945 4437 16957 4440
rect 16991 4468 17003 4471
rect 17770 4468 17776 4480
rect 16991 4440 17776 4468
rect 16991 4437 17003 4440
rect 16945 4431 17003 4437
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18524 4468 18552 4576
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19577 4607 19635 4613
rect 19577 4573 19589 4607
rect 19623 4604 19635 4607
rect 19812 4604 19840 4644
rect 19623 4576 19840 4604
rect 19623 4573 19635 4576
rect 19577 4567 19635 4573
rect 19886 4564 19892 4616
rect 19944 4613 19950 4616
rect 19944 4604 19952 4613
rect 19944 4576 19989 4604
rect 19944 4567 19952 4576
rect 19944 4564 19950 4567
rect 19702 4496 19708 4548
rect 19760 4496 19766 4548
rect 19797 4539 19855 4545
rect 19797 4505 19809 4539
rect 19843 4505 19855 4539
rect 19797 4499 19855 4505
rect 19812 4468 19840 4499
rect 18524 4440 19840 4468
rect 20456 4468 20484 4644
rect 24302 4632 24308 4684
rect 24360 4672 24366 4684
rect 24360 4644 24716 4672
rect 24360 4632 24366 4644
rect 20530 4564 20536 4616
rect 20588 4564 20594 4616
rect 22922 4613 22928 4616
rect 20800 4607 20858 4613
rect 20800 4604 20812 4607
rect 20732 4576 20812 4604
rect 20732 4548 20760 4576
rect 20800 4573 20812 4576
rect 20846 4573 20858 4607
rect 20800 4567 20858 4573
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4573 22707 4607
rect 22916 4604 22928 4613
rect 22883 4576 22928 4604
rect 22649 4567 22707 4573
rect 22916 4567 22928 4576
rect 20714 4496 20720 4548
rect 20772 4496 20778 4548
rect 22664 4480 22692 4567
rect 22922 4564 22928 4567
rect 22980 4564 22986 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24688 4604 24716 4644
rect 26418 4632 26424 4684
rect 26476 4632 26482 4684
rect 24837 4607 24895 4613
rect 24837 4604 24849 4607
rect 24688 4576 24849 4604
rect 24581 4567 24639 4573
rect 24837 4573 24849 4576
rect 24883 4573 24895 4607
rect 24837 4567 24895 4573
rect 22186 4468 22192 4480
rect 20456 4440 22192 4468
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 24596 4468 24624 4567
rect 26510 4564 26516 4616
rect 26568 4604 26574 4616
rect 26677 4607 26735 4613
rect 26677 4604 26689 4607
rect 26568 4576 26689 4604
rect 26568 4564 26574 4576
rect 26677 4573 26689 4576
rect 26723 4573 26735 4607
rect 26677 4567 26735 4573
rect 22704 4440 24624 4468
rect 22704 4428 22710 4440
rect 25590 4428 25596 4480
rect 25648 4468 25654 4480
rect 25774 4468 25780 4480
rect 25648 4440 25780 4468
rect 25648 4428 25654 4440
rect 25774 4428 25780 4440
rect 25832 4428 25838 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8294 4264 8300 4276
rect 8159 4236 8300 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 15933 4267 15991 4273
rect 15933 4264 15945 4267
rect 15896 4236 15945 4264
rect 15896 4224 15902 4236
rect 15933 4233 15945 4236
rect 15979 4233 15991 4267
rect 15933 4227 15991 4233
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 19886 4264 19892 4276
rect 17000 4236 19892 4264
rect 17000 4224 17006 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 27154 4264 27160 4276
rect 21416 4236 27160 4264
rect 21416 4224 21422 4236
rect 6932 4168 7144 4196
rect 1578 4088 1584 4140
rect 1636 4128 1642 4140
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1636 4100 1685 4128
rect 1636 4088 1642 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 1940 4131 1998 4137
rect 1940 4097 1952 4131
rect 1986 4128 1998 4131
rect 1986 4100 2774 4128
rect 1986 4097 1998 4100
rect 1940 4091 1998 4097
rect 2746 3924 2774 4100
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 4056 4131 4114 4137
rect 4056 4097 4068 4131
rect 4102 4128 4114 4131
rect 6932 4128 6960 4168
rect 7006 4137 7012 4140
rect 4102 4100 6960 4128
rect 4102 4097 4114 4100
rect 4056 4091 4114 4097
rect 7000 4091 7012 4137
rect 7006 4088 7012 4091
rect 7064 4088 7070 4140
rect 7116 4128 7144 4168
rect 8570 4156 8576 4208
rect 8628 4156 8634 4208
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 10505 4199 10563 4205
rect 10505 4196 10517 4199
rect 10468 4168 10517 4196
rect 10468 4156 10474 4168
rect 10505 4165 10517 4168
rect 10551 4165 10563 4199
rect 10505 4159 10563 4165
rect 13722 4156 13728 4208
rect 13780 4156 13786 4208
rect 13906 4156 13912 4208
rect 13964 4205 13970 4208
rect 13964 4199 13983 4205
rect 13971 4165 13983 4199
rect 13964 4159 13983 4165
rect 13964 4156 13970 4159
rect 14642 4156 14648 4208
rect 14700 4196 14706 4208
rect 14798 4199 14856 4205
rect 14798 4196 14810 4199
rect 14700 4168 14810 4196
rect 14700 4156 14706 4168
rect 14798 4165 14810 4168
rect 14844 4165 14856 4199
rect 14798 4159 14856 4165
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 17126 4205 17132 4208
rect 17098 4199 17132 4205
rect 17098 4196 17110 4199
rect 15712 4168 17110 4196
rect 15712 4156 15718 4168
rect 17098 4165 17110 4168
rect 17098 4159 17132 4165
rect 17126 4156 17132 4159
rect 17184 4156 17190 4208
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 20530 4196 20536 4208
rect 19392 4168 20536 4196
rect 19392 4156 19398 4168
rect 20530 4156 20536 4168
rect 20588 4156 20594 4208
rect 22112 4205 22140 4236
rect 27154 4224 27160 4236
rect 27212 4224 27218 4276
rect 22097 4199 22155 4205
rect 22097 4165 22109 4199
rect 22143 4165 22155 4199
rect 22097 4159 22155 4165
rect 22278 4156 22284 4208
rect 22336 4196 22342 4208
rect 22646 4196 22652 4208
rect 22336 4168 22652 4196
rect 22336 4156 22342 4168
rect 22646 4156 22652 4168
rect 22704 4156 22710 4208
rect 8588 4128 8616 4156
rect 7116 4100 8616 4128
rect 8840 4131 8898 4137
rect 8840 4097 8852 4131
rect 8886 4128 8898 4131
rect 10689 4131 10747 4137
rect 8886 4100 10364 4128
rect 8886 4097 8898 4100
rect 8840 4091 8898 4097
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 5500 4032 6745 4060
rect 5500 4020 5506 4032
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 6733 4023 6791 4029
rect 7760 4032 8585 4060
rect 3050 3952 3056 4004
rect 3108 3952 3114 4004
rect 6638 3924 6644 3936
rect 2746 3896 6644 3924
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6748 3924 6776 4023
rect 7098 3924 7104 3936
rect 6748 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3924 7162 3936
rect 7760 3924 7788 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 10336 4060 10364 4100
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 10870 4128 10876 4140
rect 10735 4100 10876 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 10870 4088 10876 4100
rect 10928 4128 10934 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 10928 4100 11897 4128
rect 10928 4088 10934 4100
rect 11885 4097 11897 4100
rect 11931 4128 11943 4131
rect 11974 4128 11980 4140
rect 11931 4100 11980 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12152 4131 12210 4137
rect 12152 4097 12164 4131
rect 12198 4128 12210 4131
rect 16758 4128 16764 4140
rect 12198 4100 16764 4128
rect 12198 4097 12210 4100
rect 12152 4091 12210 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19352 4128 19380 4156
rect 19199 4100 19380 4128
rect 19420 4131 19478 4137
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19420 4097 19432 4131
rect 19466 4128 19478 4131
rect 19702 4128 19708 4140
rect 19466 4100 19708 4128
rect 19466 4097 19478 4100
rect 19420 4091 19478 4097
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 25492 4131 25550 4137
rect 25492 4097 25504 4131
rect 25538 4128 25550 4131
rect 25774 4128 25780 4140
rect 25538 4100 25780 4128
rect 25538 4097 25550 4100
rect 25492 4091 25550 4097
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 25866 4088 25872 4140
rect 25924 4128 25930 4140
rect 25924 4100 26648 4128
rect 25924 4088 25930 4100
rect 10962 4060 10968 4072
rect 10336 4032 10968 4060
rect 8573 4023 8631 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 13320 4032 14565 4060
rect 13320 4020 13326 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 16850 4060 16856 4072
rect 15620 4032 16856 4060
rect 15620 4020 15626 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9640 3964 9965 3992
rect 9640 3952 9646 3964
rect 9953 3961 9965 3964
rect 9999 3992 10011 3995
rect 11790 3992 11796 4004
rect 9999 3964 11796 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 7156 3896 7788 3924
rect 7156 3884 7162 3896
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12250 3924 12256 3936
rect 11756 3896 12256 3924
rect 11756 3884 11762 3896
rect 12250 3884 12256 3896
rect 12308 3924 12314 3936
rect 13265 3927 13323 3933
rect 13265 3924 13277 3927
rect 12308 3896 13277 3924
rect 12308 3884 12314 3896
rect 13265 3893 13277 3896
rect 13311 3893 13323 3927
rect 13265 3887 13323 3893
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 13780 3896 13921 3924
rect 13780 3884 13786 3896
rect 13909 3893 13921 3896
rect 13955 3893 13967 3927
rect 13909 3887 13967 3893
rect 14090 3884 14096 3936
rect 14148 3884 14154 3936
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 19518 3924 19524 3936
rect 18279 3896 19524 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20530 3884 20536 3936
rect 20588 3884 20594 3936
rect 25240 3924 25268 4023
rect 26620 4001 26648 4100
rect 26605 3995 26663 4001
rect 26605 3961 26617 3995
rect 26651 3961 26663 3995
rect 26605 3955 26663 3961
rect 26418 3924 26424 3936
rect 25240 3896 26424 3924
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 4154 3680 4160 3732
rect 4212 3680 4218 3732
rect 6822 3680 6828 3732
rect 6880 3680 6886 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 13078 3720 13084 3732
rect 8628 3692 13084 3720
rect 8628 3680 8634 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 15378 3720 15384 3732
rect 13311 3692 15384 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 20530 3720 20536 3732
rect 17184 3692 20536 3720
rect 17184 3680 17190 3692
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23072 3692 23765 3720
rect 23072 3680 23078 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 28353 3723 28411 3729
rect 28353 3720 28365 3723
rect 25096 3692 28365 3720
rect 25096 3680 25102 3692
rect 28353 3689 28365 3692
rect 28399 3689 28411 3723
rect 28353 3683 28411 3689
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 5258 3652 5264 3664
rect 3375 3624 5264 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 10502 3652 10508 3664
rect 7064 3624 10508 3652
rect 7064 3612 7070 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 14458 3652 14464 3664
rect 12124 3624 14464 3652
rect 12124 3612 12130 3624
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 1949 3587 2007 3593
rect 1949 3584 1961 3587
rect 1636 3556 1961 3584
rect 1636 3544 1642 3556
rect 1949 3553 1961 3556
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 5442 3584 5448 3596
rect 3844 3556 5448 3584
rect 3844 3544 3850 3556
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 10686 3584 10692 3596
rect 6696 3556 10692 3584
rect 6696 3544 6702 3556
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10870 3544 10876 3596
rect 10928 3544 10934 3596
rect 13998 3584 14004 3596
rect 11932 3556 14004 3584
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 5718 3525 5724 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 1360 3488 4077 3516
rect 1360 3476 1366 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 5712 3516 5724 3525
rect 5679 3488 5724 3516
rect 4065 3479 4123 3485
rect 5712 3479 5724 3488
rect 5718 3476 5724 3479
rect 5776 3476 5782 3528
rect 11140 3519 11198 3525
rect 11140 3485 11152 3519
rect 11186 3516 11198 3519
rect 11932 3516 11960 3556
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 20533 3587 20591 3593
rect 20533 3584 20545 3587
rect 19300 3556 20545 3584
rect 19300 3544 19306 3556
rect 20533 3553 20545 3556
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 22278 3544 22284 3596
rect 22336 3584 22342 3596
rect 22373 3587 22431 3593
rect 22373 3584 22385 3587
rect 22336 3556 22385 3584
rect 22336 3544 22342 3556
rect 22373 3553 22385 3556
rect 22419 3553 22431 3587
rect 22373 3547 22431 3553
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 26970 3584 26976 3596
rect 26476 3556 26976 3584
rect 26476 3544 26482 3556
rect 26970 3544 26976 3556
rect 27028 3544 27034 3596
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 11186 3488 11960 3516
rect 11992 3488 12725 3516
rect 11186 3485 11198 3488
rect 11140 3479 11198 3485
rect 1394 3408 1400 3460
rect 1452 3448 1458 3460
rect 2194 3451 2252 3457
rect 2194 3448 2206 3451
rect 1452 3420 2206 3448
rect 1452 3408 1458 3420
rect 2194 3417 2206 3420
rect 2240 3417 2252 3451
rect 2194 3411 2252 3417
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 11992 3448 12020 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12713 3479 12771 3485
rect 12820 3488 13001 3516
rect 12820 3448 12848 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13170 3516 13176 3528
rect 13127 3488 13176 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 14734 3476 14740 3528
rect 14792 3476 14798 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 16908 3488 17417 3516
rect 16908 3476 16914 3488
rect 17405 3485 17417 3488
rect 17451 3516 17463 3519
rect 19334 3516 19340 3528
rect 17451 3488 19340 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 20806 3525 20812 3528
rect 20800 3516 20812 3525
rect 20767 3488 20812 3516
rect 20800 3479 20812 3488
rect 20806 3476 20812 3479
rect 20864 3476 20870 3528
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22646 3525 22652 3528
rect 22629 3519 22652 3525
rect 22629 3516 22641 3519
rect 22520 3488 22641 3516
rect 22520 3476 22526 3488
rect 22629 3485 22641 3488
rect 22629 3479 22652 3485
rect 22646 3476 22652 3479
rect 22704 3476 22710 3528
rect 25133 3519 25191 3525
rect 25133 3485 25145 3519
rect 25179 3516 25191 3519
rect 26436 3516 26464 3544
rect 25179 3488 26464 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 26878 3476 26884 3528
rect 26936 3516 26942 3528
rect 27229 3519 27287 3525
rect 27229 3516 27241 3519
rect 26936 3488 27241 3516
rect 26936 3476 26942 3488
rect 27229 3485 27241 3488
rect 27275 3485 27287 3519
rect 27229 3479 27287 3485
rect 9364 3420 12020 3448
rect 12084 3420 12848 3448
rect 9364 3408 9370 3420
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 12084 3380 12112 3420
rect 12894 3408 12900 3460
rect 12952 3408 12958 3460
rect 13354 3448 13360 3460
rect 13004 3420 13360 3448
rect 6236 3352 12112 3380
rect 12253 3383 12311 3389
rect 6236 3340 6242 3352
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12618 3380 12624 3392
rect 12299 3352 12624 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12618 3340 12624 3352
rect 12676 3380 12682 3392
rect 13004 3380 13032 3420
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 15004 3451 15062 3457
rect 15004 3417 15016 3451
rect 15050 3448 15062 3451
rect 16206 3448 16212 3460
rect 15050 3420 16212 3448
rect 15050 3417 15062 3420
rect 15004 3411 15062 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 17672 3451 17730 3457
rect 17672 3417 17684 3451
rect 17718 3448 17730 3451
rect 20898 3448 20904 3460
rect 17718 3420 20904 3448
rect 17718 3417 17730 3420
rect 17672 3411 17730 3417
rect 20898 3408 20904 3420
rect 20956 3448 20962 3460
rect 25400 3451 25458 3457
rect 20956 3420 21956 3448
rect 20956 3408 20962 3420
rect 12676 3352 13032 3380
rect 12676 3340 12682 3352
rect 15194 3340 15200 3392
rect 15252 3380 15258 3392
rect 16022 3380 16028 3392
rect 15252 3352 16028 3380
rect 15252 3340 15258 3352
rect 16022 3340 16028 3352
rect 16080 3380 16086 3392
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 16080 3352 16129 3380
rect 16080 3340 16086 3352
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16117 3343 16175 3349
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 21928 3389 21956 3420
rect 25400 3417 25412 3451
rect 25446 3448 25458 3451
rect 25590 3448 25596 3460
rect 25446 3420 25596 3448
rect 25446 3417 25458 3420
rect 25400 3411 25458 3417
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 16356 3352 18797 3380
rect 16356 3340 16362 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 21913 3383 21971 3389
rect 21913 3349 21925 3383
rect 21959 3349 21971 3383
rect 21913 3343 21971 3349
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 26513 3383 26571 3389
rect 26513 3380 26525 3383
rect 24268 3352 26525 3380
rect 24268 3340 24274 3352
rect 26513 3349 26525 3352
rect 26559 3349 26571 3383
rect 26513 3343 26571 3349
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 3602 3136 3608 3188
rect 3660 3136 3666 3188
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11149 3179 11207 3185
rect 11149 3176 11161 3179
rect 11112 3148 11161 3176
rect 11112 3136 11118 3148
rect 11149 3145 11161 3148
rect 11195 3145 11207 3179
rect 11149 3139 11207 3145
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 13722 3176 13728 3188
rect 12676 3148 13728 3176
rect 12676 3136 12682 3148
rect 13722 3136 13728 3148
rect 13780 3176 13786 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13780 3148 13829 3176
rect 13780 3136 13786 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 14826 3136 14832 3188
rect 14884 3176 14890 3188
rect 15286 3176 15292 3188
rect 14884 3148 15292 3176
rect 14884 3136 14890 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 16482 3136 16488 3188
rect 16540 3176 16546 3188
rect 16540 3148 18184 3176
rect 16540 3136 16546 3148
rect 10036 3111 10094 3117
rect 10036 3077 10048 3111
rect 10082 3108 10094 3111
rect 11698 3108 11704 3120
rect 10082 3080 11704 3108
rect 10082 3077 10094 3080
rect 10036 3071 10094 3077
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 12704 3111 12762 3117
rect 12704 3077 12716 3111
rect 12750 3108 12762 3111
rect 15194 3108 15200 3120
rect 12750 3080 15200 3108
rect 12750 3077 12762 3080
rect 12704 3071 12762 3077
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 17120 3111 17178 3117
rect 17120 3077 17132 3111
rect 17166 3108 17178 3111
rect 17678 3108 17684 3120
rect 17166 3080 17684 3108
rect 17166 3077 17178 3080
rect 17120 3071 17178 3077
rect 17678 3068 17684 3080
rect 17736 3108 17742 3120
rect 17862 3108 17868 3120
rect 17736 3080 17868 3108
rect 17736 3068 17742 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 18156 3108 18184 3148
rect 18230 3136 18236 3188
rect 18288 3136 18294 3188
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 20901 3179 20959 3185
rect 20901 3176 20913 3179
rect 20772 3148 20913 3176
rect 20772 3136 20778 3148
rect 20901 3145 20913 3148
rect 20947 3145 20959 3179
rect 20901 3139 20959 3145
rect 22922 3136 22928 3188
rect 22980 3176 22986 3188
rect 23477 3179 23535 3185
rect 23477 3176 23489 3179
rect 22980 3148 23489 3176
rect 22980 3136 22986 3148
rect 23477 3145 23489 3148
rect 23523 3145 23535 3179
rect 23477 3139 23535 3145
rect 18874 3108 18880 3120
rect 18156 3080 18880 3108
rect 18874 3068 18880 3080
rect 18932 3068 18938 3120
rect 19518 3068 19524 3120
rect 19576 3108 19582 3120
rect 19766 3111 19824 3117
rect 19766 3108 19778 3111
rect 19576 3080 19778 3108
rect 19576 3068 19582 3080
rect 19766 3077 19778 3080
rect 19812 3077 19824 3111
rect 22278 3108 22284 3120
rect 19766 3071 19824 3077
rect 22112 3080 22284 3108
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1946 3040 1952 3052
rect 1636 3012 1952 3040
rect 1636 3000 1642 3012
rect 1946 3000 1952 3012
rect 2004 3040 2010 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 2004 3012 2237 3040
rect 2004 3000 2010 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4154 3040 4160 3052
rect 3844 3012 4160 3040
rect 3844 3000 3850 3012
rect 4154 3000 4160 3012
rect 4212 3040 4218 3052
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 4212 3012 4353 3040
rect 4212 3000 4218 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4608 3043 4666 3049
rect 4608 3009 4620 3043
rect 4654 3040 4666 3043
rect 9306 3040 9312 3052
rect 4654 3012 9312 3040
rect 4654 3009 4666 3012
rect 4608 3003 4666 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 9858 3040 9864 3052
rect 9815 3012 9864 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 9858 3000 9864 3012
rect 9916 3040 9922 3052
rect 10870 3040 10876 3052
rect 9916 3012 10876 3040
rect 9916 3000 9922 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12032 3012 12449 3040
rect 12032 3000 12038 3012
rect 12437 3009 12449 3012
rect 12483 3040 12495 3043
rect 12483 3012 13584 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 13556 2972 13584 3012
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14608 3012 14657 3040
rect 14608 3000 14614 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 14734 2972 14740 2984
rect 13556 2944 14740 2972
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 14936 2904 14964 3003
rect 15010 3000 15016 3052
rect 15068 3000 15074 3052
rect 15746 3000 15752 3052
rect 15804 3000 15810 3052
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16850 3040 16856 3052
rect 15979 3012 16856 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15948 2972 15976 3003
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 20898 3040 20904 3052
rect 20772 3012 20904 3040
rect 20772 3000 20778 3012
rect 20898 3000 20904 3012
rect 20956 3000 20962 3052
rect 22112 3049 22140 3080
rect 22278 3068 22284 3080
rect 22336 3108 22342 3120
rect 22336 3080 23980 3108
rect 22336 3068 22342 3080
rect 23952 3052 23980 3080
rect 24026 3068 24032 3120
rect 24084 3108 24090 3120
rect 24210 3117 24216 3120
rect 24204 3108 24216 3117
rect 24084 3080 24216 3108
rect 24084 3068 24090 3080
rect 24204 3071 24216 3080
rect 24210 3068 24216 3071
rect 24268 3068 24274 3120
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3009 22155 3043
rect 22097 3003 22155 3009
rect 22186 3000 22192 3052
rect 22244 3040 22250 3052
rect 22364 3043 22422 3049
rect 22364 3040 22376 3043
rect 22244 3012 22376 3040
rect 22244 3000 22250 3012
rect 22364 3009 22376 3012
rect 22410 3040 22422 3043
rect 23290 3040 23296 3052
rect 22410 3012 23296 3040
rect 22410 3009 22422 3012
rect 22364 3003 22422 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23934 3000 23940 3052
rect 23992 3000 23998 3052
rect 15712 2944 15976 2972
rect 15712 2932 15718 2944
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19392 2944 19533 2972
rect 19392 2932 19398 2944
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 11112 2876 12434 2904
rect 11112 2864 11118 2876
rect 5718 2796 5724 2848
rect 5776 2796 5782 2848
rect 12406 2836 12434 2876
rect 13372 2876 14964 2904
rect 15197 2907 15255 2913
rect 13372 2836 13400 2876
rect 15197 2873 15209 2907
rect 15243 2904 15255 2907
rect 15243 2876 16896 2904
rect 15243 2873 15255 2876
rect 15197 2867 15255 2873
rect 12406 2808 13400 2836
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 16390 2836 16396 2848
rect 15804 2808 16396 2836
rect 15804 2796 15810 2808
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 16868 2836 16896 2876
rect 18138 2836 18144 2848
rect 16868 2808 18144 2836
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 24912 2808 25329 2836
rect 24912 2796 24918 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 1670 2592 1676 2644
rect 1728 2592 1734 2644
rect 3326 2592 3332 2644
rect 3384 2592 3390 2644
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 5810 2632 5816 2644
rect 5399 2604 5816 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 9398 2632 9404 2644
rect 7331 2604 9404 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 12066 2632 12072 2644
rect 11287 2604 12072 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 12802 2632 12808 2644
rect 12308 2604 12808 2632
rect 12308 2592 12314 2604
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2632 13691 2635
rect 13814 2632 13820 2644
rect 13679 2604 13820 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 17954 2592 17960 2644
rect 18012 2592 18018 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 18196 2604 18429 2632
rect 18196 2592 18202 2604
rect 18417 2601 18429 2604
rect 18463 2601 18475 2635
rect 18417 2595 18475 2601
rect 18874 2592 18880 2644
rect 18932 2592 18938 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19024 2604 22416 2632
rect 19024 2592 19030 2604
rect 12529 2567 12587 2573
rect 12529 2533 12541 2567
rect 12575 2533 12587 2567
rect 12529 2527 12587 2533
rect 1946 2456 1952 2508
rect 2004 2456 2010 2508
rect 9858 2456 9864 2508
rect 9916 2456 9922 2508
rect 12250 2456 12256 2508
rect 12308 2456 12314 2508
rect 1964 2428 1992 2456
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 1964 2400 3985 2428
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5902 2428 5908 2440
rect 5500 2400 5908 2428
rect 5500 2388 5506 2400
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6178 2437 6184 2440
rect 6172 2391 6184 2437
rect 6178 2388 6184 2391
rect 6236 2388 6242 2440
rect 10128 2431 10186 2437
rect 10128 2397 10140 2431
rect 10174 2428 10186 2431
rect 10870 2428 10876 2440
rect 10174 2400 10876 2428
rect 10174 2397 10186 2400
rect 10128 2391 10186 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11112 2400 11989 2428
rect 11112 2388 11118 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2428 12219 2431
rect 12268 2428 12296 2456
rect 12207 2400 12296 2428
rect 12345 2431 12403 2437
rect 12207 2397 12219 2400
rect 12161 2391 12219 2397
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12544 2428 12572 2527
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16264 2536 17908 2564
rect 16264 2524 16270 2536
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14792 2468 14841 2496
rect 14792 2456 14798 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17092 2468 17821 2496
rect 17092 2456 17098 2468
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12544 2400 13001 2428
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13078 2388 13084 2440
rect 13136 2388 13142 2440
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13228 2400 13277 2428
rect 13228 2388 13234 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 13495 2431 13553 2437
rect 13495 2397 13507 2431
rect 13541 2428 13553 2431
rect 14642 2428 14648 2440
rect 13541 2400 14648 2428
rect 13541 2397 13553 2400
rect 13495 2391 13553 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 17310 2388 17316 2440
rect 17368 2388 17374 2440
rect 17461 2431 17519 2437
rect 17461 2397 17473 2431
rect 17507 2428 17519 2431
rect 17589 2431 17647 2437
rect 17507 2397 17540 2428
rect 17461 2391 17540 2397
rect 17589 2397 17601 2431
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 1670 2320 1676 2372
rect 1728 2360 1734 2372
rect 2194 2363 2252 2369
rect 2194 2360 2206 2363
rect 1728 2332 2206 2360
rect 1728 2320 1734 2332
rect 2194 2329 2206 2332
rect 2240 2329 2252 2363
rect 2194 2323 2252 2329
rect 4240 2363 4298 2369
rect 4240 2329 4252 2363
rect 4286 2360 4298 2363
rect 5813 2363 5871 2369
rect 5813 2360 5825 2363
rect 4286 2332 5825 2360
rect 4286 2329 4298 2332
rect 4240 2323 4298 2329
rect 5813 2329 5825 2332
rect 5859 2360 5871 2363
rect 6454 2360 6460 2372
rect 5859 2332 6460 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 6454 2320 6460 2332
rect 6512 2320 6518 2372
rect 12253 2363 12311 2369
rect 12253 2329 12265 2363
rect 12299 2360 12311 2363
rect 15096 2363 15154 2369
rect 15096 2360 15108 2363
rect 12299 2332 15108 2360
rect 12299 2329 12311 2332
rect 12253 2323 12311 2329
rect 15096 2329 15108 2332
rect 15142 2360 15154 2363
rect 15286 2360 15292 2372
rect 15142 2332 15292 2360
rect 15142 2329 15154 2332
rect 15096 2323 15154 2329
rect 15286 2320 15292 2332
rect 15344 2320 15350 2372
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 17310 2292 17316 2304
rect 13136 2264 17316 2292
rect 13136 2252 13142 2264
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17512 2292 17540 2391
rect 17604 2360 17632 2391
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 17793 2437 17821 2468
rect 17778 2431 17836 2437
rect 17778 2397 17790 2431
rect 17824 2397 17836 2431
rect 17778 2391 17836 2397
rect 17604 2332 17816 2360
rect 17788 2304 17816 2332
rect 17678 2292 17684 2304
rect 17512 2264 17684 2292
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 17770 2252 17776 2304
rect 17828 2252 17834 2304
rect 17880 2292 17908 2536
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 20622 2564 20628 2576
rect 18380 2536 20628 2564
rect 18380 2524 18386 2536
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18509 2499 18567 2505
rect 18509 2496 18521 2499
rect 18104 2468 18521 2496
rect 18104 2456 18110 2468
rect 18509 2465 18521 2468
rect 18555 2465 18567 2499
rect 18509 2459 18567 2465
rect 18782 2456 18788 2508
rect 18840 2496 18846 2508
rect 18840 2468 21128 2496
rect 18840 2456 18846 2468
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 19150 2428 19156 2440
rect 18739 2400 19156 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 18417 2363 18475 2369
rect 18417 2329 18429 2363
rect 18463 2360 18475 2363
rect 19242 2360 19248 2372
rect 18463 2332 19248 2360
rect 18463 2329 18475 2332
rect 18417 2323 18475 2329
rect 19242 2320 19248 2332
rect 19300 2320 19306 2372
rect 20990 2292 20996 2304
rect 17880 2264 20996 2292
rect 20990 2252 20996 2264
rect 21048 2252 21054 2304
rect 21100 2292 21128 2468
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22278 2428 22284 2440
rect 21315 2400 22284 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 22388 2428 22416 2604
rect 24118 2592 24124 2644
rect 24176 2632 24182 2644
rect 28353 2635 28411 2641
rect 28353 2632 28365 2635
rect 24176 2604 28365 2632
rect 24176 2592 24182 2604
rect 28353 2601 28365 2604
rect 28399 2601 28411 2635
rect 28353 2595 28411 2601
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23992 2468 24593 2496
rect 23992 2456 23998 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 26970 2456 26976 2508
rect 27028 2456 27034 2508
rect 25682 2428 25688 2440
rect 22388 2400 25688 2428
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 25958 2388 25964 2440
rect 26016 2428 26022 2440
rect 27229 2431 27287 2437
rect 27229 2428 27241 2431
rect 26016 2400 27241 2428
rect 26016 2388 26022 2400
rect 27229 2397 27241 2400
rect 27275 2397 27287 2431
rect 27229 2391 27287 2397
rect 21536 2363 21594 2369
rect 21536 2329 21548 2363
rect 21582 2360 21594 2363
rect 22370 2360 22376 2372
rect 21582 2332 22376 2360
rect 21582 2329 21594 2332
rect 21536 2323 21594 2329
rect 22370 2320 22376 2332
rect 22428 2360 22434 2372
rect 24854 2369 24860 2372
rect 24848 2360 24860 2369
rect 22428 2332 23244 2360
rect 24815 2332 24860 2360
rect 22428 2320 22434 2332
rect 22649 2295 22707 2301
rect 22649 2292 22661 2295
rect 21100 2264 22661 2292
rect 22649 2261 22661 2264
rect 22695 2261 22707 2295
rect 23216 2292 23244 2332
rect 24848 2323 24860 2332
rect 24854 2320 24860 2323
rect 24912 2320 24918 2372
rect 25961 2295 26019 2301
rect 25961 2292 25973 2295
rect 23216 2264 25973 2292
rect 22649 2255 22707 2261
rect 25961 2261 25973 2264
rect 26007 2261 26019 2295
rect 25961 2255 26019 2261
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 2317 2091 2375 2097
rect 2317 2057 2329 2091
rect 2363 2088 2375 2091
rect 5537 2091 5595 2097
rect 2363 2060 5488 2088
rect 2363 2057 2375 2060
rect 2317 2051 2375 2057
rect 1946 1912 1952 1964
rect 2004 1952 2010 1964
rect 3697 1955 3755 1961
rect 3697 1952 3709 1955
rect 2004 1924 3709 1952
rect 2004 1912 2010 1924
rect 3697 1921 3709 1924
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 4154 1912 4160 1964
rect 4212 1912 4218 1964
rect 4424 1955 4482 1961
rect 4424 1921 4436 1955
rect 4470 1952 4482 1955
rect 5460 1952 5488 2060
rect 5537 2057 5549 2091
rect 5583 2088 5595 2091
rect 7374 2088 7380 2100
rect 5583 2060 7380 2088
rect 5583 2057 5595 2060
rect 5537 2051 5595 2057
rect 7374 2048 7380 2060
rect 7432 2048 7438 2100
rect 9306 2048 9312 2100
rect 9364 2048 9370 2100
rect 13630 2088 13636 2100
rect 11716 2060 13636 2088
rect 8196 2023 8254 2029
rect 8196 1989 8208 2023
rect 8242 2020 8254 2023
rect 9582 2020 9588 2032
rect 8242 1992 9588 2020
rect 8242 1989 8254 1992
rect 8196 1983 8254 1989
rect 9582 1980 9588 1992
rect 9640 1980 9646 2032
rect 11238 2020 11244 2032
rect 9692 1992 11244 2020
rect 9692 1952 9720 1992
rect 11238 1980 11244 1992
rect 11296 1980 11302 2032
rect 11716 2029 11744 2060
rect 13630 2048 13636 2060
rect 13688 2048 13694 2100
rect 13909 2091 13967 2097
rect 13909 2057 13921 2091
rect 13955 2088 13967 2091
rect 13998 2088 14004 2100
rect 13955 2060 14004 2088
rect 13955 2057 13967 2060
rect 13909 2051 13967 2057
rect 13998 2048 14004 2060
rect 14056 2048 14062 2100
rect 15286 2048 15292 2100
rect 15344 2088 15350 2100
rect 18325 2091 18383 2097
rect 18325 2088 18337 2091
rect 15344 2060 18337 2088
rect 15344 2048 15350 2060
rect 18325 2057 18337 2060
rect 18371 2057 18383 2091
rect 18325 2051 18383 2057
rect 20165 2091 20223 2097
rect 20165 2057 20177 2091
rect 20211 2057 20223 2091
rect 20165 2051 20223 2057
rect 11701 2023 11759 2029
rect 11701 1989 11713 2023
rect 11747 1989 11759 2023
rect 11701 1983 11759 1989
rect 11917 2023 11975 2029
rect 11917 1989 11929 2023
rect 11963 2020 11975 2023
rect 12158 2020 12164 2032
rect 11963 1992 12164 2020
rect 11963 1989 11975 1992
rect 11917 1983 11975 1989
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 12618 2020 12624 2032
rect 12406 1992 12624 2020
rect 4470 1924 5396 1952
rect 5460 1924 9720 1952
rect 9769 1955 9827 1961
rect 4470 1921 4482 1924
rect 4424 1915 4482 1921
rect 1765 1887 1823 1893
rect 1765 1853 1777 1887
rect 1811 1884 1823 1887
rect 3418 1884 3424 1896
rect 1811 1856 3424 1884
rect 1811 1853 1823 1856
rect 1765 1847 1823 1853
rect 3418 1844 3424 1856
rect 3476 1844 3482 1896
rect 5368 1884 5396 1924
rect 9769 1921 9781 1955
rect 9815 1952 9827 1955
rect 9858 1952 9864 1964
rect 9815 1924 9864 1952
rect 9815 1921 9827 1924
rect 9769 1915 9827 1921
rect 9858 1912 9864 1924
rect 9916 1912 9922 1964
rect 10036 1955 10094 1961
rect 10036 1921 10048 1955
rect 10082 1952 10094 1955
rect 12406 1952 12434 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 12796 2023 12854 2029
rect 12796 2020 12808 2023
rect 12719 1992 12808 2020
rect 10082 1924 12434 1952
rect 10082 1921 10094 1924
rect 10036 1915 10094 1921
rect 12526 1912 12532 1964
rect 12584 1912 12590 1964
rect 12719 1952 12747 1992
rect 12796 1989 12808 1992
rect 12842 2020 12854 2023
rect 13446 2020 13452 2032
rect 12842 1992 13452 2020
rect 12842 1989 12854 1992
rect 12796 1983 12854 1989
rect 13446 1980 13452 1992
rect 13504 1980 13510 2032
rect 15188 2023 15246 2029
rect 15188 1989 15200 2023
rect 15234 2020 15246 2023
rect 15746 2020 15752 2032
rect 15234 1992 15752 2020
rect 15234 1989 15246 1992
rect 15188 1983 15246 1989
rect 15746 1980 15752 1992
rect 15804 2020 15810 2032
rect 16298 2020 16304 2032
rect 15804 1992 16304 2020
rect 15804 1980 15810 1992
rect 16298 1980 16304 1992
rect 16356 1980 16362 2032
rect 17212 2023 17270 2029
rect 17212 1989 17224 2023
rect 17258 2020 17270 2023
rect 17494 2020 17500 2032
rect 17258 1992 17500 2020
rect 17258 1989 17270 1992
rect 17212 1983 17270 1989
rect 17494 1980 17500 1992
rect 17552 1980 17558 2032
rect 17678 1980 17684 2032
rect 17736 2020 17742 2032
rect 19702 2020 19708 2032
rect 17736 1992 19708 2020
rect 17736 1980 17742 1992
rect 19702 1980 19708 1992
rect 19760 1980 19766 2032
rect 20180 2020 20208 2051
rect 21266 2048 21272 2100
rect 21324 2048 21330 2100
rect 22278 2048 22284 2100
rect 22336 2048 22342 2100
rect 23290 2048 23296 2100
rect 23348 2088 23354 2100
rect 23385 2091 23443 2097
rect 23385 2088 23397 2091
rect 23348 2060 23397 2088
rect 23348 2048 23354 2060
rect 23385 2057 23397 2060
rect 23431 2057 23443 2091
rect 25225 2091 25283 2097
rect 25225 2088 25237 2091
rect 23385 2051 23443 2057
rect 23492 2060 25237 2088
rect 21634 2020 21640 2032
rect 20180 1992 21640 2020
rect 21634 1980 21640 1992
rect 21692 1980 21698 2032
rect 22296 2020 22324 2048
rect 22020 1992 22324 2020
rect 17034 1952 17040 1964
rect 12636 1924 12747 1952
rect 16868 1924 17040 1952
rect 5626 1884 5632 1896
rect 5368 1856 5632 1884
rect 5626 1844 5632 1856
rect 5684 1844 5690 1896
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 7929 1887 7987 1893
rect 7929 1884 7941 1887
rect 5960 1856 7941 1884
rect 5960 1844 5966 1856
rect 7929 1853 7941 1856
rect 7975 1853 7987 1887
rect 12636 1884 12664 1924
rect 7929 1847 7987 1853
rect 12406 1856 12664 1884
rect 14921 1887 14979 1893
rect 7944 1748 7972 1847
rect 11149 1819 11207 1825
rect 11149 1785 11161 1819
rect 11195 1816 11207 1819
rect 12406 1816 12434 1856
rect 14921 1853 14933 1887
rect 14967 1853 14979 1887
rect 14921 1847 14979 1853
rect 11195 1788 12434 1816
rect 11195 1785 11207 1788
rect 11149 1779 11207 1785
rect 8202 1748 8208 1760
rect 7944 1720 8208 1748
rect 8202 1708 8208 1720
rect 8260 1708 8266 1760
rect 11882 1708 11888 1760
rect 11940 1708 11946 1760
rect 12069 1751 12127 1757
rect 12069 1717 12081 1751
rect 12115 1748 12127 1751
rect 14550 1748 14556 1760
rect 12115 1720 14556 1748
rect 12115 1717 12127 1720
rect 12069 1711 12127 1717
rect 14550 1708 14556 1720
rect 14608 1708 14614 1760
rect 14936 1748 14964 1847
rect 16301 1819 16359 1825
rect 16301 1785 16313 1819
rect 16347 1816 16359 1819
rect 16868 1816 16896 1924
rect 17034 1912 17040 1924
rect 17092 1952 17098 1964
rect 19041 1955 19099 1961
rect 19041 1952 19053 1955
rect 17092 1924 19053 1952
rect 17092 1912 17098 1924
rect 19041 1921 19053 1924
rect 19087 1921 19099 1955
rect 19041 1915 19099 1921
rect 20625 1955 20683 1961
rect 20625 1921 20637 1955
rect 20671 1921 20683 1955
rect 20625 1915 20683 1921
rect 16945 1887 17003 1893
rect 16945 1853 16957 1887
rect 16991 1853 17003 1887
rect 16945 1847 17003 1853
rect 18785 1887 18843 1893
rect 18785 1853 18797 1887
rect 18831 1853 18843 1887
rect 18785 1847 18843 1853
rect 16347 1788 16896 1816
rect 16347 1785 16359 1788
rect 16301 1779 16359 1785
rect 15654 1748 15660 1760
rect 14936 1720 15660 1748
rect 15654 1708 15660 1720
rect 15712 1748 15718 1760
rect 16960 1748 16988 1847
rect 18800 1748 18828 1847
rect 15712 1720 18828 1748
rect 20640 1748 20668 1915
rect 20714 1912 20720 1964
rect 20772 1912 20778 1964
rect 20901 1955 20959 1961
rect 20901 1921 20913 1955
rect 20947 1921 20959 1955
rect 20901 1915 20959 1921
rect 20916 1884 20944 1915
rect 20990 1912 20996 1964
rect 21048 1912 21054 1964
rect 21082 1912 21088 1964
rect 21140 1961 21146 1964
rect 22020 1961 22048 1992
rect 22646 1980 22652 2032
rect 22704 2020 22710 2032
rect 23492 2020 23520 2060
rect 25225 2057 25237 2060
rect 25271 2057 25283 2091
rect 25225 2051 25283 2057
rect 22704 1992 23520 2020
rect 22704 1980 22710 1992
rect 23658 1980 23664 2032
rect 23716 2020 23722 2032
rect 24118 2029 24124 2032
rect 24090 2023 24124 2029
rect 24090 2020 24102 2023
rect 23716 1992 24102 2020
rect 23716 1980 23722 1992
rect 24090 1989 24102 1992
rect 24090 1983 24124 1989
rect 24118 1980 24124 1983
rect 24176 1980 24182 2032
rect 24210 1980 24216 2032
rect 24268 1980 24274 2032
rect 24854 1980 24860 2032
rect 24912 2020 24918 2032
rect 25961 2023 26019 2029
rect 25961 2020 25973 2023
rect 24912 1992 25973 2020
rect 24912 1980 24918 1992
rect 25961 1989 25973 1992
rect 26007 1989 26019 2023
rect 25961 1983 26019 1989
rect 21140 1952 21148 1961
rect 22005 1955 22063 1961
rect 21140 1924 21185 1952
rect 21140 1915 21148 1924
rect 22005 1921 22017 1955
rect 22051 1921 22063 1955
rect 22005 1915 22063 1921
rect 22272 1955 22330 1961
rect 22272 1921 22284 1955
rect 22318 1952 22330 1955
rect 23014 1952 23020 1964
rect 22318 1924 23020 1952
rect 22318 1921 22330 1924
rect 22272 1915 22330 1921
rect 21140 1912 21146 1915
rect 23014 1912 23020 1924
rect 23072 1912 23078 1964
rect 23845 1955 23903 1961
rect 23845 1921 23857 1955
rect 23891 1952 23903 1955
rect 23934 1952 23940 1964
rect 23891 1924 23940 1952
rect 23891 1921 23903 1924
rect 23845 1915 23903 1921
rect 23934 1912 23940 1924
rect 23992 1912 23998 1964
rect 24228 1952 24256 1980
rect 25685 1955 25743 1961
rect 24228 1924 24900 1952
rect 21450 1884 21456 1896
rect 20916 1856 21456 1884
rect 21450 1844 21456 1856
rect 21508 1844 21514 1896
rect 24872 1884 24900 1924
rect 25685 1921 25697 1955
rect 25731 1952 25743 1955
rect 25774 1952 25780 1964
rect 25731 1924 25780 1952
rect 25731 1921 25743 1924
rect 25685 1915 25743 1921
rect 25774 1912 25780 1924
rect 25832 1912 25838 1964
rect 25869 1955 25927 1961
rect 25869 1921 25881 1955
rect 25915 1921 25927 1955
rect 25869 1915 25927 1921
rect 26053 1955 26111 1961
rect 26053 1921 26065 1955
rect 26099 1921 26111 1955
rect 26053 1915 26111 1921
rect 25884 1884 25912 1915
rect 24872 1856 25912 1884
rect 25958 1844 25964 1896
rect 26016 1884 26022 1896
rect 26068 1884 26096 1915
rect 26016 1856 26096 1884
rect 26016 1844 26022 1856
rect 26237 1751 26295 1757
rect 26237 1748 26249 1751
rect 20640 1720 26249 1748
rect 15712 1708 15718 1720
rect 26237 1717 26249 1720
rect 26283 1717 26295 1751
rect 26237 1711 26295 1717
rect 1104 1658 28888 1680
rect 1104 1606 4423 1658
rect 4475 1606 4487 1658
rect 4539 1606 4551 1658
rect 4603 1606 4615 1658
rect 4667 1606 4679 1658
rect 4731 1606 11369 1658
rect 11421 1606 11433 1658
rect 11485 1606 11497 1658
rect 11549 1606 11561 1658
rect 11613 1606 11625 1658
rect 11677 1606 18315 1658
rect 18367 1606 18379 1658
rect 18431 1606 18443 1658
rect 18495 1606 18507 1658
rect 18559 1606 18571 1658
rect 18623 1606 25261 1658
rect 25313 1606 25325 1658
rect 25377 1606 25389 1658
rect 25441 1606 25453 1658
rect 25505 1606 25517 1658
rect 25569 1606 28888 1658
rect 1104 1584 28888 1606
rect 5626 1504 5632 1556
rect 5684 1544 5690 1556
rect 11882 1544 11888 1556
rect 5684 1516 11888 1544
rect 5684 1504 5690 1516
rect 11882 1504 11888 1516
rect 11940 1504 11946 1556
rect 14550 1504 14556 1556
rect 14608 1504 14614 1556
rect 14737 1547 14795 1553
rect 14737 1513 14749 1547
rect 14783 1544 14795 1547
rect 16666 1544 16672 1556
rect 14783 1516 16672 1544
rect 14783 1513 14795 1516
rect 14737 1507 14795 1513
rect 16666 1504 16672 1516
rect 16724 1504 16730 1556
rect 17770 1504 17776 1556
rect 17828 1544 17834 1556
rect 22554 1544 22560 1556
rect 17828 1516 19334 1544
rect 17828 1504 17834 1516
rect 14090 1436 14096 1488
rect 14148 1476 14154 1488
rect 14645 1479 14703 1485
rect 14645 1476 14657 1479
rect 14148 1448 14657 1476
rect 14148 1436 14154 1448
rect 14645 1445 14657 1448
rect 14691 1445 14703 1479
rect 14645 1439 14703 1445
rect 1946 1368 1952 1420
rect 2004 1368 2010 1420
rect 12989 1411 13047 1417
rect 12989 1377 13001 1411
rect 13035 1408 13047 1411
rect 13078 1408 13084 1420
rect 13035 1380 13084 1408
rect 13035 1377 13047 1380
rect 12989 1371 13047 1377
rect 13078 1368 13084 1380
rect 13136 1368 13142 1420
rect 14660 1380 14964 1408
rect 1964 1340 1992 1368
rect 3973 1343 4031 1349
rect 3973 1340 3985 1343
rect 1964 1312 3985 1340
rect 3973 1309 3985 1312
rect 4019 1309 4031 1343
rect 3973 1303 4031 1309
rect 8294 1300 8300 1352
rect 8352 1340 8358 1352
rect 9398 1349 9404 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 8352 1312 9137 1340
rect 8352 1300 8358 1312
rect 9125 1309 9137 1312
rect 9171 1309 9183 1343
rect 9392 1340 9404 1349
rect 9359 1312 9404 1340
rect 9125 1303 9183 1309
rect 9392 1303 9404 1312
rect 9398 1300 9404 1303
rect 9456 1300 9462 1352
rect 11974 1300 11980 1352
rect 12032 1300 12038 1352
rect 12161 1343 12219 1349
rect 12161 1309 12173 1343
rect 12207 1309 12219 1343
rect 12161 1303 12219 1309
rect 14369 1343 14427 1349
rect 14369 1309 14381 1343
rect 14415 1340 14427 1343
rect 14660 1340 14688 1380
rect 14415 1312 14688 1340
rect 14829 1343 14887 1349
rect 14415 1309 14427 1312
rect 14369 1303 14427 1309
rect 14829 1309 14841 1343
rect 14875 1309 14887 1343
rect 14936 1340 14964 1380
rect 15470 1340 15476 1352
rect 14936 1312 15476 1340
rect 14829 1303 14887 1309
rect 2222 1281 2228 1284
rect 1673 1275 1731 1281
rect 1673 1241 1685 1275
rect 1719 1272 1731 1275
rect 2216 1272 2228 1281
rect 1719 1244 2228 1272
rect 1719 1241 1731 1244
rect 1673 1235 1731 1241
rect 2216 1235 2228 1244
rect 2222 1232 2228 1235
rect 2280 1232 2286 1284
rect 4240 1275 4298 1281
rect 4240 1241 4252 1275
rect 4286 1272 4298 1275
rect 4286 1244 5764 1272
rect 4286 1241 4298 1244
rect 4240 1235 4298 1241
rect 3326 1164 3332 1216
rect 3384 1164 3390 1216
rect 5350 1164 5356 1216
rect 5408 1164 5414 1216
rect 5736 1213 5764 1244
rect 9490 1232 9496 1284
rect 9548 1272 9554 1284
rect 12176 1272 12204 1303
rect 9548 1244 12204 1272
rect 9548 1232 9554 1244
rect 12342 1232 12348 1284
rect 12400 1272 12406 1284
rect 14844 1272 14872 1303
rect 15470 1300 15476 1312
rect 15528 1300 15534 1352
rect 15746 1300 15752 1352
rect 15804 1300 15810 1352
rect 16022 1300 16028 1352
rect 16080 1300 16086 1352
rect 16114 1300 16120 1352
rect 16172 1300 16178 1352
rect 16390 1300 16396 1352
rect 16448 1340 16454 1352
rect 17497 1343 17555 1349
rect 17497 1340 17509 1343
rect 16448 1312 17509 1340
rect 16448 1300 16454 1312
rect 17497 1309 17509 1312
rect 17543 1309 17555 1343
rect 18046 1340 18052 1352
rect 17497 1303 17555 1309
rect 17604 1312 18052 1340
rect 12400 1244 14872 1272
rect 12400 1232 12406 1244
rect 15930 1232 15936 1284
rect 15988 1232 15994 1284
rect 5721 1207 5779 1213
rect 5721 1173 5733 1207
rect 5767 1204 5779 1207
rect 10318 1204 10324 1216
rect 5767 1176 10324 1204
rect 5767 1173 5779 1176
rect 5721 1167 5779 1173
rect 10318 1164 10324 1176
rect 10376 1164 10382 1216
rect 10502 1164 10508 1216
rect 10560 1164 10566 1216
rect 14734 1164 14740 1216
rect 14792 1204 14798 1216
rect 14921 1207 14979 1213
rect 14921 1204 14933 1207
rect 14792 1176 14933 1204
rect 14792 1164 14798 1176
rect 14921 1173 14933 1176
rect 14967 1173 14979 1207
rect 14921 1167 14979 1173
rect 16301 1207 16359 1213
rect 16301 1173 16313 1207
rect 16347 1204 16359 1207
rect 17604 1204 17632 1312
rect 18046 1300 18052 1312
rect 18104 1300 18110 1352
rect 17764 1275 17822 1281
rect 17764 1241 17776 1275
rect 17810 1272 17822 1275
rect 18414 1272 18420 1284
rect 17810 1244 18420 1272
rect 17810 1241 17822 1244
rect 17764 1235 17822 1241
rect 18414 1232 18420 1244
rect 18472 1232 18478 1284
rect 19306 1272 19334 1516
rect 22112 1516 22560 1544
rect 21450 1408 21456 1420
rect 21100 1380 21456 1408
rect 21100 1352 21128 1380
rect 21450 1368 21456 1380
rect 21508 1368 21514 1420
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19576 1312 19901 1340
rect 19576 1300 19582 1312
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 20257 1343 20315 1349
rect 20257 1309 20269 1343
rect 20303 1340 20315 1343
rect 20530 1340 20536 1352
rect 20303 1312 20536 1340
rect 20303 1309 20315 1312
rect 20257 1303 20315 1309
rect 20530 1300 20536 1312
rect 20588 1300 20594 1352
rect 20898 1300 20904 1352
rect 20956 1300 20962 1352
rect 21082 1300 21088 1352
rect 21140 1300 21146 1352
rect 21269 1343 21327 1349
rect 21269 1309 21281 1343
rect 21315 1340 21327 1343
rect 22112 1340 22140 1516
rect 22554 1504 22560 1516
rect 22612 1544 22618 1556
rect 25958 1544 25964 1556
rect 22612 1516 25964 1544
rect 22612 1504 22618 1516
rect 25958 1504 25964 1516
rect 26016 1504 26022 1556
rect 21315 1312 22140 1340
rect 21315 1309 21327 1312
rect 21269 1303 21327 1309
rect 22278 1300 22284 1352
rect 22336 1340 22342 1352
rect 22373 1343 22431 1349
rect 22373 1340 22385 1343
rect 22336 1312 22385 1340
rect 22336 1300 22342 1312
rect 22373 1309 22385 1312
rect 22419 1309 22431 1343
rect 22373 1303 22431 1309
rect 22640 1343 22698 1349
rect 22640 1309 22652 1343
rect 22686 1340 22698 1343
rect 23382 1340 23388 1352
rect 22686 1312 23388 1340
rect 22686 1309 22698 1312
rect 22640 1303 22698 1309
rect 23382 1300 23388 1312
rect 23440 1300 23446 1352
rect 25225 1343 25283 1349
rect 25225 1309 25237 1343
rect 25271 1340 25283 1343
rect 26970 1340 26976 1352
rect 25271 1312 26976 1340
rect 25271 1309 25283 1312
rect 25225 1303 25283 1309
rect 26970 1300 26976 1312
rect 27028 1300 27034 1352
rect 20073 1275 20131 1281
rect 20073 1272 20085 1275
rect 19306 1244 20085 1272
rect 20073 1241 20085 1244
rect 20119 1241 20131 1275
rect 20073 1235 20131 1241
rect 20162 1232 20168 1284
rect 20220 1232 20226 1284
rect 21177 1275 21235 1281
rect 21177 1241 21189 1275
rect 21223 1272 21235 1275
rect 24026 1272 24032 1284
rect 21223 1244 24032 1272
rect 21223 1241 21235 1244
rect 21177 1235 21235 1241
rect 24026 1232 24032 1244
rect 24084 1232 24090 1284
rect 25038 1232 25044 1284
rect 25096 1272 25102 1284
rect 25470 1275 25528 1281
rect 25470 1272 25482 1275
rect 25096 1244 25482 1272
rect 25096 1232 25102 1244
rect 25470 1241 25482 1244
rect 25516 1241 25528 1275
rect 25470 1235 25528 1241
rect 16347 1176 17632 1204
rect 16347 1173 16359 1176
rect 16301 1167 16359 1173
rect 17862 1164 17868 1216
rect 17920 1204 17926 1216
rect 18877 1207 18935 1213
rect 18877 1204 18889 1207
rect 17920 1176 18889 1204
rect 17920 1164 17926 1176
rect 18877 1173 18889 1176
rect 18923 1173 18935 1207
rect 18877 1167 18935 1173
rect 19242 1164 19248 1216
rect 19300 1204 19306 1216
rect 20441 1207 20499 1213
rect 20441 1204 20453 1207
rect 19300 1176 20453 1204
rect 19300 1164 19306 1176
rect 20441 1173 20453 1176
rect 20487 1173 20499 1207
rect 20441 1167 20499 1173
rect 20622 1164 20628 1216
rect 20680 1204 20686 1216
rect 21453 1207 21511 1213
rect 21453 1204 21465 1207
rect 20680 1176 21465 1204
rect 20680 1164 20686 1176
rect 21453 1173 21465 1176
rect 21499 1173 21511 1207
rect 21453 1167 21511 1173
rect 23750 1164 23756 1216
rect 23808 1164 23814 1216
rect 25774 1164 25780 1216
rect 25832 1204 25838 1216
rect 26605 1207 26663 1213
rect 26605 1204 26617 1207
rect 25832 1176 26617 1204
rect 25832 1164 25838 1176
rect 26605 1173 26617 1176
rect 26651 1173 26663 1207
rect 26605 1167 26663 1173
rect 1104 1114 29048 1136
rect 1104 1062 7896 1114
rect 7948 1062 7960 1114
rect 8012 1062 8024 1114
rect 8076 1062 8088 1114
rect 8140 1062 8152 1114
rect 8204 1062 14842 1114
rect 14894 1062 14906 1114
rect 14958 1062 14970 1114
rect 15022 1062 15034 1114
rect 15086 1062 15098 1114
rect 15150 1062 21788 1114
rect 21840 1062 21852 1114
rect 21904 1062 21916 1114
rect 21968 1062 21980 1114
rect 22032 1062 22044 1114
rect 22096 1062 28734 1114
rect 28786 1062 28798 1114
rect 28850 1062 28862 1114
rect 28914 1062 28926 1114
rect 28978 1062 28990 1114
rect 29042 1062 29048 1114
rect 1104 1040 29048 1062
rect 15930 960 15936 1012
rect 15988 1000 15994 1012
rect 21082 1000 21088 1012
rect 15988 972 21088 1000
rect 15988 960 15994 972
rect 21082 960 21088 972
rect 21140 960 21146 1012
rect 23750 1000 23756 1012
rect 22066 972 23756 1000
rect 19702 892 19708 944
rect 19760 932 19766 944
rect 22066 932 22094 972
rect 23750 960 23756 972
rect 23808 960 23814 1012
rect 19760 904 22094 932
rect 19760 892 19766 904
rect 20162 824 20168 876
rect 20220 864 20226 876
rect 23658 864 23664 876
rect 20220 836 23664 864
rect 20220 824 20226 836
rect 23658 824 23664 836
rect 23716 824 23722 876
<< via1 >>
rect 7896 32614 7948 32666
rect 7960 32614 8012 32666
rect 8024 32614 8076 32666
rect 8088 32614 8140 32666
rect 8152 32614 8204 32666
rect 14842 32614 14894 32666
rect 14906 32614 14958 32666
rect 14970 32614 15022 32666
rect 15034 32614 15086 32666
rect 15098 32614 15150 32666
rect 21788 32614 21840 32666
rect 21852 32614 21904 32666
rect 21916 32614 21968 32666
rect 21980 32614 22032 32666
rect 22044 32614 22096 32666
rect 28734 32614 28786 32666
rect 28798 32614 28850 32666
rect 28862 32614 28914 32666
rect 28926 32614 28978 32666
rect 28990 32614 29042 32666
rect 4344 32555 4396 32564
rect 4344 32521 4353 32555
rect 4353 32521 4387 32555
rect 4387 32521 4396 32555
rect 4344 32512 4396 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 8576 32555 8628 32564
rect 8576 32521 8585 32555
rect 8585 32521 8619 32555
rect 8619 32521 8628 32555
rect 8576 32512 8628 32521
rect 9496 32555 9548 32564
rect 9496 32521 9505 32555
rect 9505 32521 9539 32555
rect 9539 32521 9548 32555
rect 9496 32512 9548 32521
rect 11244 32512 11296 32564
rect 8484 32444 8536 32496
rect 1676 32376 1728 32428
rect 5172 32376 5224 32428
rect 8300 32376 8352 32428
rect 12532 32419 12584 32428
rect 12532 32385 12541 32419
rect 12541 32385 12575 32419
rect 12575 32385 12584 32419
rect 12532 32376 12584 32385
rect 14280 32419 14332 32428
rect 14280 32385 14289 32419
rect 14289 32385 14323 32419
rect 14323 32385 14332 32419
rect 14280 32376 14332 32385
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 4804 32351 4856 32360
rect 4804 32317 4813 32351
rect 4813 32317 4847 32351
rect 4847 32317 4856 32351
rect 4804 32308 4856 32317
rect 8208 32351 8260 32360
rect 8208 32317 8217 32351
rect 8217 32317 8251 32351
rect 8251 32317 8260 32351
rect 8208 32308 8260 32317
rect 9496 32351 9548 32360
rect 9496 32317 9505 32351
rect 9505 32317 9539 32351
rect 9539 32317 9548 32351
rect 9496 32308 9548 32317
rect 11152 32308 11204 32360
rect 3332 32240 3384 32292
rect 5172 32283 5224 32292
rect 5172 32249 5181 32283
rect 5181 32249 5215 32283
rect 5215 32249 5224 32283
rect 5172 32240 5224 32249
rect 8392 32240 8444 32292
rect 8576 32283 8628 32292
rect 8576 32249 8585 32283
rect 8585 32249 8619 32283
rect 8619 32249 8628 32283
rect 8576 32240 8628 32249
rect 4896 32172 4948 32224
rect 10140 32215 10192 32224
rect 10140 32181 10149 32215
rect 10149 32181 10183 32215
rect 10183 32181 10192 32215
rect 10140 32172 10192 32181
rect 11244 32240 11296 32292
rect 15752 32419 15804 32428
rect 15752 32385 15761 32419
rect 15761 32385 15795 32419
rect 15795 32385 15804 32419
rect 15752 32376 15804 32385
rect 13084 32172 13136 32224
rect 15108 32172 15160 32224
rect 4423 32070 4475 32122
rect 4487 32070 4539 32122
rect 4551 32070 4603 32122
rect 4615 32070 4667 32122
rect 4679 32070 4731 32122
rect 11369 32070 11421 32122
rect 11433 32070 11485 32122
rect 11497 32070 11549 32122
rect 11561 32070 11613 32122
rect 11625 32070 11677 32122
rect 18315 32070 18367 32122
rect 18379 32070 18431 32122
rect 18443 32070 18495 32122
rect 18507 32070 18559 32122
rect 18571 32070 18623 32122
rect 25261 32070 25313 32122
rect 25325 32070 25377 32122
rect 25389 32070 25441 32122
rect 25453 32070 25505 32122
rect 25517 32070 25569 32122
rect 2780 31968 2832 32020
rect 5264 31968 5316 32020
rect 3332 31875 3384 31884
rect 3332 31841 3341 31875
rect 3341 31841 3375 31875
rect 3375 31841 3384 31875
rect 3332 31832 3384 31841
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 5172 31900 5224 31952
rect 12532 31968 12584 32020
rect 9036 31832 9088 31884
rect 11888 31900 11940 31952
rect 9496 31832 9548 31884
rect 10968 31832 11020 31884
rect 4436 31807 4488 31816
rect 4436 31773 4439 31807
rect 4439 31773 4488 31807
rect 4436 31764 4488 31773
rect 4804 31764 4856 31816
rect 7564 31764 7616 31816
rect 8208 31807 8260 31816
rect 8208 31773 8217 31807
rect 8217 31773 8251 31807
rect 8251 31773 8260 31807
rect 8208 31764 8260 31773
rect 8576 31807 8628 31816
rect 8576 31773 8585 31807
rect 8585 31773 8619 31807
rect 8619 31773 8628 31807
rect 8576 31764 8628 31773
rect 4712 31696 4764 31748
rect 5908 31671 5960 31680
rect 5908 31637 5917 31671
rect 5917 31637 5951 31671
rect 5951 31637 5960 31671
rect 5908 31628 5960 31637
rect 11152 31764 11204 31816
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 11704 31832 11756 31884
rect 10232 31671 10284 31680
rect 10232 31637 10241 31671
rect 10241 31637 10275 31671
rect 10275 31637 10284 31671
rect 10232 31628 10284 31637
rect 12348 31807 12400 31816
rect 12348 31773 12357 31807
rect 12357 31773 12391 31807
rect 12391 31773 12400 31807
rect 12348 31764 12400 31773
rect 13084 31764 13136 31816
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 15108 31807 15160 31816
rect 15108 31773 15117 31807
rect 15117 31773 15151 31807
rect 15151 31773 15160 31807
rect 15108 31764 15160 31773
rect 16396 31807 16448 31816
rect 16396 31773 16405 31807
rect 16405 31773 16439 31807
rect 16439 31773 16448 31807
rect 16396 31764 16448 31773
rect 12164 31628 12216 31680
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 5080 31424 5132 31476
rect 5908 31424 5960 31476
rect 6920 31424 6972 31476
rect 1492 31288 1544 31340
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 2596 31331 2648 31340
rect 2596 31297 2605 31331
rect 2605 31297 2639 31331
rect 2639 31297 2648 31331
rect 2596 31288 2648 31297
rect 4804 31331 4856 31340
rect 4804 31297 4813 31331
rect 4813 31297 4847 31331
rect 4847 31297 4856 31331
rect 4804 31288 4856 31297
rect 6552 31288 6604 31340
rect 7656 31288 7708 31340
rect 10232 31424 10284 31476
rect 11152 31467 11204 31476
rect 11152 31433 11161 31467
rect 11161 31433 11195 31467
rect 11195 31433 11204 31467
rect 12072 31467 12124 31476
rect 11152 31424 11204 31433
rect 12072 31433 12081 31467
rect 12081 31433 12115 31467
rect 12115 31433 12124 31467
rect 12072 31424 12124 31433
rect 13728 31424 13780 31476
rect 11060 31356 11112 31408
rect 12348 31356 12400 31408
rect 11152 31331 11204 31340
rect 11152 31297 11161 31331
rect 11161 31297 11195 31331
rect 11195 31297 11204 31331
rect 11152 31288 11204 31297
rect 11980 31288 12032 31340
rect 3884 31220 3936 31272
rect 7564 31220 7616 31272
rect 9956 31263 10008 31272
rect 9956 31229 9965 31263
rect 9965 31229 9999 31263
rect 9999 31229 10008 31263
rect 9956 31220 10008 31229
rect 11520 31220 11572 31272
rect 12164 31220 12216 31272
rect 13176 31220 13228 31272
rect 5172 31195 5224 31204
rect 5172 31161 5181 31195
rect 5181 31161 5215 31195
rect 5215 31161 5224 31195
rect 5172 31152 5224 31161
rect 5908 31152 5960 31204
rect 12072 31195 12124 31204
rect 12072 31161 12081 31195
rect 12081 31161 12115 31195
rect 12115 31161 12124 31195
rect 12072 31152 12124 31161
rect 14372 31152 14424 31204
rect 15200 31152 15252 31204
rect 3792 31084 3844 31136
rect 4252 31084 4304 31136
rect 4436 31084 4488 31136
rect 6368 31084 6420 31136
rect 12624 31084 12676 31136
rect 14004 31084 14056 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 2596 30880 2648 30932
rect 7656 30923 7708 30932
rect 7656 30889 7665 30923
rect 7665 30889 7699 30923
rect 7699 30889 7708 30923
rect 7656 30880 7708 30889
rect 8300 30812 8352 30864
rect 12072 30880 12124 30932
rect 5632 30744 5684 30796
rect 7564 30744 7616 30796
rect 9588 30812 9640 30864
rect 9956 30744 10008 30796
rect 11060 30744 11112 30796
rect 4252 30719 4304 30728
rect 4252 30685 4261 30719
rect 4261 30685 4295 30719
rect 4295 30685 4304 30719
rect 4252 30676 4304 30685
rect 4344 30676 4396 30728
rect 6552 30676 6604 30728
rect 7656 30719 7708 30728
rect 7656 30685 7665 30719
rect 7665 30685 7699 30719
rect 7699 30685 7708 30719
rect 7656 30676 7708 30685
rect 6000 30608 6052 30660
rect 4160 30540 4212 30592
rect 9588 30540 9640 30592
rect 14372 30744 14424 30796
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 13176 30676 13228 30728
rect 14004 30676 14056 30728
rect 15200 30719 15252 30728
rect 15200 30685 15209 30719
rect 15209 30685 15243 30719
rect 15243 30685 15252 30719
rect 15200 30676 15252 30685
rect 13268 30608 13320 30660
rect 12716 30540 12768 30592
rect 13176 30540 13228 30592
rect 13728 30583 13780 30592
rect 13728 30549 13737 30583
rect 13737 30549 13771 30583
rect 13771 30549 13780 30583
rect 13728 30540 13780 30549
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 6920 30379 6972 30388
rect 6920 30345 6929 30379
rect 6929 30345 6963 30379
rect 6963 30345 6972 30379
rect 6920 30336 6972 30345
rect 1860 30268 1912 30320
rect 3976 30268 4028 30320
rect 2136 30243 2188 30252
rect 2136 30209 2145 30243
rect 2145 30209 2179 30243
rect 2179 30209 2188 30243
rect 2136 30200 2188 30209
rect 2228 30243 2280 30252
rect 2228 30209 2237 30243
rect 2237 30209 2271 30243
rect 2271 30209 2280 30243
rect 2228 30200 2280 30209
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 2872 30243 2924 30252
rect 2872 30209 2881 30243
rect 2881 30209 2915 30243
rect 2915 30209 2924 30243
rect 2872 30200 2924 30209
rect 7472 30268 7524 30320
rect 5448 30243 5500 30252
rect 5448 30209 5457 30243
rect 5457 30209 5491 30243
rect 5491 30209 5500 30243
rect 5448 30200 5500 30209
rect 6184 30200 6236 30252
rect 6552 30243 6604 30252
rect 6552 30209 6561 30243
rect 6561 30209 6595 30243
rect 6595 30209 6604 30243
rect 6552 30200 6604 30209
rect 7564 30200 7616 30252
rect 9956 30243 10008 30252
rect 9956 30209 9965 30243
rect 9965 30209 9999 30243
rect 9999 30209 10008 30243
rect 9956 30200 10008 30209
rect 11060 30200 11112 30252
rect 12716 30379 12768 30388
rect 12716 30345 12725 30379
rect 12725 30345 12759 30379
rect 12759 30345 12768 30379
rect 12716 30336 12768 30345
rect 13728 30336 13780 30388
rect 11704 30243 11756 30252
rect 11704 30209 11713 30243
rect 11713 30209 11747 30243
rect 11747 30209 11756 30243
rect 11704 30200 11756 30209
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 14004 30243 14056 30252
rect 14004 30209 14013 30243
rect 14013 30209 14047 30243
rect 14047 30209 14056 30243
rect 14832 30243 14884 30252
rect 14004 30200 14056 30209
rect 14832 30209 14841 30243
rect 14841 30209 14875 30243
rect 14875 30209 14884 30243
rect 14832 30200 14884 30209
rect 5632 30175 5684 30184
rect 5632 30141 5641 30175
rect 5641 30141 5675 30175
rect 5675 30141 5684 30175
rect 5632 30132 5684 30141
rect 13176 30175 13228 30184
rect 4344 30064 4396 30116
rect 5080 30064 5132 30116
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 14372 30175 14424 30184
rect 6920 30107 6972 30116
rect 6920 30073 6929 30107
rect 6929 30073 6963 30107
rect 6963 30073 6972 30107
rect 6920 30064 6972 30073
rect 7656 30064 7708 30116
rect 12900 30064 12952 30116
rect 14372 30141 14381 30175
rect 14381 30141 14415 30175
rect 14415 30141 14424 30175
rect 14372 30132 14424 30141
rect 13820 30064 13872 30116
rect 15200 30107 15252 30116
rect 15200 30073 15209 30107
rect 15209 30073 15243 30107
rect 15243 30073 15252 30107
rect 15200 30064 15252 30073
rect 1584 29996 1636 30048
rect 2504 29996 2556 30048
rect 4252 29996 4304 30048
rect 10416 29996 10468 30048
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 5172 29792 5224 29844
rect 2228 29724 2280 29776
rect 4252 29724 4304 29776
rect 7380 29792 7432 29844
rect 14464 29792 14516 29844
rect 1952 29588 2004 29640
rect 2412 29588 2464 29640
rect 4252 29631 4304 29640
rect 4252 29597 4261 29631
rect 4261 29597 4295 29631
rect 4295 29597 4304 29631
rect 4252 29588 4304 29597
rect 3884 29520 3936 29572
rect 5908 29724 5960 29776
rect 6920 29724 6972 29776
rect 11060 29724 11112 29776
rect 12900 29767 12952 29776
rect 12900 29733 12909 29767
rect 12909 29733 12943 29767
rect 12943 29733 12952 29767
rect 12900 29724 12952 29733
rect 9956 29699 10008 29708
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 10692 29656 10744 29708
rect 14832 29699 14884 29708
rect 14832 29665 14841 29699
rect 14841 29665 14875 29699
rect 14875 29665 14884 29699
rect 14832 29656 14884 29665
rect 5540 29588 5592 29640
rect 6460 29588 6512 29640
rect 7472 29631 7524 29640
rect 7472 29597 7481 29631
rect 7481 29597 7515 29631
rect 7515 29597 7524 29631
rect 7472 29588 7524 29597
rect 7564 29588 7616 29640
rect 8300 29631 8352 29640
rect 8300 29597 8344 29631
rect 8344 29597 8352 29631
rect 8300 29588 8352 29597
rect 1584 29452 1636 29504
rect 3424 29452 3476 29504
rect 5816 29520 5868 29572
rect 5632 29495 5684 29504
rect 5632 29461 5641 29495
rect 5641 29461 5675 29495
rect 5675 29461 5684 29495
rect 5632 29452 5684 29461
rect 6828 29452 6880 29504
rect 11060 29452 11112 29504
rect 11888 29520 11940 29572
rect 13176 29588 13228 29640
rect 13820 29588 13872 29640
rect 15200 29631 15252 29640
rect 15200 29597 15209 29631
rect 15209 29597 15243 29631
rect 15243 29597 15252 29631
rect 15200 29588 15252 29597
rect 14188 29520 14240 29572
rect 12716 29452 12768 29504
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 1768 29248 1820 29300
rect 2412 29180 2464 29232
rect 2872 29248 2924 29300
rect 11060 29291 11112 29300
rect 11060 29257 11069 29291
rect 11069 29257 11103 29291
rect 11103 29257 11112 29291
rect 11060 29248 11112 29257
rect 5632 29180 5684 29232
rect 16396 29248 16448 29300
rect 2596 29155 2648 29164
rect 2596 29121 2605 29155
rect 2605 29121 2639 29155
rect 2639 29121 2648 29155
rect 2596 29112 2648 29121
rect 5448 29155 5500 29164
rect 5448 29121 5457 29155
rect 5457 29121 5491 29155
rect 5491 29121 5500 29155
rect 5448 29112 5500 29121
rect 6920 29155 6972 29164
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 6920 29112 6972 29121
rect 3976 29044 4028 29096
rect 6736 29044 6788 29096
rect 7012 29087 7064 29096
rect 7012 29053 7021 29087
rect 7021 29053 7055 29087
rect 7055 29053 7064 29087
rect 7012 29044 7064 29053
rect 14372 29180 14424 29232
rect 10692 29155 10744 29164
rect 10692 29121 10701 29155
rect 10701 29121 10735 29155
rect 10735 29121 10744 29155
rect 10692 29112 10744 29121
rect 11060 29155 11112 29164
rect 11060 29121 11069 29155
rect 11069 29121 11103 29155
rect 11103 29121 11112 29155
rect 11060 29112 11112 29121
rect 11704 29155 11756 29164
rect 11704 29121 11713 29155
rect 11713 29121 11747 29155
rect 11747 29121 11756 29155
rect 11704 29112 11756 29121
rect 5540 28976 5592 29028
rect 6092 28976 6144 29028
rect 5724 28908 5776 28960
rect 6644 28908 6696 28960
rect 7656 28976 7708 29028
rect 9312 29019 9364 29028
rect 9312 28985 9321 29019
rect 9321 28985 9355 29019
rect 9355 28985 9364 29019
rect 9312 28976 9364 28985
rect 10140 28976 10192 29028
rect 13820 29112 13872 29164
rect 12348 29087 12400 29096
rect 12348 29053 12357 29087
rect 12357 29053 12391 29087
rect 12391 29053 12400 29087
rect 12348 29044 12400 29053
rect 14188 29087 14240 29096
rect 14188 29053 14197 29087
rect 14197 29053 14231 29087
rect 14231 29053 14240 29087
rect 14188 29044 14240 29053
rect 15200 29019 15252 29028
rect 15200 28985 15209 29019
rect 15209 28985 15243 29019
rect 15243 28985 15252 29019
rect 15200 28976 15252 28985
rect 11060 28908 11112 28960
rect 12716 28951 12768 28960
rect 12716 28917 12725 28951
rect 12725 28917 12759 28951
rect 12759 28917 12768 28951
rect 12716 28908 12768 28917
rect 13820 28908 13872 28960
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 7564 28704 7616 28756
rect 15752 28704 15804 28756
rect 5172 28636 5224 28688
rect 7288 28636 7340 28688
rect 8392 28636 8444 28688
rect 2044 28543 2096 28552
rect 2044 28509 2053 28543
rect 2053 28509 2087 28543
rect 2087 28509 2096 28543
rect 2044 28500 2096 28509
rect 3424 28500 3476 28552
rect 9128 28568 9180 28620
rect 9496 28568 9548 28620
rect 2688 28432 2740 28484
rect 6092 28543 6144 28552
rect 6092 28509 6101 28543
rect 6101 28509 6135 28543
rect 6135 28509 6144 28543
rect 6092 28500 6144 28509
rect 6644 28543 6696 28552
rect 6644 28509 6653 28543
rect 6653 28509 6687 28543
rect 6687 28509 6696 28543
rect 6644 28500 6696 28509
rect 4344 28432 4396 28484
rect 7564 28543 7616 28552
rect 7564 28509 7573 28543
rect 7573 28509 7607 28543
rect 7607 28509 7616 28543
rect 7564 28500 7616 28509
rect 9588 28500 9640 28552
rect 14372 28636 14424 28688
rect 12716 28611 12768 28620
rect 12716 28577 12725 28611
rect 12725 28577 12759 28611
rect 12759 28577 12768 28611
rect 12716 28568 12768 28577
rect 12348 28543 12400 28552
rect 3516 28364 3568 28416
rect 5172 28364 5224 28416
rect 5448 28364 5500 28416
rect 7472 28407 7524 28416
rect 7472 28373 7481 28407
rect 7481 28373 7515 28407
rect 7515 28373 7524 28407
rect 7472 28364 7524 28373
rect 7748 28432 7800 28484
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 11704 28432 11756 28484
rect 8576 28364 8628 28416
rect 11796 28364 11848 28416
rect 14188 28568 14240 28620
rect 13820 28364 13872 28416
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 4160 28160 4212 28212
rect 4252 28160 4304 28212
rect 8852 28160 8904 28212
rect 1676 28024 1728 28076
rect 1952 28024 2004 28076
rect 3424 28092 3476 28144
rect 5908 28135 5960 28144
rect 5908 28101 5917 28135
rect 5917 28101 5951 28135
rect 5951 28101 5960 28135
rect 5908 28092 5960 28101
rect 6920 28092 6972 28144
rect 2504 28024 2556 28076
rect 3516 28024 3568 28076
rect 4252 27956 4304 28008
rect 4988 28067 5040 28076
rect 4988 28033 4997 28067
rect 4997 28033 5031 28067
rect 5031 28033 5040 28067
rect 4988 28024 5040 28033
rect 5724 28067 5776 28076
rect 5724 28033 5733 28067
rect 5733 28033 5767 28067
rect 5767 28033 5776 28067
rect 5724 28024 5776 28033
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 7472 28024 7524 28076
rect 7196 27956 7248 28008
rect 8300 27956 8352 28008
rect 10048 27956 10100 28008
rect 12348 28024 12400 28076
rect 13176 28067 13228 28076
rect 13176 28033 13185 28067
rect 13185 28033 13219 28067
rect 13219 28033 13228 28067
rect 13176 28024 13228 28033
rect 17592 28024 17644 28076
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 14556 27956 14608 28008
rect 8944 27931 8996 27940
rect 8944 27897 8953 27931
rect 8953 27897 8987 27931
rect 8987 27897 8996 27931
rect 8944 27888 8996 27897
rect 13728 27888 13780 27940
rect 6920 27863 6972 27872
rect 6920 27829 6929 27863
rect 6929 27829 6963 27863
rect 6963 27829 6972 27863
rect 6920 27820 6972 27829
rect 12992 27863 13044 27872
rect 12992 27829 13001 27863
rect 13001 27829 13035 27863
rect 13035 27829 13044 27863
rect 12992 27820 13044 27829
rect 16304 27863 16356 27872
rect 16304 27829 16313 27863
rect 16313 27829 16347 27863
rect 16347 27829 16356 27863
rect 16304 27820 16356 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 2596 27616 2648 27668
rect 4068 27616 4120 27668
rect 6552 27616 6604 27668
rect 8852 27616 8904 27668
rect 10600 27659 10652 27668
rect 10600 27625 10609 27659
rect 10609 27625 10643 27659
rect 10643 27625 10652 27659
rect 10600 27616 10652 27625
rect 6092 27548 6144 27600
rect 9036 27548 9088 27600
rect 2044 27412 2096 27464
rect 8576 27480 8628 27532
rect 11796 27616 11848 27668
rect 11980 27523 12032 27532
rect 11980 27489 11989 27523
rect 11989 27489 12023 27523
rect 12023 27489 12032 27523
rect 11980 27480 12032 27489
rect 4068 27455 4120 27464
rect 4068 27421 4077 27455
rect 4077 27421 4111 27455
rect 4111 27421 4120 27455
rect 4068 27412 4120 27421
rect 3976 27344 4028 27396
rect 5632 27412 5684 27464
rect 4160 27276 4212 27328
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 8484 27412 8536 27464
rect 10600 27455 10652 27464
rect 10600 27421 10609 27455
rect 10609 27421 10643 27455
rect 10643 27421 10652 27455
rect 10600 27412 10652 27421
rect 11888 27455 11940 27464
rect 11888 27421 11897 27455
rect 11897 27421 11931 27455
rect 11931 27421 11940 27455
rect 11888 27412 11940 27421
rect 7748 27344 7800 27396
rect 9404 27344 9456 27396
rect 13176 27412 13228 27464
rect 18328 27412 18380 27464
rect 10140 27276 10192 27328
rect 14372 27276 14424 27328
rect 14464 27276 14516 27328
rect 20720 27455 20772 27464
rect 20720 27421 20729 27455
rect 20729 27421 20763 27455
rect 20763 27421 20772 27455
rect 20720 27412 20772 27421
rect 20260 27344 20312 27396
rect 22560 27276 22612 27328
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 1860 27072 1912 27124
rect 4068 27072 4120 27124
rect 4160 27072 4212 27124
rect 7472 27072 7524 27124
rect 7564 27072 7616 27124
rect 9404 27072 9456 27124
rect 11704 27115 11756 27124
rect 11704 27081 11713 27115
rect 11713 27081 11747 27115
rect 11747 27081 11756 27115
rect 11704 27072 11756 27081
rect 13544 27115 13596 27124
rect 13544 27081 13553 27115
rect 13553 27081 13587 27115
rect 13587 27081 13596 27115
rect 13544 27072 13596 27081
rect 13820 27072 13872 27124
rect 14464 27072 14516 27124
rect 2688 26936 2740 26988
rect 5448 27004 5500 27056
rect 7104 27004 7156 27056
rect 1860 26911 1912 26920
rect 1860 26877 1869 26911
rect 1869 26877 1903 26911
rect 1903 26877 1912 26911
rect 1860 26868 1912 26877
rect 2412 26868 2464 26920
rect 4712 26911 4764 26920
rect 4712 26877 4721 26911
rect 4721 26877 4755 26911
rect 4755 26877 4764 26911
rect 4712 26868 4764 26877
rect 5172 26800 5224 26852
rect 6092 26936 6144 26988
rect 6368 26936 6420 26988
rect 7656 27004 7708 27056
rect 6460 26868 6512 26920
rect 7748 26936 7800 26988
rect 20720 27004 20772 27056
rect 12072 26979 12124 26988
rect 12072 26945 12081 26979
rect 12081 26945 12115 26979
rect 12115 26945 12124 26979
rect 12072 26936 12124 26945
rect 12992 26936 13044 26988
rect 13728 26936 13780 26988
rect 14372 26979 14424 26988
rect 14372 26945 14381 26979
rect 14381 26945 14415 26979
rect 14415 26945 14424 26979
rect 14372 26936 14424 26945
rect 18328 26979 18380 26988
rect 18328 26945 18337 26979
rect 18337 26945 18371 26979
rect 18371 26945 18380 26979
rect 18328 26936 18380 26945
rect 19156 26979 19208 26988
rect 19156 26945 19165 26979
rect 19165 26945 19199 26979
rect 19199 26945 19208 26979
rect 19156 26936 19208 26945
rect 20628 26936 20680 26988
rect 22836 26936 22888 26988
rect 8300 26868 8352 26920
rect 10048 26868 10100 26920
rect 12716 26868 12768 26920
rect 21824 26868 21876 26920
rect 9864 26800 9916 26852
rect 4160 26775 4212 26784
rect 4160 26741 4169 26775
rect 4169 26741 4203 26775
rect 4203 26741 4212 26775
rect 4160 26732 4212 26741
rect 4712 26732 4764 26784
rect 5632 26732 5684 26784
rect 5724 26732 5776 26784
rect 8208 26732 8260 26784
rect 20260 26732 20312 26784
rect 24400 26775 24452 26784
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 2412 26528 2464 26580
rect 5356 26503 5408 26512
rect 5356 26469 5365 26503
rect 5365 26469 5399 26503
rect 5399 26469 5408 26503
rect 5356 26460 5408 26469
rect 2044 26392 2096 26444
rect 2688 26392 2740 26444
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 4252 26367 4304 26376
rect 4252 26333 4286 26367
rect 4286 26333 4304 26367
rect 4252 26324 4304 26333
rect 7104 26460 7156 26512
rect 8300 26528 8352 26580
rect 8852 26528 8904 26580
rect 9588 26571 9640 26580
rect 9588 26537 9597 26571
rect 9597 26537 9631 26571
rect 9631 26537 9640 26571
rect 9588 26528 9640 26537
rect 13544 26571 13596 26580
rect 13544 26537 13553 26571
rect 13553 26537 13587 26571
rect 13587 26537 13596 26571
rect 13544 26528 13596 26537
rect 17592 26571 17644 26580
rect 17592 26537 17601 26571
rect 17601 26537 17635 26571
rect 17635 26537 17644 26571
rect 17592 26528 17644 26537
rect 22836 26528 22888 26580
rect 9956 26460 10008 26512
rect 5540 26392 5592 26444
rect 8208 26435 8260 26444
rect 8208 26401 8217 26435
rect 8217 26401 8251 26435
rect 8251 26401 8260 26435
rect 8208 26392 8260 26401
rect 6000 26367 6052 26376
rect 6000 26333 6009 26367
rect 6009 26333 6043 26367
rect 6043 26333 6052 26367
rect 6000 26324 6052 26333
rect 4804 26256 4856 26308
rect 6736 26299 6788 26308
rect 6736 26265 6745 26299
rect 6745 26265 6779 26299
rect 6779 26265 6788 26299
rect 6736 26256 6788 26265
rect 8484 26324 8536 26376
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 9680 26324 9732 26376
rect 10048 26324 10100 26376
rect 8852 26256 8904 26308
rect 12992 26392 13044 26444
rect 21456 26392 21508 26444
rect 21824 26435 21876 26444
rect 21824 26401 21833 26435
rect 21833 26401 21867 26435
rect 21867 26401 21876 26435
rect 21824 26392 21876 26401
rect 12716 26367 12768 26376
rect 12716 26333 12725 26367
rect 12725 26333 12759 26367
rect 12759 26333 12768 26367
rect 12716 26324 12768 26333
rect 18328 26324 18380 26376
rect 25136 26324 25188 26376
rect 10232 26256 10284 26308
rect 2688 26188 2740 26240
rect 5356 26188 5408 26240
rect 9772 26188 9824 26240
rect 10048 26231 10100 26240
rect 10048 26197 10057 26231
rect 10057 26197 10091 26231
rect 10091 26197 10100 26231
rect 10048 26188 10100 26197
rect 12072 26188 12124 26240
rect 12164 26188 12216 26240
rect 17408 26256 17460 26308
rect 22560 26256 22612 26308
rect 25044 26256 25096 26308
rect 26148 26256 26200 26308
rect 17684 26188 17736 26240
rect 18328 26188 18380 26240
rect 19156 26188 19208 26240
rect 23204 26231 23256 26240
rect 23204 26197 23213 26231
rect 23213 26197 23247 26231
rect 23247 26197 23256 26231
rect 23204 26188 23256 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 5356 25984 5408 26036
rect 5448 25984 5500 26036
rect 1676 25891 1728 25900
rect 1676 25857 1685 25891
rect 1685 25857 1719 25891
rect 1719 25857 1728 25891
rect 1676 25848 1728 25857
rect 4068 25848 4120 25900
rect 5632 25891 5684 25900
rect 5632 25857 5641 25891
rect 5641 25857 5675 25891
rect 5675 25857 5684 25891
rect 5632 25848 5684 25857
rect 6552 25959 6604 25968
rect 6552 25925 6561 25959
rect 6561 25925 6595 25959
rect 6595 25925 6604 25959
rect 6552 25916 6604 25925
rect 6828 26027 6880 26036
rect 6828 25993 6837 26027
rect 6837 25993 6871 26027
rect 6871 25993 6880 26027
rect 6828 25984 6880 25993
rect 8944 26027 8996 26036
rect 8944 25993 8953 26027
rect 8953 25993 8987 26027
rect 8987 25993 8996 26027
rect 8944 25984 8996 25993
rect 9772 25984 9824 26036
rect 11796 25984 11848 26036
rect 13544 26027 13596 26036
rect 13544 25993 13553 26027
rect 13553 25993 13587 26027
rect 13587 25993 13596 26027
rect 13544 25984 13596 25993
rect 26148 25984 26200 26036
rect 7196 25916 7248 25968
rect 9220 25916 9272 25968
rect 12348 25916 12400 25968
rect 13268 25916 13320 25968
rect 16580 25916 16632 25968
rect 19248 25916 19300 25968
rect 25596 25916 25648 25968
rect 6920 25848 6972 25900
rect 7104 25891 7156 25900
rect 7104 25857 7113 25891
rect 7113 25857 7147 25891
rect 7147 25857 7156 25891
rect 7104 25848 7156 25857
rect 8852 25891 8904 25900
rect 8852 25857 8861 25891
rect 8861 25857 8895 25891
rect 8895 25857 8904 25891
rect 8852 25848 8904 25857
rect 10416 25848 10468 25900
rect 10968 25891 11020 25900
rect 10968 25857 10977 25891
rect 10977 25857 11011 25891
rect 11011 25857 11020 25891
rect 10968 25848 11020 25857
rect 12716 25848 12768 25900
rect 12992 25848 13044 25900
rect 16028 25891 16080 25900
rect 16028 25857 16037 25891
rect 16037 25857 16071 25891
rect 16071 25857 16080 25891
rect 16028 25848 16080 25857
rect 17224 25848 17276 25900
rect 18328 25891 18380 25900
rect 18328 25857 18337 25891
rect 18337 25857 18371 25891
rect 18371 25857 18380 25891
rect 18328 25848 18380 25857
rect 2044 25780 2096 25832
rect 4804 25823 4856 25832
rect 4804 25789 4813 25823
rect 4813 25789 4847 25823
rect 4847 25789 4856 25823
rect 4804 25780 4856 25789
rect 4988 25823 5040 25832
rect 4988 25789 4997 25823
rect 4997 25789 5031 25823
rect 5031 25789 5040 25823
rect 4988 25780 5040 25789
rect 5172 25780 5224 25832
rect 25136 25780 25188 25832
rect 3976 25644 4028 25696
rect 4252 25712 4304 25764
rect 12624 25712 12676 25764
rect 5632 25644 5684 25696
rect 6000 25644 6052 25696
rect 12256 25644 12308 25696
rect 15844 25687 15896 25696
rect 15844 25653 15853 25687
rect 15853 25653 15887 25687
rect 15887 25653 15896 25687
rect 15844 25644 15896 25653
rect 19708 25687 19760 25696
rect 19708 25653 19717 25687
rect 19717 25653 19751 25687
rect 19751 25653 19760 25687
rect 19708 25644 19760 25653
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 1952 25440 2004 25492
rect 3424 25440 3476 25492
rect 5816 25440 5868 25492
rect 4988 25304 5040 25356
rect 5172 25304 5224 25356
rect 2044 25279 2096 25288
rect 2044 25245 2053 25279
rect 2053 25245 2087 25279
rect 2087 25245 2096 25279
rect 2044 25236 2096 25245
rect 4252 25236 4304 25288
rect 5356 25236 5408 25288
rect 5816 25304 5868 25356
rect 7104 25440 7156 25492
rect 7380 25440 7432 25492
rect 8576 25440 8628 25492
rect 11888 25440 11940 25492
rect 17684 25440 17736 25492
rect 7012 25372 7064 25424
rect 8208 25372 8260 25424
rect 8484 25372 8536 25424
rect 10416 25372 10468 25424
rect 7656 25304 7708 25356
rect 8576 25304 8628 25356
rect 7196 25236 7248 25288
rect 4528 25211 4580 25220
rect 4528 25177 4537 25211
rect 4537 25177 4571 25211
rect 4571 25177 4580 25211
rect 4528 25168 4580 25177
rect 6092 25211 6144 25220
rect 6092 25177 6101 25211
rect 6101 25177 6135 25211
rect 6135 25177 6144 25211
rect 6092 25168 6144 25177
rect 8300 25279 8352 25288
rect 8300 25245 8309 25279
rect 8309 25245 8343 25279
rect 8343 25245 8352 25279
rect 12256 25347 12308 25356
rect 12256 25313 12265 25347
rect 12265 25313 12299 25347
rect 12299 25313 12308 25347
rect 12256 25304 12308 25313
rect 8300 25236 8352 25245
rect 7656 25168 7708 25220
rect 8944 25168 8996 25220
rect 9680 25168 9732 25220
rect 11704 25168 11756 25220
rect 8208 25100 8260 25152
rect 10048 25100 10100 25152
rect 10968 25100 11020 25152
rect 12072 25211 12124 25220
rect 12072 25177 12107 25211
rect 12107 25177 12124 25211
rect 12348 25236 12400 25288
rect 25964 25483 26016 25492
rect 25964 25449 25973 25483
rect 25973 25449 26007 25483
rect 26007 25449 26016 25483
rect 25964 25440 26016 25449
rect 26976 25279 27028 25288
rect 26976 25245 26985 25279
rect 26985 25245 27019 25279
rect 27019 25245 27028 25279
rect 26976 25236 27028 25245
rect 12072 25168 12124 25177
rect 12440 25168 12492 25220
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 25688 25211 25740 25220
rect 25688 25177 25697 25211
rect 25697 25177 25731 25211
rect 25731 25177 25740 25211
rect 25688 25168 25740 25177
rect 27252 25211 27304 25220
rect 27252 25177 27286 25211
rect 27286 25177 27304 25211
rect 27252 25168 27304 25177
rect 27528 25100 27580 25152
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 3792 24896 3844 24948
rect 3148 24871 3200 24880
rect 3148 24837 3157 24871
rect 3157 24837 3191 24871
rect 3191 24837 3200 24871
rect 3148 24828 3200 24837
rect 2688 24760 2740 24812
rect 2964 24803 3016 24812
rect 2964 24769 2973 24803
rect 2973 24769 3007 24803
rect 3007 24769 3016 24803
rect 2964 24760 3016 24769
rect 3884 24760 3936 24812
rect 4528 24896 4580 24948
rect 5632 24896 5684 24948
rect 6092 24896 6144 24948
rect 7656 24896 7708 24948
rect 10232 24939 10284 24948
rect 10232 24905 10241 24939
rect 10241 24905 10275 24939
rect 10275 24905 10284 24939
rect 10232 24896 10284 24905
rect 11060 24896 11112 24948
rect 4620 24803 4672 24812
rect 4620 24769 4629 24803
rect 4629 24769 4663 24803
rect 4663 24769 4672 24803
rect 4620 24760 4672 24769
rect 7564 24828 7616 24880
rect 12164 24828 12216 24880
rect 12440 24828 12492 24880
rect 1860 24692 1912 24744
rect 4988 24692 5040 24744
rect 4068 24624 4120 24676
rect 4620 24624 4672 24676
rect 4896 24624 4948 24676
rect 5448 24760 5500 24812
rect 5816 24760 5868 24812
rect 10140 24760 10192 24812
rect 7748 24692 7800 24744
rect 10968 24760 11020 24812
rect 11060 24760 11112 24812
rect 11796 24760 11848 24812
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 6184 24624 6236 24676
rect 10508 24692 10560 24744
rect 11980 24692 12032 24744
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 16488 24760 16540 24812
rect 17040 24803 17092 24812
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 15568 24692 15620 24744
rect 16028 24692 16080 24744
rect 10232 24624 10284 24676
rect 9680 24556 9732 24608
rect 12716 24599 12768 24608
rect 12716 24565 12725 24599
rect 12725 24565 12759 24599
rect 12759 24565 12768 24599
rect 12716 24556 12768 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 2136 24352 2188 24404
rect 3884 24352 3936 24404
rect 9312 24352 9364 24404
rect 10232 24395 10284 24404
rect 10232 24361 10241 24395
rect 10241 24361 10275 24395
rect 10275 24361 10284 24395
rect 10232 24352 10284 24361
rect 16580 24395 16632 24404
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 16580 24352 16632 24361
rect 1492 24148 1544 24200
rect 848 24080 900 24132
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 2228 24148 2280 24200
rect 2320 24191 2372 24200
rect 2320 24157 2329 24191
rect 2329 24157 2363 24191
rect 2363 24157 2372 24191
rect 2320 24148 2372 24157
rect 4160 24284 4212 24336
rect 4344 24284 4396 24336
rect 3148 24216 3200 24268
rect 10692 24284 10744 24336
rect 11704 24216 11756 24268
rect 11980 24216 12032 24268
rect 2688 24148 2740 24200
rect 4528 24191 4580 24200
rect 4528 24157 4537 24191
rect 4537 24157 4571 24191
rect 4571 24157 4580 24191
rect 4528 24148 4580 24157
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 1860 24012 1912 24064
rect 2044 24012 2096 24064
rect 4068 24080 4120 24132
rect 5724 24148 5776 24200
rect 8300 24148 8352 24200
rect 9956 24148 10008 24200
rect 10508 24148 10560 24200
rect 12072 24148 12124 24200
rect 12256 24148 12308 24200
rect 2320 24012 2372 24064
rect 4528 24012 4580 24064
rect 6276 24080 6328 24132
rect 6644 24080 6696 24132
rect 10968 24080 11020 24132
rect 12624 24080 12676 24132
rect 20720 24216 20772 24268
rect 13268 24148 13320 24200
rect 16488 24191 16540 24200
rect 16488 24157 16497 24191
rect 16497 24157 16531 24191
rect 16531 24157 16540 24191
rect 16488 24148 16540 24157
rect 16120 24080 16172 24132
rect 17040 24148 17092 24200
rect 24584 24148 24636 24200
rect 25136 24148 25188 24200
rect 26976 24191 27028 24200
rect 26976 24157 26985 24191
rect 26985 24157 27019 24191
rect 27019 24157 27028 24191
rect 26976 24148 27028 24157
rect 19156 24080 19208 24132
rect 23204 24080 23256 24132
rect 27344 24080 27396 24132
rect 5724 24012 5776 24064
rect 21548 24012 21600 24064
rect 24124 24012 24176 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 4988 23808 5040 23860
rect 5448 23808 5500 23860
rect 6368 23808 6420 23860
rect 7012 23808 7064 23860
rect 7840 23851 7892 23860
rect 7840 23817 7849 23851
rect 7849 23817 7883 23851
rect 7883 23817 7892 23851
rect 7840 23808 7892 23817
rect 8300 23808 8352 23860
rect 2596 23783 2648 23792
rect 2596 23749 2605 23783
rect 2605 23749 2639 23783
rect 2639 23749 2648 23783
rect 2596 23740 2648 23749
rect 4712 23740 4764 23792
rect 3608 23672 3660 23724
rect 4988 23672 5040 23724
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5816 23740 5868 23792
rect 7104 23740 7156 23792
rect 10600 23740 10652 23792
rect 5264 23672 5316 23681
rect 5448 23715 5500 23724
rect 5448 23681 5457 23715
rect 5457 23681 5491 23715
rect 5491 23681 5500 23715
rect 5448 23672 5500 23681
rect 7196 23672 7248 23724
rect 9772 23672 9824 23724
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 11152 23672 11204 23724
rect 5816 23604 5868 23656
rect 6460 23604 6512 23656
rect 8392 23536 8444 23588
rect 10140 23604 10192 23656
rect 10508 23604 10560 23656
rect 12256 23604 12308 23656
rect 14740 23740 14792 23792
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 16304 23672 16356 23724
rect 21180 23604 21232 23656
rect 24400 23740 24452 23792
rect 24584 23604 24636 23656
rect 4160 23468 4212 23520
rect 6460 23468 6512 23520
rect 6644 23468 6696 23520
rect 6920 23511 6972 23520
rect 6920 23477 6929 23511
rect 6929 23477 6963 23511
rect 6963 23477 6972 23511
rect 6920 23468 6972 23477
rect 7840 23468 7892 23520
rect 12072 23468 12124 23520
rect 15568 23468 15620 23520
rect 16028 23468 16080 23520
rect 26056 23468 26108 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 1584 23264 1636 23316
rect 11704 23264 11756 23316
rect 11980 23264 12032 23316
rect 12348 23264 12400 23316
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 5356 23196 5408 23248
rect 9036 23196 9088 23248
rect 9956 23196 10008 23248
rect 5540 23128 5592 23180
rect 5632 23171 5684 23180
rect 5632 23137 5641 23171
rect 5641 23137 5675 23171
rect 5675 23137 5684 23171
rect 5632 23128 5684 23137
rect 6184 23128 6236 23180
rect 6644 23128 6696 23180
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 10416 23128 10468 23180
rect 24584 23128 24636 23180
rect 4160 22992 4212 23044
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 10600 23060 10652 23112
rect 10876 23060 10928 23112
rect 12348 23103 12400 23112
rect 12348 23069 12357 23103
rect 12357 23069 12391 23103
rect 12391 23069 12400 23103
rect 12348 23060 12400 23069
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 18236 23060 18288 23112
rect 20720 23060 20772 23112
rect 6184 22992 6236 23044
rect 12900 22992 12952 23044
rect 14556 22992 14608 23044
rect 17960 22992 18012 23044
rect 6644 22924 6696 22976
rect 9680 22924 9732 22976
rect 12808 22967 12860 22976
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 13360 22967 13412 22976
rect 13360 22933 13369 22967
rect 13369 22933 13403 22967
rect 13403 22933 13412 22967
rect 13360 22924 13412 22933
rect 18144 22924 18196 22976
rect 21640 22924 21692 22976
rect 26056 22924 26108 22976
rect 27252 22967 27304 22976
rect 27252 22933 27261 22967
rect 27261 22933 27295 22967
rect 27295 22933 27304 22967
rect 27252 22924 27304 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 4896 22720 4948 22772
rect 10508 22720 10560 22772
rect 11704 22763 11756 22772
rect 11704 22729 11713 22763
rect 11713 22729 11747 22763
rect 11747 22729 11756 22763
rect 11704 22720 11756 22729
rect 13360 22720 13412 22772
rect 13728 22652 13780 22704
rect 4896 22584 4948 22636
rect 2504 22516 2556 22568
rect 6644 22516 6696 22568
rect 1400 22380 1452 22432
rect 7012 22627 7064 22636
rect 7012 22593 7021 22627
rect 7021 22593 7055 22627
rect 7055 22593 7064 22627
rect 7012 22584 7064 22593
rect 7196 22584 7248 22636
rect 7380 22516 7432 22568
rect 9404 22584 9456 22636
rect 11704 22584 11756 22636
rect 12072 22584 12124 22636
rect 12164 22627 12216 22636
rect 12164 22593 12173 22627
rect 12173 22593 12207 22627
rect 12207 22593 12216 22627
rect 12164 22584 12216 22593
rect 12900 22627 12952 22636
rect 12900 22593 12909 22627
rect 12909 22593 12943 22627
rect 12943 22593 12952 22627
rect 12900 22584 12952 22593
rect 16028 22720 16080 22772
rect 17960 22720 18012 22772
rect 18788 22720 18840 22772
rect 20720 22652 20772 22704
rect 20076 22584 20128 22636
rect 21640 22584 21692 22636
rect 23388 22584 23440 22636
rect 23940 22652 23992 22704
rect 24124 22695 24176 22704
rect 24124 22661 24158 22695
rect 24158 22661 24176 22695
rect 24124 22652 24176 22661
rect 24584 22584 24636 22636
rect 11704 22380 11756 22432
rect 13912 22448 13964 22500
rect 14096 22380 14148 22432
rect 15752 22380 15804 22432
rect 20628 22380 20680 22432
rect 25136 22380 25188 22432
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 7012 22176 7064 22228
rect 10876 22176 10928 22228
rect 11244 22176 11296 22228
rect 9772 22108 9824 22160
rect 10048 22108 10100 22160
rect 10416 22108 10468 22160
rect 1952 22083 2004 22092
rect 1952 22049 1961 22083
rect 1961 22049 1995 22083
rect 1995 22049 2004 22083
rect 1952 22040 2004 22049
rect 5080 22040 5132 22092
rect 7288 22040 7340 22092
rect 7380 22040 7432 22092
rect 8576 22040 8628 22092
rect 9956 22040 10008 22092
rect 12808 22040 12860 22092
rect 24584 22083 24636 22092
rect 24584 22049 24593 22083
rect 24593 22049 24627 22083
rect 24627 22049 24636 22083
rect 24584 22040 24636 22049
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2136 22015 2188 22024
rect 2136 21981 2145 22015
rect 2145 21981 2179 22015
rect 2179 21981 2188 22015
rect 2136 21972 2188 21981
rect 2320 22015 2372 22024
rect 2320 21981 2329 22015
rect 2329 21981 2363 22015
rect 2363 21981 2372 22015
rect 2320 21972 2372 21981
rect 4068 21972 4120 22024
rect 5724 21972 5776 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 6736 22015 6788 22024
rect 6736 21981 6745 22015
rect 6745 21981 6779 22015
rect 6779 21981 6788 22015
rect 6736 21972 6788 21981
rect 3884 21904 3936 21956
rect 6920 21904 6972 21956
rect 7288 21904 7340 21956
rect 7472 21904 7524 21956
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 5356 21879 5408 21888
rect 5356 21845 5365 21879
rect 5365 21845 5399 21879
rect 5399 21845 5408 21879
rect 5356 21836 5408 21845
rect 7012 21836 7064 21888
rect 7840 21836 7892 21888
rect 8852 21836 8904 21888
rect 9128 21836 9180 21888
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 12072 21904 12124 21956
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 12440 21836 12492 21888
rect 14188 21836 14240 21888
rect 18236 21972 18288 22024
rect 21640 21972 21692 22024
rect 25964 21972 26016 22024
rect 18144 21904 18196 21956
rect 24492 21904 24544 21956
rect 25136 21904 25188 21956
rect 26884 21904 26936 21956
rect 27528 21904 27580 21956
rect 17776 21879 17828 21888
rect 17776 21845 17785 21879
rect 17785 21845 17819 21879
rect 17819 21845 17828 21879
rect 17776 21836 17828 21845
rect 20168 21836 20220 21888
rect 21548 21836 21600 21888
rect 22284 21836 22336 21888
rect 23296 21836 23348 21888
rect 26148 21836 26200 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 2320 21632 2372 21684
rect 6552 21632 6604 21684
rect 13636 21632 13688 21684
rect 2136 21564 2188 21616
rect 3148 21539 3200 21548
rect 3148 21505 3157 21539
rect 3157 21505 3191 21539
rect 3191 21505 3200 21539
rect 3148 21496 3200 21505
rect 4344 21496 4396 21548
rect 5816 21496 5868 21548
rect 6644 21496 6696 21548
rect 7104 21496 7156 21548
rect 7196 21496 7248 21548
rect 5264 21360 5316 21412
rect 11704 21496 11756 21548
rect 9220 21428 9272 21480
rect 9404 21428 9456 21480
rect 7104 21292 7156 21344
rect 9496 21292 9548 21344
rect 10600 21292 10652 21344
rect 17776 21632 17828 21684
rect 12256 21496 12308 21548
rect 18696 21564 18748 21616
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 20536 21564 20588 21616
rect 21456 21564 21508 21616
rect 23112 21564 23164 21616
rect 20352 21539 20404 21548
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 15844 21428 15896 21437
rect 20352 21505 20386 21539
rect 20386 21505 20404 21539
rect 20352 21496 20404 21505
rect 23296 21496 23348 21548
rect 23480 21539 23532 21548
rect 23480 21505 23514 21539
rect 23514 21505 23532 21539
rect 23480 21496 23532 21505
rect 25964 21564 26016 21616
rect 15292 21360 15344 21412
rect 15660 21360 15712 21412
rect 19340 21428 19392 21480
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 19248 21292 19300 21344
rect 19800 21292 19852 21344
rect 20076 21292 20128 21344
rect 22744 21292 22796 21344
rect 24860 21292 24912 21344
rect 25596 21292 25648 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 6920 21088 6972 21140
rect 7196 21088 7248 21140
rect 10232 21088 10284 21140
rect 11060 21088 11112 21140
rect 12348 21088 12400 21140
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 1492 20748 1544 20800
rect 5356 20748 5408 20800
rect 6276 20859 6328 20868
rect 6276 20825 6285 20859
rect 6285 20825 6319 20859
rect 6319 20825 6328 20859
rect 6276 20816 6328 20825
rect 7288 20884 7340 20936
rect 9312 20884 9364 20936
rect 6920 20748 6972 20800
rect 7196 20816 7248 20868
rect 9588 20859 9640 20868
rect 9588 20825 9597 20859
rect 9597 20825 9631 20859
rect 9631 20825 9640 20859
rect 9588 20816 9640 20825
rect 9772 20859 9824 20868
rect 9772 20825 9781 20859
rect 9781 20825 9815 20859
rect 9815 20825 9824 20859
rect 9772 20816 9824 20825
rect 7288 20791 7340 20800
rect 7288 20757 7297 20791
rect 7297 20757 7331 20791
rect 7331 20757 7340 20791
rect 7288 20748 7340 20757
rect 7472 20748 7524 20800
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 11152 20884 11204 20936
rect 12992 20884 13044 20936
rect 11612 20859 11664 20868
rect 11612 20825 11646 20859
rect 11646 20825 11664 20859
rect 11612 20816 11664 20825
rect 11704 20816 11756 20868
rect 16488 21088 16540 21140
rect 14188 20952 14240 21004
rect 11796 20748 11848 20800
rect 13820 20748 13872 20800
rect 16764 20884 16816 20936
rect 19340 20884 19392 20936
rect 20720 20884 20772 20936
rect 22744 21088 22796 21140
rect 23204 20884 23256 20936
rect 25964 20884 26016 20936
rect 15568 20816 15620 20868
rect 22376 20816 22428 20868
rect 25136 20816 25188 20868
rect 16212 20748 16264 20800
rect 18052 20748 18104 20800
rect 21640 20748 21692 20800
rect 23848 20791 23900 20800
rect 23848 20757 23857 20791
rect 23857 20757 23891 20791
rect 23891 20757 23900 20791
rect 23848 20748 23900 20757
rect 26516 20748 26568 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 4252 20544 4304 20596
rect 5172 20544 5224 20596
rect 5448 20544 5500 20596
rect 6276 20544 6328 20596
rect 6828 20544 6880 20596
rect 10324 20544 10376 20596
rect 10508 20587 10560 20596
rect 10508 20553 10517 20587
rect 10517 20553 10551 20587
rect 10551 20553 10560 20587
rect 10508 20544 10560 20553
rect 12164 20544 12216 20596
rect 16120 20587 16172 20596
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 3240 20476 3292 20528
rect 4988 20408 5040 20460
rect 4252 20383 4304 20392
rect 4252 20349 4261 20383
rect 4261 20349 4295 20383
rect 4295 20349 4304 20383
rect 4252 20340 4304 20349
rect 4804 20340 4856 20392
rect 5448 20340 5500 20392
rect 5908 20408 5960 20460
rect 8116 20476 8168 20528
rect 9680 20476 9732 20528
rect 10416 20476 10468 20528
rect 12716 20476 12768 20528
rect 13912 20476 13964 20528
rect 7472 20451 7524 20460
rect 7472 20417 7481 20451
rect 7481 20417 7515 20451
rect 7515 20417 7524 20451
rect 7472 20408 7524 20417
rect 6276 20340 6328 20392
rect 7104 20340 7156 20392
rect 9312 20408 9364 20460
rect 9496 20451 9548 20460
rect 9496 20417 9505 20451
rect 9505 20417 9539 20451
rect 9539 20417 9548 20451
rect 9496 20408 9548 20417
rect 14188 20408 14240 20460
rect 15568 20408 15620 20460
rect 6736 20272 6788 20324
rect 7748 20272 7800 20324
rect 4804 20204 4856 20256
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 10508 20340 10560 20392
rect 11060 20340 11112 20392
rect 11612 20340 11664 20392
rect 11980 20383 12032 20392
rect 11980 20349 11989 20383
rect 11989 20349 12023 20383
rect 12023 20349 12032 20383
rect 11980 20340 12032 20349
rect 9588 20204 9640 20256
rect 10416 20204 10468 20256
rect 10876 20272 10928 20324
rect 12164 20383 12216 20392
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 12256 20340 12308 20392
rect 15660 20340 15712 20392
rect 16764 20340 16816 20392
rect 19340 20476 19392 20528
rect 18236 20408 18288 20460
rect 21640 20476 21692 20528
rect 19892 20408 19944 20460
rect 23204 20476 23256 20528
rect 22284 20451 22336 20460
rect 22284 20417 22318 20451
rect 22318 20417 22336 20451
rect 22284 20408 22336 20417
rect 25964 20476 26016 20528
rect 24400 20408 24452 20460
rect 19984 20383 20036 20392
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 15936 20315 15988 20324
rect 15936 20281 15945 20315
rect 15945 20281 15979 20315
rect 15979 20281 15988 20315
rect 15936 20272 15988 20281
rect 11980 20204 12032 20256
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 16396 20204 16448 20256
rect 23664 20272 23716 20324
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 25136 20204 25188 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 4988 20000 5040 20052
rect 5632 20000 5684 20052
rect 5724 20043 5776 20052
rect 5724 20009 5733 20043
rect 5733 20009 5767 20043
rect 5767 20009 5776 20043
rect 5724 20000 5776 20009
rect 6092 20000 6144 20052
rect 7196 20000 7248 20052
rect 8852 20000 8904 20052
rect 9680 20000 9732 20052
rect 9864 20000 9916 20052
rect 10232 20043 10284 20052
rect 10232 20009 10241 20043
rect 10241 20009 10275 20043
rect 10275 20009 10284 20043
rect 10232 20000 10284 20009
rect 10416 20000 10468 20052
rect 10784 20000 10836 20052
rect 17132 20000 17184 20052
rect 17408 20000 17460 20052
rect 23204 20000 23256 20052
rect 23480 20000 23532 20052
rect 2228 19932 2280 19984
rect 7656 19932 7708 19984
rect 5172 19864 5224 19916
rect 5356 19796 5408 19848
rect 5540 19864 5592 19916
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 12440 19932 12492 19984
rect 9864 19864 9916 19916
rect 10876 19864 10928 19916
rect 16764 19907 16816 19916
rect 16764 19873 16773 19907
rect 16773 19873 16807 19907
rect 16807 19873 16816 19907
rect 16764 19864 16816 19873
rect 19984 19864 20036 19916
rect 3332 19660 3384 19712
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 6552 19771 6604 19780
rect 6552 19737 6561 19771
rect 6561 19737 6595 19771
rect 6595 19737 6604 19771
rect 6552 19728 6604 19737
rect 5632 19660 5684 19712
rect 7104 19728 7156 19780
rect 6736 19703 6788 19712
rect 6736 19669 6761 19703
rect 6761 19669 6788 19703
rect 6736 19660 6788 19669
rect 7196 19660 7248 19712
rect 7840 19660 7892 19712
rect 8116 19728 8168 19780
rect 9864 19771 9916 19780
rect 9864 19737 9873 19771
rect 9873 19737 9907 19771
rect 9907 19737 9916 19771
rect 9864 19728 9916 19737
rect 10968 19796 11020 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 20720 19796 20772 19848
rect 22652 19839 22704 19848
rect 22652 19805 22661 19839
rect 22661 19805 22695 19839
rect 22695 19805 22704 19839
rect 22652 19796 22704 19805
rect 25964 19796 26016 19848
rect 26976 19796 27028 19848
rect 10140 19728 10192 19780
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 11520 19728 11572 19780
rect 12348 19728 12400 19780
rect 15568 19728 15620 19780
rect 16396 19728 16448 19780
rect 19064 19728 19116 19780
rect 23388 19728 23440 19780
rect 25780 19728 25832 19780
rect 10416 19660 10468 19712
rect 11336 19703 11388 19712
rect 11336 19669 11345 19703
rect 11345 19669 11379 19703
rect 11379 19669 11388 19703
rect 11336 19660 11388 19669
rect 13268 19660 13320 19712
rect 15660 19660 15712 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 22652 19660 22704 19712
rect 25228 19660 25280 19712
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 3700 19456 3752 19508
rect 3976 19388 4028 19440
rect 7380 19388 7432 19440
rect 7656 19456 7708 19508
rect 10048 19456 10100 19508
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 10784 19456 10836 19508
rect 10140 19388 10192 19440
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 5172 19320 5224 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 3424 19184 3476 19236
rect 5080 19252 5132 19304
rect 6644 19252 6696 19304
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 7656 19320 7708 19372
rect 8668 19320 8720 19372
rect 9312 19320 9364 19372
rect 6368 19184 6420 19236
rect 8116 19184 8168 19236
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 9772 19252 9824 19304
rect 10692 19320 10744 19372
rect 11060 19388 11112 19440
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 11244 19388 11296 19440
rect 12256 19388 12308 19440
rect 11888 19320 11940 19372
rect 14004 19456 14056 19508
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 13636 19320 13688 19372
rect 15660 19456 15712 19508
rect 16212 19456 16264 19508
rect 16764 19456 16816 19508
rect 19340 19456 19392 19508
rect 23296 19456 23348 19508
rect 15568 19431 15620 19440
rect 15568 19397 15577 19431
rect 15577 19397 15611 19431
rect 15611 19397 15620 19431
rect 15568 19388 15620 19397
rect 17224 19431 17276 19440
rect 17224 19397 17233 19431
rect 17233 19397 17267 19431
rect 17267 19397 17276 19431
rect 17224 19388 17276 19397
rect 16948 19320 17000 19372
rect 17040 19320 17092 19372
rect 22468 19388 22520 19440
rect 23388 19388 23440 19440
rect 9956 19184 10008 19236
rect 17224 19252 17276 19304
rect 23204 19320 23256 19372
rect 24952 19320 25004 19372
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 11888 19184 11940 19236
rect 12992 19184 13044 19236
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 5264 19116 5316 19168
rect 8484 19116 8536 19168
rect 9772 19116 9824 19168
rect 11520 19116 11572 19168
rect 16120 19116 16172 19168
rect 19248 19184 19300 19236
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 25964 19116 26016 19168
rect 26332 19116 26384 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 4344 18955 4396 18964
rect 4344 18921 4353 18955
rect 4353 18921 4387 18955
rect 4387 18921 4396 18955
rect 4344 18912 4396 18921
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 7104 18912 7156 18964
rect 8484 18912 8536 18964
rect 10416 18912 10468 18964
rect 14004 18912 14056 18964
rect 16028 18912 16080 18964
rect 20444 18912 20496 18964
rect 4804 18844 4856 18896
rect 3056 18776 3108 18828
rect 4344 18776 4396 18828
rect 4896 18776 4948 18828
rect 5540 18776 5592 18828
rect 5908 18776 5960 18828
rect 3516 18640 3568 18692
rect 5816 18708 5868 18760
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 7288 18776 7340 18828
rect 8300 18776 8352 18828
rect 10968 18844 11020 18896
rect 14648 18844 14700 18896
rect 17960 18844 18012 18896
rect 20812 18844 20864 18896
rect 23572 18844 23624 18896
rect 8116 18708 8168 18760
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 7472 18640 7524 18692
rect 7748 18640 7800 18692
rect 8484 18640 8536 18692
rect 8852 18640 8904 18692
rect 4988 18572 5040 18624
rect 5908 18615 5960 18624
rect 5908 18581 5917 18615
rect 5917 18581 5951 18615
rect 5951 18581 5960 18615
rect 5908 18572 5960 18581
rect 6644 18615 6696 18624
rect 6644 18581 6653 18615
rect 6653 18581 6687 18615
rect 6687 18581 6696 18615
rect 6644 18572 6696 18581
rect 7564 18572 7616 18624
rect 10416 18640 10468 18692
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 10140 18572 10192 18624
rect 10876 18572 10928 18624
rect 11244 18708 11296 18760
rect 16120 18776 16172 18828
rect 12808 18708 12860 18760
rect 14280 18708 14332 18760
rect 15384 18708 15436 18760
rect 16580 18776 16632 18828
rect 18788 18776 18840 18828
rect 12900 18640 12952 18692
rect 14004 18640 14056 18692
rect 16120 18640 16172 18692
rect 16304 18683 16356 18692
rect 16304 18649 16313 18683
rect 16313 18649 16347 18683
rect 16347 18649 16356 18683
rect 16304 18640 16356 18649
rect 16580 18640 16632 18692
rect 16672 18640 16724 18692
rect 17224 18640 17276 18692
rect 18880 18708 18932 18760
rect 20076 18751 20128 18760
rect 20076 18717 20085 18751
rect 20085 18717 20119 18751
rect 20119 18717 20128 18751
rect 20076 18708 20128 18717
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 17408 18640 17460 18692
rect 17592 18640 17644 18692
rect 20720 18708 20772 18760
rect 25044 18776 25096 18828
rect 25964 18776 26016 18828
rect 21456 18708 21508 18760
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 23480 18708 23532 18760
rect 13912 18572 13964 18624
rect 14740 18572 14792 18624
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 18236 18572 18288 18624
rect 21272 18640 21324 18692
rect 19984 18572 20036 18624
rect 20720 18572 20772 18624
rect 22192 18572 22244 18624
rect 24768 18640 24820 18692
rect 26332 18640 26384 18692
rect 27160 18572 27212 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 2964 18368 3016 18420
rect 6000 18368 6052 18420
rect 6184 18368 6236 18420
rect 9864 18368 9916 18420
rect 8852 18300 8904 18352
rect 8944 18343 8996 18352
rect 8944 18309 8953 18343
rect 8953 18309 8987 18343
rect 8987 18309 8996 18343
rect 8944 18300 8996 18309
rect 9956 18300 10008 18352
rect 12624 18368 12676 18420
rect 13084 18368 13136 18420
rect 15476 18368 15528 18420
rect 3332 18232 3384 18284
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 3424 18164 3476 18216
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 6552 18028 6604 18080
rect 7196 18232 7248 18284
rect 8668 18232 8720 18284
rect 9312 18232 9364 18284
rect 13820 18300 13872 18352
rect 14096 18300 14148 18352
rect 16028 18300 16080 18352
rect 10416 18275 10468 18284
rect 10416 18241 10426 18275
rect 10426 18241 10460 18275
rect 10460 18241 10468 18275
rect 10416 18232 10468 18241
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 10968 18232 11020 18284
rect 14556 18232 14608 18284
rect 15476 18232 15528 18284
rect 12716 18164 12768 18216
rect 8576 18096 8628 18148
rect 16212 18096 16264 18148
rect 16580 18096 16632 18148
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17316 18275 17368 18284
rect 17316 18241 17351 18275
rect 17351 18241 17368 18275
rect 17316 18232 17368 18241
rect 20076 18368 20128 18420
rect 20628 18300 20680 18352
rect 21364 18300 21416 18352
rect 22100 18300 22152 18352
rect 17960 18232 18012 18284
rect 18144 18275 18196 18284
rect 18144 18241 18154 18275
rect 18154 18241 18188 18275
rect 18188 18241 18196 18275
rect 18144 18232 18196 18241
rect 18236 18232 18288 18284
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 19340 18275 19392 18284
rect 19340 18241 19349 18275
rect 19349 18241 19383 18275
rect 19383 18241 19392 18275
rect 19340 18232 19392 18241
rect 21088 18232 21140 18284
rect 23480 18300 23532 18352
rect 23848 18300 23900 18352
rect 24768 18300 24820 18352
rect 26884 18300 26936 18352
rect 24860 18275 24912 18284
rect 24860 18241 24869 18275
rect 24869 18241 24903 18275
rect 24903 18241 24912 18275
rect 24860 18232 24912 18241
rect 17408 18096 17460 18148
rect 9680 18028 9732 18080
rect 10140 18028 10192 18080
rect 13452 18028 13504 18080
rect 14648 18028 14700 18080
rect 15936 18028 15988 18080
rect 17684 18028 17736 18080
rect 17960 18028 18012 18080
rect 23020 18207 23072 18216
rect 23020 18173 23029 18207
rect 23029 18173 23063 18207
rect 23063 18173 23072 18207
rect 23020 18164 23072 18173
rect 24124 18164 24176 18216
rect 20444 18028 20496 18080
rect 23940 18028 23992 18080
rect 24400 18071 24452 18080
rect 24400 18037 24409 18071
rect 24409 18037 24443 18071
rect 24443 18037 24452 18071
rect 24400 18028 24452 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 2688 17824 2740 17876
rect 3148 17824 3200 17876
rect 5724 17867 5776 17876
rect 5724 17833 5733 17867
rect 5733 17833 5767 17867
rect 5767 17833 5776 17867
rect 5724 17824 5776 17833
rect 6368 17824 6420 17876
rect 7288 17824 7340 17876
rect 10876 17824 10928 17876
rect 10416 17756 10468 17808
rect 1676 17688 1728 17740
rect 4252 17688 4304 17740
rect 4804 17688 4856 17740
rect 5724 17688 5776 17740
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 4988 17620 5040 17672
rect 6920 17688 6972 17740
rect 2596 17552 2648 17604
rect 5080 17484 5132 17536
rect 5448 17552 5500 17604
rect 6828 17620 6880 17672
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 6460 17595 6512 17604
rect 6460 17561 6469 17595
rect 6469 17561 6503 17595
rect 6503 17561 6512 17595
rect 8208 17620 8260 17672
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 10048 17620 10100 17672
rect 6460 17552 6512 17561
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 9496 17595 9548 17604
rect 9496 17561 9505 17595
rect 9505 17561 9539 17595
rect 9539 17561 9548 17595
rect 9496 17552 9548 17561
rect 6920 17484 6972 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 9128 17484 9180 17536
rect 9588 17484 9640 17536
rect 9680 17484 9732 17536
rect 10140 17484 10192 17536
rect 11152 17620 11204 17672
rect 12440 17824 12492 17876
rect 14188 17824 14240 17876
rect 18696 17824 18748 17876
rect 19616 17824 19668 17876
rect 22836 17824 22888 17876
rect 12256 17688 12308 17740
rect 12624 17663 12676 17672
rect 12624 17629 12633 17663
rect 12633 17629 12667 17663
rect 12667 17629 12676 17663
rect 12624 17620 12676 17629
rect 12900 17620 12952 17672
rect 13452 17731 13504 17740
rect 13452 17697 13461 17731
rect 13461 17697 13495 17731
rect 13495 17697 13504 17731
rect 13452 17688 13504 17697
rect 17040 17756 17092 17808
rect 24860 17756 24912 17808
rect 18880 17688 18932 17740
rect 12348 17595 12400 17604
rect 12348 17561 12357 17595
rect 12357 17561 12391 17595
rect 12391 17561 12400 17595
rect 12348 17552 12400 17561
rect 13176 17552 13228 17604
rect 14188 17552 14240 17604
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 14556 17620 14608 17672
rect 16856 17620 16908 17672
rect 18972 17620 19024 17672
rect 26976 17731 27028 17740
rect 26976 17697 26985 17731
rect 26985 17697 27019 17731
rect 27019 17697 27028 17731
rect 26976 17688 27028 17697
rect 20628 17620 20680 17672
rect 23020 17620 23072 17672
rect 25872 17620 25924 17672
rect 14004 17484 14056 17536
rect 14372 17484 14424 17536
rect 16028 17484 16080 17536
rect 16488 17552 16540 17604
rect 16672 17484 16724 17536
rect 16948 17484 17000 17536
rect 17408 17484 17460 17536
rect 20168 17552 20220 17604
rect 22100 17552 22152 17604
rect 22468 17552 22520 17604
rect 23940 17552 23992 17604
rect 17960 17484 18012 17536
rect 20904 17484 20956 17536
rect 20996 17484 21048 17536
rect 24032 17484 24084 17536
rect 26424 17527 26476 17536
rect 26424 17493 26433 17527
rect 26433 17493 26467 17527
rect 26467 17493 26476 17527
rect 26424 17484 26476 17493
rect 27528 17484 27580 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 3056 17280 3108 17332
rect 3240 17323 3292 17332
rect 3240 17289 3249 17323
rect 3249 17289 3283 17323
rect 3283 17289 3292 17323
rect 3240 17280 3292 17289
rect 3332 17280 3384 17332
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2596 17144 2648 17196
rect 2872 17144 2924 17196
rect 3516 17187 3568 17196
rect 3516 17153 3526 17187
rect 3526 17153 3560 17187
rect 3560 17153 3568 17187
rect 3516 17144 3568 17153
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 7012 17280 7064 17332
rect 8208 17323 8260 17332
rect 5080 17212 5132 17264
rect 6092 17212 6144 17264
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 7564 17212 7616 17264
rect 4804 17076 4856 17128
rect 6000 17144 6052 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 2688 17008 2740 17060
rect 5448 17008 5500 17060
rect 1952 16940 2004 16992
rect 3792 16940 3844 16992
rect 5080 16940 5132 16992
rect 6276 17076 6328 17128
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 10048 17280 10100 17332
rect 10324 17280 10376 17332
rect 12716 17323 12768 17332
rect 12716 17289 12725 17323
rect 12725 17289 12759 17323
rect 12759 17289 12768 17323
rect 12716 17280 12768 17289
rect 14188 17280 14240 17332
rect 14740 17280 14792 17332
rect 17592 17280 17644 17332
rect 10968 17212 11020 17264
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 14004 17212 14056 17264
rect 17960 17212 18012 17264
rect 8484 17144 8536 17196
rect 9496 17144 9548 17196
rect 7564 17076 7616 17085
rect 8484 17008 8536 17060
rect 5724 16940 5776 16992
rect 9956 17076 10008 17128
rect 12256 17144 12308 17196
rect 12348 17144 12400 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 14740 17144 14792 17196
rect 17040 17144 17092 17196
rect 17776 17144 17828 17196
rect 18696 17212 18748 17264
rect 14464 17076 14516 17128
rect 11704 17008 11756 17060
rect 14372 17008 14424 17060
rect 14648 17076 14700 17128
rect 11244 16940 11296 16992
rect 11980 16940 12032 16992
rect 14280 16940 14332 16992
rect 16120 17076 16172 17128
rect 19340 17212 19392 17264
rect 22284 17280 22336 17332
rect 20168 17187 20220 17196
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20444 17187 20496 17196
rect 23296 17212 23348 17264
rect 24952 17212 25004 17264
rect 26148 17212 26200 17264
rect 20444 17153 20479 17187
rect 20479 17153 20496 17187
rect 20444 17144 20496 17153
rect 20996 17144 21048 17196
rect 23664 17144 23716 17196
rect 25872 17144 25924 17196
rect 20904 17076 20956 17128
rect 21640 17076 21692 17128
rect 18052 17008 18104 17060
rect 17224 16940 17276 16992
rect 19892 17008 19944 17060
rect 20628 17008 20680 17060
rect 23296 17008 23348 17060
rect 24492 17008 24544 17060
rect 19156 16940 19208 16992
rect 19340 16940 19392 16992
rect 23020 16940 23072 16992
rect 23112 16940 23164 16992
rect 26884 16940 26936 16992
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 1676 16736 1728 16788
rect 5724 16736 5776 16788
rect 6184 16736 6236 16788
rect 6736 16736 6788 16788
rect 8208 16736 8260 16788
rect 10324 16736 10376 16788
rect 11152 16736 11204 16788
rect 11336 16736 11388 16788
rect 17132 16736 17184 16788
rect 18788 16736 18840 16788
rect 18880 16736 18932 16788
rect 19708 16736 19760 16788
rect 2596 16668 2648 16720
rect 4712 16668 4764 16720
rect 7104 16668 7156 16720
rect 2964 16600 3016 16652
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 5264 16600 5316 16652
rect 9128 16668 9180 16720
rect 9588 16668 9640 16720
rect 9772 16668 9824 16720
rect 664 16532 716 16584
rect 2228 16532 2280 16584
rect 2596 16532 2648 16584
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 4252 16532 4304 16584
rect 3148 16507 3200 16516
rect 3148 16473 3157 16507
rect 3157 16473 3191 16507
rect 3191 16473 3200 16507
rect 3148 16464 3200 16473
rect 6184 16532 6236 16584
rect 7104 16532 7156 16584
rect 5632 16507 5684 16516
rect 5632 16473 5641 16507
rect 5641 16473 5675 16507
rect 5675 16473 5684 16507
rect 5632 16464 5684 16473
rect 6000 16464 6052 16516
rect 6368 16464 6420 16516
rect 10232 16600 10284 16652
rect 7564 16532 7616 16584
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 8668 16532 8720 16584
rect 8300 16507 8352 16516
rect 8300 16473 8309 16507
rect 8309 16473 8343 16507
rect 8343 16473 8352 16507
rect 8300 16464 8352 16473
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 4804 16396 4856 16448
rect 6828 16396 6880 16448
rect 7012 16396 7064 16448
rect 7564 16396 7616 16448
rect 8944 16464 8996 16516
rect 9312 16532 9364 16584
rect 9588 16532 9640 16584
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10692 16532 10744 16584
rect 12532 16668 12584 16720
rect 17224 16668 17276 16720
rect 19156 16668 19208 16720
rect 12256 16600 12308 16652
rect 14740 16600 14792 16652
rect 16120 16600 16172 16652
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 17776 16532 17828 16584
rect 19524 16575 19576 16584
rect 19892 16668 19944 16720
rect 20444 16736 20496 16788
rect 20812 16779 20864 16788
rect 20812 16745 20821 16779
rect 20821 16745 20855 16779
rect 20855 16745 20864 16779
rect 20812 16736 20864 16745
rect 19524 16541 19540 16575
rect 19540 16541 19574 16575
rect 19574 16541 19576 16575
rect 19524 16532 19576 16541
rect 11888 16464 11940 16516
rect 15844 16464 15896 16516
rect 18880 16464 18932 16516
rect 11796 16396 11848 16448
rect 12072 16396 12124 16448
rect 15660 16396 15712 16448
rect 16304 16396 16356 16448
rect 17316 16396 17368 16448
rect 19432 16396 19484 16448
rect 20444 16532 20496 16584
rect 21088 16575 21140 16584
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 19708 16464 19760 16516
rect 20720 16464 20772 16516
rect 22100 16464 22152 16516
rect 22376 16532 22428 16584
rect 24216 16736 24268 16788
rect 22560 16668 22612 16720
rect 23756 16668 23808 16720
rect 23204 16600 23256 16652
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 23388 16532 23440 16584
rect 26976 16643 27028 16652
rect 26976 16609 26985 16643
rect 26985 16609 27019 16643
rect 27019 16609 27028 16643
rect 26976 16600 27028 16609
rect 24308 16532 24360 16584
rect 24584 16575 24636 16584
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 25136 16532 25188 16584
rect 24860 16507 24912 16516
rect 24860 16473 24894 16507
rect 24894 16473 24912 16507
rect 24860 16464 24912 16473
rect 26240 16464 26292 16516
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 22836 16439 22888 16448
rect 22836 16405 22845 16439
rect 22845 16405 22879 16439
rect 22879 16405 22888 16439
rect 22836 16396 22888 16405
rect 23296 16396 23348 16448
rect 27068 16396 27120 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 1860 16192 1912 16244
rect 5816 16192 5868 16244
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 2780 16056 2832 16108
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 5080 16099 5132 16108
rect 5080 16065 5089 16099
rect 5089 16065 5123 16099
rect 5123 16065 5132 16099
rect 5080 16056 5132 16065
rect 5448 16124 5500 16176
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6184 16124 6236 16176
rect 6092 16056 6144 16108
rect 6276 16056 6328 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7564 16124 7616 16176
rect 5540 15988 5592 16040
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7012 16056 7064 16108
rect 8208 16056 8260 16108
rect 8116 16031 8168 16040
rect 8116 15997 8125 16031
rect 8125 15997 8159 16031
rect 8159 15997 8168 16031
rect 8116 15988 8168 15997
rect 2780 15920 2832 15972
rect 3148 15920 3200 15972
rect 5632 15920 5684 15972
rect 6184 15920 6236 15972
rect 9680 16192 9732 16244
rect 10324 16192 10376 16244
rect 10692 16192 10744 16244
rect 8852 16124 8904 16176
rect 11980 16192 12032 16244
rect 8760 16056 8812 16108
rect 9036 16056 9088 16108
rect 9772 16056 9824 16108
rect 10048 16056 10100 16108
rect 9312 15988 9364 16040
rect 10232 16056 10284 16108
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 9220 15920 9272 15972
rect 10416 15920 10468 15972
rect 11336 16056 11388 16108
rect 5724 15852 5776 15904
rect 6552 15852 6604 15904
rect 6828 15852 6880 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 8852 15852 8904 15904
rect 10232 15852 10284 15904
rect 12348 16124 12400 16176
rect 14740 16192 14792 16244
rect 13728 16124 13780 16176
rect 14556 16124 14608 16176
rect 17960 16192 18012 16244
rect 18604 16192 18656 16244
rect 19524 16192 19576 16244
rect 22376 16192 22428 16244
rect 22468 16192 22520 16244
rect 26332 16192 26384 16244
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15384 16056 15436 16108
rect 18144 16124 18196 16176
rect 19064 16124 19116 16176
rect 19340 16167 19392 16176
rect 19340 16133 19350 16167
rect 19350 16133 19384 16167
rect 19384 16133 19392 16167
rect 19340 16124 19392 16133
rect 19984 16124 20036 16176
rect 17776 16056 17828 16108
rect 17224 15988 17276 16040
rect 18696 16056 18748 16108
rect 19156 16089 19208 16108
rect 19156 16056 19166 16089
rect 19166 16056 19200 16089
rect 19200 16056 19208 16089
rect 19616 16099 19668 16108
rect 19616 16065 19625 16099
rect 19625 16065 19659 16099
rect 19659 16065 19668 16099
rect 19616 16056 19668 16065
rect 20168 16124 20220 16176
rect 20904 16167 20956 16176
rect 20904 16133 20913 16167
rect 20913 16133 20947 16167
rect 20947 16133 20956 16167
rect 20904 16124 20956 16133
rect 20996 16124 21048 16176
rect 21364 16056 21416 16108
rect 21640 16056 21692 16108
rect 21088 15988 21140 16040
rect 23480 16056 23532 16108
rect 25596 16124 25648 16176
rect 24584 16056 24636 16108
rect 25872 16056 25924 16108
rect 26976 16056 27028 16108
rect 23020 15988 23072 16040
rect 24768 15988 24820 16040
rect 25136 15988 25188 16040
rect 19340 15920 19392 15972
rect 12624 15852 12676 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 15752 15852 15804 15904
rect 17776 15852 17828 15904
rect 18144 15852 18196 15904
rect 20168 15852 20220 15904
rect 20352 15852 20404 15904
rect 20628 15852 20680 15904
rect 20996 15852 21048 15904
rect 21180 15852 21232 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 23020 15852 23072 15904
rect 23940 15852 23992 15904
rect 24584 15852 24636 15904
rect 26608 15895 26660 15904
rect 26608 15861 26617 15895
rect 26617 15861 26651 15895
rect 26651 15861 26660 15895
rect 26608 15852 26660 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1768 15648 1820 15700
rect 3976 15648 4028 15700
rect 4896 15648 4948 15700
rect 6552 15648 6604 15700
rect 6828 15648 6880 15700
rect 7104 15580 7156 15632
rect 8392 15648 8444 15700
rect 8484 15648 8536 15700
rect 9220 15648 9272 15700
rect 10048 15648 10100 15700
rect 10140 15691 10192 15700
rect 10140 15657 10149 15691
rect 10149 15657 10183 15691
rect 10183 15657 10192 15691
rect 10140 15648 10192 15657
rect 5632 15512 5684 15564
rect 5724 15555 5776 15564
rect 5724 15521 5733 15555
rect 5733 15521 5767 15555
rect 5767 15521 5776 15555
rect 5724 15512 5776 15521
rect 2412 15444 2464 15496
rect 2964 15308 3016 15360
rect 3976 15419 4028 15428
rect 3976 15385 3985 15419
rect 3985 15385 4019 15419
rect 4019 15385 4028 15419
rect 3976 15376 4028 15385
rect 5080 15444 5132 15496
rect 6092 15444 6144 15496
rect 7472 15512 7524 15564
rect 6828 15487 6880 15496
rect 6828 15453 6837 15487
rect 6837 15453 6871 15487
rect 6871 15453 6880 15487
rect 6828 15444 6880 15453
rect 15844 15648 15896 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 17500 15648 17552 15700
rect 13360 15580 13412 15632
rect 14372 15623 14424 15632
rect 14372 15589 14381 15623
rect 14381 15589 14415 15623
rect 14415 15589 14424 15623
rect 14372 15580 14424 15589
rect 16672 15580 16724 15632
rect 20628 15648 20680 15700
rect 20720 15648 20772 15700
rect 22376 15691 22428 15700
rect 22376 15657 22385 15691
rect 22385 15657 22419 15691
rect 22419 15657 22428 15691
rect 22376 15648 22428 15657
rect 8300 15444 8352 15496
rect 9036 15444 9088 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10324 15555 10376 15564
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 10508 15512 10560 15564
rect 5816 15308 5868 15360
rect 6000 15308 6052 15360
rect 8116 15308 8168 15360
rect 10232 15376 10284 15428
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10876 15444 10928 15496
rect 12348 15512 12400 15564
rect 11612 15487 11664 15496
rect 11612 15453 11635 15487
rect 11635 15453 11664 15487
rect 11060 15376 11112 15428
rect 11612 15444 11664 15453
rect 14188 15444 14240 15496
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16304 15444 16356 15496
rect 16856 15487 16908 15496
rect 16856 15453 16865 15487
rect 16865 15453 16899 15487
rect 16899 15453 16908 15487
rect 16856 15444 16908 15453
rect 17408 15512 17460 15564
rect 17316 15444 17368 15496
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 18236 15512 18288 15564
rect 18972 15512 19024 15564
rect 20720 15512 20772 15564
rect 11980 15376 12032 15428
rect 14280 15376 14332 15428
rect 20260 15444 20312 15496
rect 21088 15444 21140 15496
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 22928 15512 22980 15564
rect 26424 15648 26476 15700
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 10508 15308 10560 15360
rect 11704 15308 11756 15360
rect 14004 15308 14056 15360
rect 14556 15308 14608 15360
rect 16120 15308 16172 15360
rect 17868 15308 17920 15360
rect 18236 15308 18288 15360
rect 18328 15351 18380 15360
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 19616 15308 19668 15360
rect 19800 15376 19852 15428
rect 20720 15376 20772 15428
rect 20904 15308 20956 15360
rect 21732 15419 21784 15428
rect 21732 15385 21767 15419
rect 21767 15385 21784 15419
rect 21732 15376 21784 15385
rect 22376 15444 22428 15496
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 22744 15419 22796 15428
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 23204 15376 23256 15428
rect 23388 15376 23440 15428
rect 23480 15376 23532 15428
rect 24400 15376 24452 15428
rect 25780 15444 25832 15496
rect 26332 15444 26384 15496
rect 24860 15419 24912 15428
rect 24860 15385 24894 15419
rect 24894 15385 24912 15419
rect 24860 15376 24912 15385
rect 22284 15308 22336 15360
rect 26148 15376 26200 15428
rect 26608 15376 26660 15428
rect 25596 15308 25648 15360
rect 27436 15308 27488 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 1860 15104 1912 15156
rect 2412 15104 2464 15156
rect 6644 15104 6696 15156
rect 7288 15104 7340 15156
rect 1768 15036 1820 15088
rect 3792 15036 3844 15088
rect 6368 15036 6420 15088
rect 7104 15036 7156 15088
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 4988 14968 5040 15020
rect 5264 14968 5316 15020
rect 7840 14968 7892 15020
rect 5356 14900 5408 14952
rect 6184 14900 6236 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 5724 14832 5776 14884
rect 8576 14968 8628 15020
rect 1768 14764 1820 14816
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 2412 14807 2464 14816
rect 2412 14773 2421 14807
rect 2421 14773 2455 14807
rect 2455 14773 2464 14807
rect 2412 14764 2464 14773
rect 2596 14764 2648 14816
rect 4896 14764 4948 14816
rect 6736 14764 6788 14816
rect 8024 14764 8076 14816
rect 8576 14764 8628 14816
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10048 14968 10100 15020
rect 9220 14832 9272 14884
rect 9864 14832 9916 14884
rect 10232 14832 10284 14884
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 16120 15104 16172 15156
rect 21364 15104 21416 15156
rect 22560 15147 22612 15156
rect 22560 15113 22585 15147
rect 22585 15113 22612 15147
rect 22560 15104 22612 15113
rect 13084 15036 13136 15088
rect 15752 15036 15804 15088
rect 16580 15036 16632 15088
rect 16764 15036 16816 15088
rect 19248 15036 19300 15088
rect 10416 15011 10468 15020
rect 10416 14977 10425 15011
rect 10425 14977 10459 15011
rect 10459 14977 10468 15011
rect 10416 14968 10468 14977
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 10784 14968 10836 15020
rect 11152 14968 11204 15020
rect 12164 14968 12216 15020
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 15568 14968 15620 15020
rect 16672 14968 16724 15020
rect 19892 15036 19944 15088
rect 20076 15079 20128 15088
rect 20076 15045 20110 15079
rect 20110 15045 20128 15079
rect 20076 15036 20128 15045
rect 20628 15036 20680 15088
rect 24308 15104 24360 15156
rect 24952 15036 25004 15088
rect 26516 15036 26568 15088
rect 16764 14900 16816 14952
rect 17684 14943 17736 14952
rect 17684 14909 17693 14943
rect 17693 14909 17727 14943
rect 17727 14909 17736 14943
rect 17684 14900 17736 14909
rect 19524 14900 19576 14952
rect 22008 14968 22060 15020
rect 23480 14968 23532 15020
rect 23572 15011 23624 15020
rect 23572 14977 23581 15011
rect 23581 14977 23615 15011
rect 23615 14977 23624 15011
rect 23572 14968 23624 14977
rect 23756 15011 23808 15020
rect 23756 14977 23763 15011
rect 23763 14977 23808 15011
rect 23756 14968 23808 14977
rect 24124 14968 24176 15020
rect 24400 14968 24452 15020
rect 26332 14968 26384 15020
rect 22100 14900 22152 14952
rect 22560 14900 22612 14952
rect 23204 14900 23256 14952
rect 13636 14832 13688 14884
rect 10508 14764 10560 14816
rect 13912 14764 13964 14816
rect 16948 14764 17000 14816
rect 18972 14832 19024 14884
rect 21640 14832 21692 14884
rect 17960 14764 18012 14816
rect 20904 14764 20956 14816
rect 21180 14807 21232 14816
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 22652 14764 22704 14816
rect 22744 14807 22796 14816
rect 22744 14773 22753 14807
rect 22753 14773 22787 14807
rect 22787 14773 22796 14807
rect 22744 14764 22796 14773
rect 26792 14764 26844 14816
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2964 14560 3016 14612
rect 5448 14560 5500 14612
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 10416 14560 10468 14612
rect 10600 14560 10652 14612
rect 4896 14492 4948 14544
rect 5632 14492 5684 14544
rect 7380 14492 7432 14544
rect 7656 14492 7708 14544
rect 572 14356 624 14408
rect 1860 14356 1912 14408
rect 4988 14424 5040 14476
rect 5356 14356 5408 14408
rect 5632 14356 5684 14408
rect 6736 14424 6788 14476
rect 6828 14424 6880 14476
rect 3976 14288 4028 14340
rect 5540 14288 5592 14340
rect 7012 14356 7064 14408
rect 7288 14424 7340 14476
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7656 14356 7708 14408
rect 11060 14492 11112 14544
rect 16580 14560 16632 14612
rect 17776 14603 17828 14612
rect 17776 14569 17785 14603
rect 17785 14569 17819 14603
rect 17819 14569 17828 14603
rect 17776 14560 17828 14569
rect 21272 14560 21324 14612
rect 21456 14560 21508 14612
rect 22376 14560 22428 14612
rect 11888 14492 11940 14544
rect 13820 14492 13872 14544
rect 18052 14492 18104 14544
rect 18880 14492 18932 14544
rect 19708 14535 19760 14544
rect 19708 14501 19717 14535
rect 19717 14501 19751 14535
rect 19751 14501 19760 14535
rect 19708 14492 19760 14501
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 6368 14288 6420 14340
rect 3240 14220 3292 14272
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 6000 14220 6052 14272
rect 6828 14220 6880 14272
rect 9036 14356 9088 14408
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 9680 14288 9732 14340
rect 10784 14288 10836 14340
rect 11244 14399 11296 14408
rect 11244 14365 11251 14399
rect 11251 14365 11296 14399
rect 11244 14356 11296 14365
rect 14280 14424 14332 14476
rect 14372 14424 14424 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 16764 14424 16816 14476
rect 21272 14424 21324 14476
rect 22284 14424 22336 14476
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 16672 14356 16724 14408
rect 17408 14356 17460 14408
rect 19708 14356 19760 14408
rect 21180 14356 21232 14408
rect 9588 14220 9640 14272
rect 10508 14220 10560 14272
rect 11612 14220 11664 14272
rect 14188 14288 14240 14340
rect 14372 14288 14424 14340
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 13820 14220 13872 14272
rect 14556 14220 14608 14272
rect 15936 14288 15988 14340
rect 20536 14288 20588 14340
rect 21088 14288 21140 14340
rect 22100 14356 22152 14408
rect 16764 14220 16816 14272
rect 17040 14220 17092 14272
rect 18052 14263 18104 14272
rect 18052 14229 18061 14263
rect 18061 14229 18095 14263
rect 18095 14229 18104 14263
rect 18052 14220 18104 14229
rect 18328 14220 18380 14272
rect 20996 14220 21048 14272
rect 23204 14356 23256 14408
rect 24124 14356 24176 14408
rect 24400 14356 24452 14408
rect 26516 14424 26568 14476
rect 26976 14467 27028 14476
rect 26976 14433 26985 14467
rect 26985 14433 27019 14467
rect 27019 14433 27028 14467
rect 26976 14424 27028 14433
rect 25228 14356 25280 14408
rect 22652 14331 22704 14340
rect 22652 14297 22686 14331
rect 22686 14297 22704 14331
rect 22652 14288 22704 14297
rect 23296 14288 23348 14340
rect 24308 14288 24360 14340
rect 26056 14288 26108 14340
rect 27068 14288 27120 14340
rect 23664 14220 23716 14272
rect 24400 14220 24452 14272
rect 28356 14263 28408 14272
rect 28356 14229 28365 14263
rect 28365 14229 28399 14263
rect 28399 14229 28408 14263
rect 28356 14220 28408 14229
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 5264 14016 5316 14068
rect 5908 14016 5960 14068
rect 4528 13948 4580 14000
rect 8300 14016 8352 14068
rect 11796 14016 11848 14068
rect 12348 14016 12400 14068
rect 12808 14016 12860 14068
rect 13452 14016 13504 14068
rect 13636 14016 13688 14068
rect 14556 14016 14608 14068
rect 2412 13880 2464 13932
rect 4068 13880 4120 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 8392 13991 8444 14000
rect 8392 13957 8401 13991
rect 8401 13957 8435 13991
rect 8435 13957 8444 13991
rect 8392 13948 8444 13957
rect 11888 13948 11940 14000
rect 13544 13991 13596 14000
rect 13544 13957 13553 13991
rect 13553 13957 13587 13991
rect 13587 13957 13596 13991
rect 13544 13948 13596 13957
rect 7748 13880 7800 13932
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 8484 13880 8536 13932
rect 8944 13880 8996 13932
rect 9036 13880 9088 13932
rect 10784 13880 10836 13932
rect 11612 13880 11664 13932
rect 12440 13880 12492 13932
rect 14280 13880 14332 13932
rect 14832 13948 14884 14000
rect 15752 13948 15804 14000
rect 16764 14016 16816 14068
rect 16948 14016 17000 14068
rect 18328 14016 18380 14068
rect 18512 14016 18564 14068
rect 19340 14016 19392 14068
rect 20352 14016 20404 14068
rect 17960 13948 18012 14000
rect 4252 13812 4304 13864
rect 5264 13812 5316 13864
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 6552 13812 6604 13864
rect 5448 13744 5500 13796
rect 5816 13787 5868 13796
rect 5816 13753 5825 13787
rect 5825 13753 5859 13787
rect 5859 13753 5868 13787
rect 5816 13744 5868 13753
rect 6736 13744 6788 13796
rect 9496 13812 9548 13864
rect 11152 13812 11204 13864
rect 13544 13812 13596 13864
rect 13268 13744 13320 13796
rect 14280 13744 14332 13796
rect 4988 13676 5040 13728
rect 5264 13676 5316 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 16304 13880 16356 13932
rect 18328 13923 18380 13932
rect 18328 13889 18337 13923
rect 18337 13889 18371 13923
rect 18371 13889 18380 13923
rect 18328 13880 18380 13889
rect 18696 13880 18748 13932
rect 19524 13948 19576 14000
rect 18880 13880 18932 13932
rect 20260 13880 20312 13932
rect 20628 13923 20680 13932
rect 20628 13889 20637 13923
rect 20637 13889 20671 13923
rect 20671 13889 20680 13923
rect 20628 13880 20680 13889
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 14832 13855 14884 13864
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 15016 13744 15068 13796
rect 19892 13812 19944 13864
rect 22376 14059 22428 14068
rect 22376 14025 22385 14059
rect 22385 14025 22419 14059
rect 22419 14025 22428 14059
rect 22376 14016 22428 14025
rect 22836 14016 22888 14068
rect 24860 14016 24912 14068
rect 25780 14016 25832 14068
rect 26700 14016 26752 14068
rect 22468 13948 22520 14000
rect 23296 13991 23348 14000
rect 23296 13957 23305 13991
rect 23305 13957 23339 13991
rect 23339 13957 23348 13991
rect 23296 13948 23348 13957
rect 26148 13991 26200 14000
rect 26148 13957 26157 13991
rect 26157 13957 26191 13991
rect 26191 13957 26200 13991
rect 26148 13948 26200 13957
rect 26240 13991 26292 14000
rect 26240 13957 26249 13991
rect 26249 13957 26283 13991
rect 26283 13957 26292 13991
rect 26240 13948 26292 13957
rect 17224 13744 17276 13796
rect 17776 13744 17828 13796
rect 18512 13744 18564 13796
rect 20996 13744 21048 13796
rect 21456 13812 21508 13864
rect 23664 13880 23716 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24216 13880 24268 13932
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 27528 13812 27580 13864
rect 15568 13676 15620 13728
rect 16396 13676 16448 13728
rect 17316 13676 17368 13728
rect 19524 13676 19576 13728
rect 20076 13676 20128 13728
rect 20904 13676 20956 13728
rect 21364 13676 21416 13728
rect 23388 13676 23440 13728
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 23756 13676 23808 13728
rect 24032 13676 24084 13728
rect 27068 13744 27120 13796
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 5724 13472 5776 13524
rect 6828 13472 6880 13524
rect 7380 13472 7432 13524
rect 8668 13472 8720 13524
rect 9588 13472 9640 13524
rect 10692 13472 10744 13524
rect 10876 13472 10928 13524
rect 9220 13404 9272 13456
rect 11244 13404 11296 13456
rect 4804 13336 4856 13388
rect 5724 13336 5776 13388
rect 3240 13268 3292 13320
rect 4528 13268 4580 13320
rect 4988 13268 5040 13320
rect 5448 13268 5500 13320
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 4252 13132 4304 13184
rect 5264 13132 5316 13184
rect 5816 13132 5868 13184
rect 6460 13268 6512 13320
rect 7288 13336 7340 13388
rect 14096 13472 14148 13524
rect 16120 13472 16172 13524
rect 16856 13472 16908 13524
rect 17592 13472 17644 13524
rect 18512 13472 18564 13524
rect 23572 13472 23624 13524
rect 23664 13515 23716 13524
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 26240 13472 26292 13524
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 7196 13268 7248 13320
rect 7564 13268 7616 13320
rect 8484 13268 8536 13320
rect 9312 13200 9364 13252
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9772 13268 9824 13320
rect 11244 13268 11296 13320
rect 12900 13404 12952 13456
rect 13268 13336 13320 13388
rect 13728 13404 13780 13456
rect 13820 13404 13872 13456
rect 14648 13404 14700 13456
rect 17960 13404 18012 13456
rect 20076 13404 20128 13456
rect 22744 13404 22796 13456
rect 20260 13336 20312 13388
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 8576 13132 8628 13184
rect 9634 13132 9686 13184
rect 10508 13200 10560 13252
rect 14188 13268 14240 13320
rect 14832 13268 14884 13320
rect 15752 13268 15804 13320
rect 16856 13268 16908 13320
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 18144 13268 18196 13320
rect 19064 13268 19116 13320
rect 20352 13268 20404 13320
rect 22008 13268 22060 13320
rect 23572 13311 23624 13320
rect 23572 13277 23581 13311
rect 23581 13277 23615 13311
rect 23615 13277 23624 13311
rect 23572 13268 23624 13277
rect 23664 13268 23716 13320
rect 10876 13132 10928 13184
rect 11612 13175 11664 13184
rect 11612 13141 11621 13175
rect 11621 13141 11655 13175
rect 11655 13141 11664 13175
rect 11612 13132 11664 13141
rect 13360 13132 13412 13184
rect 14740 13200 14792 13252
rect 15568 13200 15620 13252
rect 16488 13200 16540 13252
rect 14464 13175 14516 13184
rect 14464 13141 14489 13175
rect 14489 13141 14516 13175
rect 14464 13132 14516 13141
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 15016 13132 15068 13184
rect 16028 13132 16080 13184
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 18512 13132 18564 13184
rect 19248 13132 19300 13184
rect 20812 13200 20864 13252
rect 24492 13268 24544 13320
rect 26424 13336 26476 13388
rect 24124 13200 24176 13252
rect 24768 13200 24820 13252
rect 24952 13243 25004 13252
rect 24952 13209 24986 13243
rect 24986 13209 25004 13243
rect 24952 13200 25004 13209
rect 25044 13200 25096 13252
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 22744 13132 22796 13184
rect 22836 13132 22888 13184
rect 25872 13132 25924 13184
rect 26608 13200 26660 13252
rect 27804 13200 27856 13252
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 5540 12928 5592 12980
rect 6092 12928 6144 12980
rect 4528 12860 4580 12912
rect 5080 12860 5132 12912
rect 7656 12928 7708 12980
rect 9220 12928 9272 12980
rect 12164 12928 12216 12980
rect 13820 12928 13872 12980
rect 4252 12724 4304 12776
rect 6092 12792 6144 12844
rect 6276 12792 6328 12844
rect 6552 12792 6604 12844
rect 8668 12860 8720 12912
rect 10968 12860 11020 12912
rect 12716 12860 12768 12912
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 5724 12724 5776 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 8300 12724 8352 12776
rect 8484 12724 8536 12776
rect 6920 12656 6972 12708
rect 8392 12656 8444 12708
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9588 12792 9640 12844
rect 11612 12792 11664 12844
rect 12808 12792 12860 12844
rect 13360 12792 13412 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 9864 12724 9916 12776
rect 10140 12656 10192 12708
rect 12624 12656 12676 12708
rect 14096 12724 14148 12776
rect 16488 12928 16540 12980
rect 17592 12928 17644 12980
rect 18696 12928 18748 12980
rect 19248 12928 19300 12980
rect 21088 12928 21140 12980
rect 16212 12860 16264 12912
rect 17776 12903 17828 12912
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 15844 12835 15896 12844
rect 15844 12801 15851 12835
rect 15851 12801 15896 12835
rect 15844 12792 15896 12801
rect 13452 12656 13504 12708
rect 16120 12835 16172 12844
rect 16120 12801 16134 12835
rect 16134 12801 16168 12835
rect 16168 12801 16172 12835
rect 16120 12792 16172 12801
rect 16304 12792 16356 12844
rect 17776 12869 17785 12903
rect 17785 12869 17819 12903
rect 17819 12869 17828 12903
rect 17776 12860 17828 12869
rect 18328 12860 18380 12912
rect 19156 12860 19208 12912
rect 19432 12903 19484 12912
rect 19432 12869 19441 12903
rect 19441 12869 19475 12903
rect 19475 12869 19484 12903
rect 19432 12860 19484 12869
rect 16856 12767 16908 12776
rect 16856 12733 16865 12767
rect 16865 12733 16899 12767
rect 16899 12733 16908 12767
rect 16856 12724 16908 12733
rect 20628 12860 20680 12912
rect 17868 12724 17920 12776
rect 5172 12588 5224 12640
rect 6552 12588 6604 12640
rect 7196 12588 7248 12640
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 11888 12588 11940 12640
rect 13636 12588 13688 12640
rect 13728 12588 13780 12640
rect 17684 12656 17736 12708
rect 19156 12656 19208 12708
rect 19892 12792 19944 12844
rect 25136 12928 25188 12980
rect 24676 12860 24728 12912
rect 22376 12835 22428 12844
rect 22376 12801 22386 12835
rect 22386 12801 22420 12835
rect 22420 12801 22428 12835
rect 22376 12792 22428 12801
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 22744 12835 22796 12844
rect 22744 12801 22758 12835
rect 22758 12801 22792 12835
rect 22792 12801 22796 12835
rect 22744 12792 22796 12801
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 16304 12631 16356 12640
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 17592 12588 17644 12640
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 18052 12588 18104 12640
rect 18328 12588 18380 12640
rect 19432 12588 19484 12640
rect 23664 12724 23716 12776
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 24860 12792 24912 12844
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 24584 12656 24636 12708
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 22284 12588 22336 12640
rect 23480 12588 23532 12640
rect 26884 12792 26936 12844
rect 26148 12631 26200 12640
rect 26148 12597 26157 12631
rect 26157 12597 26191 12631
rect 26191 12597 26200 12631
rect 26148 12588 26200 12597
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 4252 12384 4304 12436
rect 4804 12316 4856 12368
rect 5172 12316 5224 12368
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 6000 12384 6052 12436
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 6552 12384 6604 12436
rect 7104 12384 7156 12436
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 10324 12384 10376 12436
rect 10968 12384 11020 12436
rect 11612 12384 11664 12436
rect 10876 12316 10928 12368
rect 11244 12316 11296 12368
rect 11980 12316 12032 12368
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 756 12180 808 12232
rect 3976 12180 4028 12232
rect 4252 12180 4304 12232
rect 4988 12248 5040 12300
rect 4712 12180 4764 12232
rect 5356 12180 5408 12232
rect 6644 12223 6696 12232
rect 5080 12112 5132 12164
rect 5448 12112 5500 12164
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7288 12248 7340 12300
rect 8392 12248 8444 12300
rect 9312 12248 9364 12300
rect 10692 12248 10744 12300
rect 14096 12384 14148 12436
rect 16396 12384 16448 12436
rect 16764 12384 16816 12436
rect 16948 12384 17000 12436
rect 17132 12427 17184 12436
rect 17132 12393 17141 12427
rect 17141 12393 17175 12427
rect 17175 12393 17184 12427
rect 17132 12384 17184 12393
rect 20260 12384 20312 12436
rect 16672 12316 16724 12368
rect 17500 12316 17552 12368
rect 17868 12316 17920 12368
rect 6460 12112 6512 12164
rect 7104 12180 7156 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 8668 12180 8720 12232
rect 9772 12180 9824 12232
rect 10416 12180 10468 12232
rect 11152 12180 11204 12232
rect 11704 12180 11756 12232
rect 6092 12044 6144 12096
rect 9864 12112 9916 12164
rect 9956 12112 10008 12164
rect 16212 12248 16264 12300
rect 19248 12248 19300 12300
rect 21180 12384 21232 12436
rect 21548 12384 21600 12436
rect 23388 12384 23440 12436
rect 23480 12427 23532 12436
rect 23480 12393 23489 12427
rect 23489 12393 23523 12427
rect 23523 12393 23532 12427
rect 23480 12384 23532 12393
rect 23572 12384 23624 12436
rect 25412 12384 25464 12436
rect 27344 12384 27396 12436
rect 22468 12316 22520 12368
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 17132 12180 17184 12232
rect 17408 12180 17460 12232
rect 17684 12180 17736 12232
rect 16488 12112 16540 12164
rect 16948 12112 17000 12164
rect 17592 12112 17644 12164
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 18604 12112 18656 12164
rect 19524 12112 19576 12164
rect 20996 12180 21048 12232
rect 21180 12180 21232 12232
rect 20168 12112 20220 12164
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 22652 12223 22704 12232
rect 22652 12189 22666 12223
rect 22666 12189 22700 12223
rect 22700 12189 22704 12223
rect 22652 12180 22704 12189
rect 7104 12044 7156 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 10324 12044 10376 12096
rect 11152 12044 11204 12096
rect 11980 12044 12032 12096
rect 15292 12044 15344 12096
rect 16672 12044 16724 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 18696 12044 18748 12096
rect 22284 12044 22336 12096
rect 23020 12112 23072 12164
rect 23296 12155 23348 12164
rect 23296 12121 23305 12155
rect 23305 12121 23339 12155
rect 23339 12121 23348 12155
rect 23296 12112 23348 12121
rect 24768 12180 24820 12232
rect 28356 12180 28408 12232
rect 25412 12155 25464 12164
rect 25412 12121 25446 12155
rect 25446 12121 25464 12155
rect 25412 12112 25464 12121
rect 25504 12112 25556 12164
rect 25596 12044 25648 12096
rect 26516 12087 26568 12096
rect 26516 12053 26525 12087
rect 26525 12053 26559 12087
rect 26559 12053 26568 12087
rect 26516 12044 26568 12053
rect 26608 12044 26660 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 1768 11568 1820 11620
rect 4344 11772 4396 11824
rect 5448 11704 5500 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6184 11840 6236 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 10140 11840 10192 11892
rect 11704 11840 11756 11892
rect 6460 11772 6512 11824
rect 6736 11815 6788 11824
rect 6736 11781 6745 11815
rect 6745 11781 6779 11815
rect 6779 11781 6788 11815
rect 6736 11772 6788 11781
rect 14188 11840 14240 11892
rect 14740 11840 14792 11892
rect 19432 11840 19484 11892
rect 7564 11704 7616 11756
rect 4252 11636 4304 11688
rect 4896 11636 4948 11688
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 5264 11679 5316 11688
rect 5264 11645 5273 11679
rect 5273 11645 5307 11679
rect 5307 11645 5316 11679
rect 5264 11636 5316 11645
rect 9404 11704 9456 11756
rect 10324 11704 10376 11756
rect 11796 11704 11848 11756
rect 14096 11704 14148 11756
rect 15200 11815 15252 11824
rect 15200 11781 15209 11815
rect 15209 11781 15243 11815
rect 15243 11781 15252 11815
rect 15200 11772 15252 11781
rect 16212 11772 16264 11824
rect 4712 11568 4764 11620
rect 5724 11568 5776 11620
rect 6552 11568 6604 11620
rect 3424 11500 3476 11552
rect 3976 11500 4028 11552
rect 4896 11500 4948 11552
rect 7564 11500 7616 11552
rect 10692 11636 10744 11688
rect 13912 11636 13964 11688
rect 14832 11704 14884 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15660 11704 15712 11756
rect 18972 11772 19024 11824
rect 19064 11772 19116 11824
rect 19708 11772 19760 11824
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 17500 11704 17552 11756
rect 17960 11747 18012 11756
rect 17960 11713 17994 11747
rect 17994 11713 18012 11747
rect 17960 11704 18012 11713
rect 15936 11636 15988 11688
rect 16488 11636 16540 11688
rect 9220 11500 9272 11552
rect 9864 11500 9916 11552
rect 10784 11500 10836 11552
rect 11244 11500 11296 11552
rect 12808 11500 12860 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 14924 11568 14976 11620
rect 17132 11568 17184 11620
rect 19616 11747 19668 11756
rect 19616 11713 19626 11747
rect 19626 11713 19660 11747
rect 19660 11713 19668 11747
rect 21088 11840 21140 11892
rect 22652 11840 22704 11892
rect 23020 11840 23072 11892
rect 23572 11840 23624 11892
rect 24216 11840 24268 11892
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 19616 11704 19668 11713
rect 20536 11772 20588 11824
rect 20260 11704 20312 11756
rect 21456 11704 21508 11756
rect 20168 11636 20220 11688
rect 20352 11636 20404 11688
rect 22560 11772 22612 11824
rect 22744 11772 22796 11824
rect 22192 11704 22244 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23572 11704 23624 11756
rect 23756 11772 23808 11824
rect 26608 11840 26660 11892
rect 27160 11840 27212 11892
rect 25596 11772 25648 11824
rect 26792 11772 26844 11824
rect 26884 11772 26936 11824
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 22100 11636 22152 11688
rect 23664 11679 23716 11688
rect 23664 11645 23673 11679
rect 23673 11645 23707 11679
rect 23707 11645 23716 11679
rect 23664 11636 23716 11645
rect 24768 11636 24820 11688
rect 26148 11704 26200 11756
rect 27252 11704 27304 11756
rect 26332 11636 26384 11688
rect 27068 11636 27120 11688
rect 27528 11747 27580 11756
rect 27528 11713 27537 11747
rect 27537 11713 27571 11747
rect 27571 11713 27580 11747
rect 27528 11704 27580 11713
rect 16948 11500 17000 11552
rect 17500 11500 17552 11552
rect 23572 11568 23624 11620
rect 17868 11500 17920 11552
rect 19708 11500 19760 11552
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 22652 11500 22704 11552
rect 23388 11500 23440 11552
rect 27712 11543 27764 11552
rect 27712 11509 27721 11543
rect 27721 11509 27755 11543
rect 27755 11509 27764 11543
rect 27712 11500 27764 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 4160 11296 4212 11348
rect 5172 11296 5224 11348
rect 5264 11296 5316 11348
rect 6368 11296 6420 11348
rect 9588 11296 9640 11348
rect 9864 11339 9916 11348
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 4344 11228 4396 11280
rect 5448 11228 5500 11280
rect 6092 11228 6144 11280
rect 7564 11228 7616 11280
rect 4160 11135 4212 11144
rect 4160 11101 4199 11135
rect 4199 11101 4212 11135
rect 4160 11092 4212 11101
rect 3516 11024 3568 11076
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5816 11024 5868 11076
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 7104 11160 7156 11212
rect 7472 11160 7524 11212
rect 9496 11228 9548 11280
rect 10692 11296 10744 11348
rect 11152 11296 11204 11348
rect 12348 11296 12400 11348
rect 13452 11296 13504 11348
rect 15200 11296 15252 11348
rect 12256 11228 12308 11280
rect 18236 11296 18288 11348
rect 20628 11296 20680 11348
rect 23020 11296 23072 11348
rect 25044 11296 25096 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 17224 11228 17276 11280
rect 18972 11228 19024 11280
rect 20076 11228 20128 11280
rect 20444 11228 20496 11280
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 8944 11092 8996 11144
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 5448 10956 5500 11008
rect 6920 11024 6972 11076
rect 7196 11024 7248 11076
rect 7288 11024 7340 11076
rect 8208 11067 8260 11076
rect 8208 11033 8217 11067
rect 8217 11033 8251 11067
rect 8251 11033 8260 11067
rect 8208 11024 8260 11033
rect 9036 11024 9088 11076
rect 14096 11092 14148 11144
rect 15292 11160 15344 11212
rect 17316 11160 17368 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 19524 11160 19576 11212
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 15384 11092 15436 11144
rect 16212 11092 16264 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17132 11092 17184 11144
rect 8576 10956 8628 11008
rect 8760 10956 8812 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 10324 10956 10376 11008
rect 10416 10956 10468 11008
rect 11152 10956 11204 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 15476 11067 15528 11076
rect 15476 11033 15485 11067
rect 15485 11033 15519 11067
rect 15519 11033 15528 11067
rect 15476 11024 15528 11033
rect 17316 11024 17368 11076
rect 17408 11024 17460 11076
rect 19892 11092 19944 11144
rect 20720 11092 20772 11144
rect 21088 11135 21140 11144
rect 21088 11101 21097 11135
rect 21097 11101 21131 11135
rect 21131 11101 21140 11135
rect 21088 11092 21140 11101
rect 22192 11228 22244 11280
rect 22560 11228 22612 11280
rect 21364 11160 21416 11212
rect 23020 11160 23072 11212
rect 23664 11228 23716 11280
rect 24860 11228 24912 11280
rect 24952 11228 25004 11280
rect 25964 11228 26016 11280
rect 27344 11271 27396 11280
rect 27344 11237 27353 11271
rect 27353 11237 27387 11271
rect 27387 11237 27396 11271
rect 27344 11228 27396 11237
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 22836 11135 22888 11144
rect 22836 11101 22843 11135
rect 22843 11101 22888 11135
rect 22836 11092 22888 11101
rect 23296 11160 23348 11212
rect 18144 11024 18196 11076
rect 18696 11024 18748 11076
rect 18880 11024 18932 11076
rect 19984 11024 20036 11076
rect 21456 11024 21508 11076
rect 22376 11024 22428 11076
rect 24032 11024 24084 11076
rect 24676 11092 24728 11144
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 25228 11160 25280 11212
rect 26056 11024 26108 11076
rect 16212 10956 16264 11008
rect 16856 10956 16908 11008
rect 17500 10956 17552 11008
rect 20076 10956 20128 11008
rect 23296 10999 23348 11008
rect 23296 10965 23305 10999
rect 23305 10965 23339 10999
rect 23339 10965 23348 10999
rect 23296 10956 23348 10965
rect 24308 10956 24360 11008
rect 24492 10956 24544 11008
rect 24952 10956 25004 11008
rect 26148 10956 26200 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 5448 10752 5500 10804
rect 5632 10752 5684 10804
rect 5908 10752 5960 10804
rect 7748 10752 7800 10804
rect 2596 10727 2648 10736
rect 2596 10693 2605 10727
rect 2605 10693 2639 10727
rect 2639 10693 2648 10727
rect 2596 10684 2648 10693
rect 7380 10684 7432 10736
rect 8484 10684 8536 10736
rect 9496 10752 9548 10804
rect 10324 10752 10376 10804
rect 11704 10752 11756 10804
rect 13912 10752 13964 10804
rect 15476 10752 15528 10804
rect 16120 10752 16172 10804
rect 16396 10752 16448 10804
rect 17776 10684 17828 10736
rect 19340 10752 19392 10804
rect 19156 10684 19208 10736
rect 19984 10684 20036 10736
rect 4252 10616 4304 10668
rect 5172 10616 5224 10668
rect 6184 10616 6236 10668
rect 6644 10616 6696 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7748 10616 7800 10668
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 3424 10548 3476 10600
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 9588 10616 9640 10668
rect 9864 10616 9916 10668
rect 10324 10616 10376 10668
rect 11612 10616 11664 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 13912 10616 13964 10668
rect 15660 10616 15712 10668
rect 15844 10616 15896 10668
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 16028 10616 16080 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 9680 10548 9732 10600
rect 14004 10548 14056 10600
rect 1584 10412 1636 10464
rect 5908 10412 5960 10464
rect 7472 10412 7524 10464
rect 14096 10480 14148 10532
rect 18880 10616 18932 10668
rect 19156 10548 19208 10600
rect 19616 10548 19668 10600
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 21364 10752 21416 10804
rect 22008 10684 22060 10736
rect 21548 10616 21600 10668
rect 22008 10548 22060 10600
rect 19524 10480 19576 10532
rect 21456 10480 21508 10532
rect 9220 10412 9272 10464
rect 10324 10412 10376 10464
rect 14188 10412 14240 10464
rect 14740 10412 14792 10464
rect 18512 10412 18564 10464
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 23848 10752 23900 10804
rect 24124 10752 24176 10804
rect 24768 10752 24820 10804
rect 25320 10752 25372 10804
rect 25872 10752 25924 10804
rect 27528 10752 27580 10804
rect 22192 10727 22244 10736
rect 22192 10693 22201 10727
rect 22201 10693 22235 10727
rect 22235 10693 22244 10727
rect 22192 10684 22244 10693
rect 22376 10684 22428 10736
rect 24400 10684 24452 10736
rect 22836 10616 22888 10668
rect 23388 10616 23440 10668
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 23664 10659 23716 10668
rect 23664 10625 23673 10659
rect 23673 10625 23707 10659
rect 23707 10625 23716 10659
rect 23664 10616 23716 10625
rect 24860 10616 24912 10668
rect 25136 10616 25188 10668
rect 25320 10616 25372 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 24952 10548 25004 10600
rect 26240 10548 26292 10600
rect 27068 10548 27120 10600
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 22652 10455 22704 10464
rect 22652 10421 22661 10455
rect 22661 10421 22695 10455
rect 22695 10421 22704 10455
rect 22652 10412 22704 10421
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 25044 10412 25096 10464
rect 25228 10412 25280 10464
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 3516 10208 3568 10260
rect 4160 10208 4212 10260
rect 4804 10208 4856 10260
rect 6644 10208 6696 10260
rect 7196 10208 7248 10260
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 10600 10251 10652 10260
rect 10600 10217 10609 10251
rect 10609 10217 10643 10251
rect 10643 10217 10652 10251
rect 10600 10208 10652 10217
rect 4068 10140 4120 10192
rect 4712 10140 4764 10192
rect 7288 10140 7340 10192
rect 8392 10140 8444 10192
rect 17316 10208 17368 10260
rect 18144 10208 18196 10260
rect 18788 10208 18840 10260
rect 20536 10208 20588 10260
rect 20996 10208 21048 10260
rect 21272 10208 21324 10260
rect 22008 10208 22060 10260
rect 23204 10208 23256 10260
rect 23388 10208 23440 10260
rect 25780 10208 25832 10260
rect 26792 10208 26844 10260
rect 13728 10140 13780 10192
rect 848 10004 900 10056
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4344 10004 4396 10056
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 5172 10072 5224 10124
rect 4896 10004 4948 10056
rect 6184 10004 6236 10056
rect 7380 10072 7432 10124
rect 6644 10004 6696 10056
rect 7104 10004 7156 10056
rect 7288 10004 7340 10056
rect 7564 10004 7616 10056
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10324 10072 10376 10124
rect 11152 10072 11204 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 9864 10047 9916 10056
rect 9864 10013 9895 10047
rect 9895 10013 9916 10047
rect 9864 10004 9916 10013
rect 5908 9936 5960 9988
rect 6460 9936 6512 9988
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 13728 10004 13780 10056
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 9680 9868 9732 9920
rect 11796 9936 11848 9988
rect 12900 9936 12952 9988
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 19340 10140 19392 10192
rect 19616 10140 19668 10192
rect 23572 10140 23624 10192
rect 24032 10140 24084 10192
rect 24676 10140 24728 10192
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 19340 10004 19392 10056
rect 19524 10047 19576 10056
rect 19524 10013 19534 10047
rect 19534 10013 19568 10047
rect 19568 10013 19576 10047
rect 19524 10004 19576 10013
rect 19892 10047 19944 10056
rect 19892 10013 19906 10047
rect 19906 10013 19940 10047
rect 19940 10013 19944 10047
rect 19892 10004 19944 10013
rect 20352 10004 20404 10056
rect 14480 9936 14532 9988
rect 14832 9936 14884 9988
rect 16764 9936 16816 9988
rect 17776 9979 17828 9988
rect 17776 9945 17785 9979
rect 17785 9945 17819 9979
rect 17819 9945 17828 9979
rect 17776 9936 17828 9945
rect 18052 9936 18104 9988
rect 19156 9868 19208 9920
rect 21088 10004 21140 10056
rect 20536 9979 20588 9988
rect 20536 9945 20545 9979
rect 20545 9945 20579 9979
rect 20579 9945 20588 9979
rect 20536 9936 20588 9945
rect 20812 9936 20864 9988
rect 19892 9868 19944 9920
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 21640 10072 21692 10124
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 22284 10004 22336 10056
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 23204 10004 23256 10056
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 24768 10004 24820 10056
rect 26884 10004 26936 10056
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 22468 9936 22520 9988
rect 23204 9868 23256 9920
rect 25872 9936 25924 9988
rect 26884 9868 26936 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 2596 9664 2648 9716
rect 4712 9664 4764 9716
rect 5080 9596 5132 9648
rect 7380 9707 7432 9716
rect 7380 9673 7405 9707
rect 7405 9673 7432 9707
rect 7380 9664 7432 9673
rect 7564 9664 7616 9716
rect 10416 9664 10468 9716
rect 10692 9664 10744 9716
rect 13912 9664 13964 9716
rect 15200 9707 15252 9716
rect 15200 9673 15209 9707
rect 15209 9673 15243 9707
rect 15243 9673 15252 9707
rect 15200 9664 15252 9673
rect 17776 9664 17828 9716
rect 19524 9664 19576 9716
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 5172 9528 5224 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 4436 9460 4488 9512
rect 4712 9503 4764 9512
rect 4712 9469 4721 9503
rect 4721 9469 4755 9503
rect 4755 9469 4764 9503
rect 4712 9460 4764 9469
rect 5080 9460 5132 9512
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 5908 9528 5960 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 7104 9596 7156 9648
rect 9220 9596 9272 9648
rect 8484 9528 8536 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 11152 9528 11204 9580
rect 11796 9528 11848 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 6644 9460 6696 9512
rect 6000 9392 6052 9444
rect 6460 9392 6512 9444
rect 8392 9460 8444 9512
rect 12532 9596 12584 9648
rect 13820 9596 13872 9648
rect 12256 9460 12308 9512
rect 7196 9324 7248 9376
rect 7748 9392 7800 9444
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 12900 9528 12952 9580
rect 13360 9528 13412 9580
rect 16028 9596 16080 9648
rect 17592 9596 17644 9648
rect 18052 9596 18104 9648
rect 18144 9596 18196 9648
rect 15476 9528 15528 9580
rect 16672 9528 16724 9580
rect 17684 9528 17736 9580
rect 19892 9639 19944 9648
rect 19892 9605 19901 9639
rect 19901 9605 19935 9639
rect 19935 9605 19944 9639
rect 19892 9596 19944 9605
rect 20260 9664 20312 9716
rect 21364 9664 21416 9716
rect 23664 9664 23716 9716
rect 17224 9460 17276 9512
rect 18512 9460 18564 9512
rect 14280 9392 14332 9444
rect 15476 9392 15528 9444
rect 16304 9392 16356 9444
rect 17960 9392 18012 9444
rect 18696 9392 18748 9444
rect 19524 9392 19576 9444
rect 19892 9460 19944 9512
rect 20444 9460 20496 9512
rect 20996 9528 21048 9580
rect 22468 9528 22520 9580
rect 23848 9596 23900 9648
rect 24124 9596 24176 9648
rect 25504 9664 25556 9716
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 23388 9528 23440 9580
rect 20812 9392 20864 9444
rect 23020 9392 23072 9444
rect 14372 9324 14424 9376
rect 15292 9324 15344 9376
rect 16672 9324 16724 9376
rect 19156 9324 19208 9376
rect 20536 9324 20588 9376
rect 22560 9324 22612 9376
rect 23112 9324 23164 9376
rect 25504 9571 25556 9580
rect 25504 9537 25513 9571
rect 25513 9537 25547 9571
rect 25547 9537 25556 9571
rect 25504 9528 25556 9537
rect 26332 9528 26384 9580
rect 25964 9460 26016 9512
rect 26056 9460 26108 9512
rect 25412 9392 25464 9444
rect 25504 9392 25556 9444
rect 27896 9392 27948 9444
rect 26516 9324 26568 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 1860 9120 1912 9172
rect 3332 9120 3384 9172
rect 4804 9120 4856 9172
rect 5816 9120 5868 9172
rect 6828 9120 6880 9172
rect 9312 9120 9364 9172
rect 9772 9120 9824 9172
rect 15200 9120 15252 9172
rect 16856 9120 16908 9172
rect 16948 9120 17000 9172
rect 18512 9120 18564 9172
rect 19248 9120 19300 9172
rect 19524 9163 19576 9172
rect 19524 9129 19533 9163
rect 19533 9129 19567 9163
rect 19567 9129 19576 9163
rect 19524 9120 19576 9129
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 5264 8984 5316 9036
rect 4804 8916 4856 8968
rect 5724 8916 5776 8968
rect 1952 8848 2004 8900
rect 5172 8848 5224 8900
rect 4896 8780 4948 8832
rect 5356 8780 5408 8832
rect 7012 9052 7064 9104
rect 11704 9052 11756 9104
rect 13452 9052 13504 9104
rect 13544 9052 13596 9104
rect 14648 9052 14700 9104
rect 15108 9052 15160 9104
rect 6644 8984 6696 9036
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7196 8984 7248 9036
rect 6368 8848 6420 8900
rect 7380 8916 7432 8968
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 8944 8916 8996 8968
rect 11888 8916 11940 8968
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 14740 8984 14792 9036
rect 14004 8916 14056 8968
rect 14556 8916 14608 8968
rect 7288 8848 7340 8900
rect 10784 8848 10836 8900
rect 12164 8848 12216 8900
rect 14464 8848 14516 8900
rect 14648 8848 14700 8900
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 16212 9095 16264 9104
rect 16212 9061 16221 9095
rect 16221 9061 16255 9095
rect 16255 9061 16264 9095
rect 16212 9052 16264 9061
rect 16304 9052 16356 9104
rect 23296 9120 23348 9172
rect 24032 9163 24084 9172
rect 24032 9129 24041 9163
rect 24041 9129 24075 9163
rect 24075 9129 24084 9163
rect 24032 9120 24084 9129
rect 25780 9120 25832 9172
rect 27252 9120 27304 9172
rect 19340 8984 19392 9036
rect 19892 9052 19944 9104
rect 20720 9052 20772 9104
rect 16488 8916 16540 8968
rect 17224 8916 17276 8968
rect 9864 8780 9916 8832
rect 11980 8780 12032 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 13452 8780 13504 8832
rect 15384 8780 15436 8832
rect 16488 8780 16540 8832
rect 17592 8848 17644 8900
rect 17500 8780 17552 8832
rect 18328 8959 18380 8968
rect 18328 8925 18338 8959
rect 18338 8925 18372 8959
rect 18372 8925 18380 8959
rect 18328 8916 18380 8925
rect 18420 8916 18472 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 18880 8916 18932 8968
rect 19248 8916 19300 8968
rect 20444 8984 20496 9036
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 20076 8916 20128 8968
rect 23388 8916 23440 8968
rect 25136 8916 25188 8968
rect 26700 8916 26752 8968
rect 26976 8916 27028 8968
rect 19432 8891 19484 8900
rect 19432 8857 19441 8891
rect 19441 8857 19475 8891
rect 19475 8857 19484 8891
rect 19432 8848 19484 8857
rect 20628 8848 20680 8900
rect 21088 8891 21140 8900
rect 21088 8857 21122 8891
rect 21122 8857 21140 8891
rect 21088 8848 21140 8857
rect 19892 8823 19944 8832
rect 19892 8789 19901 8823
rect 19901 8789 19935 8823
rect 19935 8789 19944 8823
rect 19892 8780 19944 8789
rect 20076 8780 20128 8832
rect 20260 8780 20312 8832
rect 20996 8780 21048 8832
rect 22192 8823 22244 8832
rect 22192 8789 22201 8823
rect 22201 8789 22235 8823
rect 22235 8789 22244 8823
rect 22192 8780 22244 8789
rect 23112 8848 23164 8900
rect 22836 8780 22888 8832
rect 24400 8848 24452 8900
rect 25320 8891 25372 8900
rect 25320 8857 25354 8891
rect 25354 8857 25372 8891
rect 25320 8848 25372 8857
rect 26608 8848 26660 8900
rect 27160 8891 27212 8900
rect 27160 8857 27172 8891
rect 27172 8857 27212 8891
rect 27160 8848 27212 8857
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 5448 8576 5500 8628
rect 6828 8576 6880 8628
rect 7012 8576 7064 8628
rect 7288 8576 7340 8628
rect 7748 8576 7800 8628
rect 12440 8576 12492 8628
rect 13728 8576 13780 8628
rect 5264 8440 5316 8492
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 5632 8440 5684 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6460 8440 6512 8492
rect 6000 8372 6052 8424
rect 6644 8372 6696 8424
rect 6920 8440 6972 8492
rect 10508 8508 10560 8560
rect 12164 8508 12216 8560
rect 16120 8576 16172 8628
rect 16856 8576 16908 8628
rect 17960 8576 18012 8628
rect 19340 8576 19392 8628
rect 19892 8576 19944 8628
rect 20996 8576 21048 8628
rect 22008 8576 22060 8628
rect 23572 8576 23624 8628
rect 24860 8576 24912 8628
rect 25136 8576 25188 8628
rect 25596 8576 25648 8628
rect 25872 8576 25924 8628
rect 20352 8508 20404 8560
rect 20812 8508 20864 8560
rect 24952 8508 25004 8560
rect 5540 8347 5592 8356
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 5724 8304 5776 8356
rect 6552 8304 6604 8356
rect 7748 8440 7800 8492
rect 11152 8440 11204 8492
rect 12532 8440 12584 8492
rect 12992 8440 13044 8492
rect 14004 8440 14056 8492
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18328 8483 18380 8492
rect 18328 8449 18356 8483
rect 18356 8449 18380 8483
rect 18328 8440 18380 8449
rect 18788 8440 18840 8492
rect 19340 8483 19392 8492
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 19800 8440 19852 8492
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 20628 8440 20680 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22560 8440 22612 8492
rect 25596 8440 25648 8492
rect 9220 8372 9272 8424
rect 9588 8372 9640 8424
rect 17500 8372 17552 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 6920 8236 6972 8288
rect 13452 8304 13504 8356
rect 10324 8236 10376 8288
rect 10416 8236 10468 8288
rect 13636 8236 13688 8288
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 16212 8304 16264 8356
rect 17132 8304 17184 8356
rect 17960 8304 18012 8356
rect 18880 8304 18932 8356
rect 19248 8236 19300 8288
rect 20168 8304 20220 8356
rect 24124 8347 24176 8356
rect 24124 8313 24133 8347
rect 24133 8313 24167 8347
rect 24167 8313 24176 8347
rect 24124 8304 24176 8313
rect 19892 8279 19944 8288
rect 19892 8245 19901 8279
rect 19901 8245 19935 8279
rect 19935 8245 19944 8279
rect 19892 8236 19944 8245
rect 22560 8236 22612 8288
rect 23388 8236 23440 8288
rect 27068 8236 27120 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 4988 8032 5040 8084
rect 9496 8032 9548 8084
rect 5356 7964 5408 8016
rect 11796 7964 11848 8016
rect 6736 7896 6788 7948
rect 940 7828 992 7880
rect 4344 7828 4396 7880
rect 5080 7828 5132 7880
rect 6000 7828 6052 7880
rect 6460 7828 6512 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 10692 7828 10744 7880
rect 12532 7896 12584 7948
rect 12900 7964 12952 8016
rect 12808 7871 12860 7880
rect 12808 7837 12815 7871
rect 12815 7837 12860 7871
rect 4252 7692 4304 7744
rect 5540 7692 5592 7744
rect 6552 7692 6604 7744
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 12808 7828 12860 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13360 7964 13412 8016
rect 13912 7828 13964 7880
rect 14372 7828 14424 7880
rect 15568 7828 15620 7880
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16580 7964 16632 8016
rect 19064 7964 19116 8016
rect 20812 8032 20864 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 23204 8032 23256 8084
rect 27896 8032 27948 8084
rect 20904 7964 20956 8016
rect 22100 7964 22152 8016
rect 23296 7964 23348 8016
rect 24308 7964 24360 8016
rect 18880 7896 18932 7948
rect 21548 7896 21600 7948
rect 15568 7692 15620 7744
rect 15752 7692 15804 7744
rect 17132 7760 17184 7812
rect 18236 7760 18288 7812
rect 18512 7828 18564 7880
rect 19708 7828 19760 7880
rect 19892 7828 19944 7880
rect 21824 7871 21876 7880
rect 21824 7837 21831 7871
rect 21831 7837 21876 7871
rect 21824 7828 21876 7837
rect 22100 7871 22152 7880
rect 22100 7837 22114 7871
rect 22114 7837 22148 7871
rect 22148 7837 22152 7871
rect 22100 7828 22152 7837
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 22928 7871 22980 7880
rect 22928 7837 22935 7871
rect 22935 7837 22980 7871
rect 22928 7828 22980 7837
rect 24860 7828 24912 7880
rect 25780 7828 25832 7880
rect 26700 7828 26752 7880
rect 17408 7692 17460 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 19064 7692 19116 7744
rect 20076 7803 20128 7812
rect 20076 7769 20110 7803
rect 20110 7769 20128 7803
rect 20076 7760 20128 7769
rect 20628 7760 20680 7812
rect 20352 7692 20404 7744
rect 22652 7760 22704 7812
rect 23756 7760 23808 7812
rect 26516 7760 26568 7812
rect 27344 7760 27396 7812
rect 26332 7692 26384 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 8852 7488 8904 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 3884 7352 3936 7404
rect 5724 7420 5776 7472
rect 7196 7420 7248 7472
rect 8300 7420 8352 7472
rect 9128 7420 9180 7472
rect 9404 7420 9456 7472
rect 6092 7352 6144 7404
rect 8392 7352 8444 7404
rect 7012 7284 7064 7336
rect 9680 7259 9732 7268
rect 9680 7225 9689 7259
rect 9689 7225 9723 7259
rect 9723 7225 9732 7259
rect 9680 7216 9732 7225
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 12256 7488 12308 7540
rect 13084 7420 13136 7472
rect 10784 7284 10836 7336
rect 12624 7352 12676 7404
rect 12808 7352 12860 7404
rect 13268 7420 13320 7472
rect 15384 7420 15436 7472
rect 13544 7352 13596 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 16028 7488 16080 7540
rect 17040 7488 17092 7540
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17132 7463 17184 7472
rect 17132 7429 17141 7463
rect 17141 7429 17175 7463
rect 17175 7429 17184 7463
rect 17132 7420 17184 7429
rect 18972 7420 19024 7472
rect 19892 7420 19944 7472
rect 2780 7148 2832 7200
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 4160 7148 4212 7200
rect 4804 7148 4856 7200
rect 10324 7148 10376 7200
rect 10876 7148 10928 7200
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 15292 7284 15344 7336
rect 17316 7395 17368 7404
rect 17316 7361 17330 7395
rect 17330 7361 17364 7395
rect 17364 7361 17368 7395
rect 17316 7352 17368 7361
rect 17684 7352 17736 7404
rect 18512 7352 18564 7404
rect 19984 7352 20036 7404
rect 17868 7284 17920 7336
rect 18972 7284 19024 7336
rect 19248 7284 19300 7336
rect 14096 7216 14148 7268
rect 15200 7216 15252 7268
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 14372 7148 14424 7200
rect 17960 7216 18012 7268
rect 20628 7488 20680 7540
rect 22376 7488 22428 7540
rect 24216 7488 24268 7540
rect 26608 7531 26660 7540
rect 26608 7497 26617 7531
rect 26617 7497 26651 7531
rect 26651 7497 26660 7531
rect 26608 7488 26660 7497
rect 20444 7463 20496 7472
rect 20444 7429 20453 7463
rect 20453 7429 20487 7463
rect 20487 7429 20496 7463
rect 20444 7420 20496 7429
rect 22192 7420 22244 7472
rect 20260 7352 20312 7404
rect 21640 7352 21692 7404
rect 25044 7352 25096 7404
rect 25872 7352 25924 7404
rect 20720 7284 20772 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 23572 7284 23624 7336
rect 17408 7148 17460 7200
rect 19064 7148 19116 7200
rect 24124 7216 24176 7268
rect 27160 7148 27212 7200
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 9220 6944 9272 6996
rect 10140 6944 10192 6996
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 2964 6808 3016 6860
rect 2688 6740 2740 6792
rect 6092 6808 6144 6860
rect 7656 6876 7708 6928
rect 10876 6876 10928 6928
rect 12072 6876 12124 6928
rect 13452 6944 13504 6996
rect 14280 6944 14332 6996
rect 15568 6944 15620 6996
rect 14372 6876 14424 6928
rect 16120 6876 16172 6928
rect 21732 6944 21784 6996
rect 21916 6876 21968 6928
rect 22376 6876 22428 6928
rect 23296 6876 23348 6928
rect 23940 6944 23992 6996
rect 25136 6944 25188 6996
rect 26240 6987 26292 6996
rect 26240 6953 26249 6987
rect 26249 6953 26283 6987
rect 26283 6953 26292 6987
rect 26240 6944 26292 6953
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 7012 6740 7064 6792
rect 8944 6740 8996 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 12256 6808 12308 6860
rect 5816 6672 5868 6724
rect 6276 6672 6328 6724
rect 7472 6672 7524 6724
rect 3148 6604 3200 6656
rect 4896 6604 4948 6656
rect 5356 6604 5408 6656
rect 8300 6604 8352 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 12808 6740 12860 6792
rect 16212 6808 16264 6860
rect 16672 6808 16724 6860
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 11888 6715 11940 6724
rect 11888 6681 11897 6715
rect 11897 6681 11931 6715
rect 11931 6681 11940 6715
rect 11888 6672 11940 6681
rect 12532 6672 12584 6724
rect 12716 6672 12768 6724
rect 16764 6740 16816 6792
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 17224 6808 17276 6860
rect 20168 6808 20220 6860
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 20628 6783 20680 6792
rect 20628 6749 20661 6783
rect 20661 6749 20680 6783
rect 20628 6740 20680 6749
rect 21180 6740 21232 6792
rect 21732 6808 21784 6860
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 12348 6604 12400 6656
rect 13544 6647 13596 6656
rect 13544 6613 13574 6647
rect 13574 6613 13596 6647
rect 13544 6604 13596 6613
rect 13728 6647 13780 6656
rect 13728 6613 13737 6647
rect 13737 6613 13771 6647
rect 13771 6613 13780 6647
rect 13728 6604 13780 6613
rect 15936 6604 15988 6656
rect 18696 6672 18748 6724
rect 18972 6672 19024 6724
rect 20076 6672 20128 6724
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 19892 6604 19944 6656
rect 20536 6715 20588 6724
rect 20536 6681 20545 6715
rect 20545 6681 20579 6715
rect 20579 6681 20588 6715
rect 20536 6672 20588 6681
rect 21824 6740 21876 6792
rect 22836 6740 22888 6792
rect 21916 6672 21968 6724
rect 20904 6604 20956 6656
rect 23480 6604 23532 6656
rect 24768 6740 24820 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 26332 6808 26384 6860
rect 26700 6851 26752 6860
rect 26700 6817 26709 6851
rect 26709 6817 26743 6851
rect 26743 6817 26752 6851
rect 26700 6808 26752 6817
rect 23664 6715 23716 6724
rect 23664 6681 23673 6715
rect 23673 6681 23707 6715
rect 23707 6681 23716 6715
rect 23664 6672 23716 6681
rect 26516 6740 26568 6792
rect 26240 6672 26292 6724
rect 25044 6604 25096 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 4804 6400 4856 6452
rect 5448 6400 5500 6452
rect 5908 6400 5960 6452
rect 8208 6400 8260 6452
rect 3700 6332 3752 6384
rect 3884 6332 3936 6384
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 2780 6264 2832 6316
rect 7380 6332 7432 6384
rect 7656 6332 7708 6384
rect 10600 6332 10652 6384
rect 12256 6332 12308 6384
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6460 6264 6512 6316
rect 6828 6264 6880 6316
rect 8944 6264 8996 6316
rect 9220 6264 9272 6316
rect 10416 6264 10468 6316
rect 12348 6264 12400 6316
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 14464 6332 14516 6384
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 15660 6400 15712 6452
rect 16396 6400 16448 6452
rect 17592 6400 17644 6452
rect 14556 6264 14608 6316
rect 7012 6196 7064 6248
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15292 6264 15344 6316
rect 15660 6196 15712 6248
rect 15108 6128 15160 6180
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 20904 6332 20956 6384
rect 24584 6400 24636 6452
rect 24676 6443 24728 6452
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 24768 6400 24820 6452
rect 26056 6400 26108 6452
rect 26424 6400 26476 6452
rect 17592 6307 17644 6316
rect 17592 6273 17626 6307
rect 17626 6273 17644 6307
rect 17592 6264 17644 6273
rect 18144 6264 18196 6316
rect 19248 6264 19300 6316
rect 20444 6264 20496 6316
rect 20536 6264 20588 6316
rect 23112 6332 23164 6384
rect 16212 6128 16264 6180
rect 21548 6196 21600 6248
rect 20260 6128 20312 6180
rect 22928 6128 22980 6180
rect 8300 6060 8352 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9312 6060 9364 6112
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 14004 6060 14056 6112
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 17500 6060 17552 6112
rect 19340 6060 19392 6112
rect 22284 6060 22336 6112
rect 24584 6196 24636 6248
rect 24860 6196 24912 6248
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 24584 6060 24636 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 3056 5856 3108 5908
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 3792 5856 3844 5908
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5356 5720 5408 5772
rect 7012 5856 7064 5908
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 5448 5652 5500 5704
rect 5724 5652 5776 5704
rect 8392 5856 8444 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 13544 5856 13596 5908
rect 14280 5856 14332 5908
rect 15108 5856 15160 5908
rect 15384 5856 15436 5908
rect 18696 5899 18748 5908
rect 18696 5865 18705 5899
rect 18705 5865 18739 5899
rect 18739 5865 18748 5899
rect 18696 5856 18748 5865
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 12808 5831 12860 5840
rect 12808 5797 12817 5831
rect 12817 5797 12851 5831
rect 12851 5797 12860 5831
rect 12808 5788 12860 5797
rect 13268 5788 13320 5840
rect 13912 5788 13964 5840
rect 14004 5788 14056 5840
rect 14648 5788 14700 5840
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 13728 5720 13780 5772
rect 9036 5652 9088 5704
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 5540 5584 5592 5636
rect 7104 5584 7156 5636
rect 7564 5584 7616 5636
rect 12072 5652 12124 5704
rect 2780 5516 2832 5568
rect 3884 5516 3936 5568
rect 9312 5516 9364 5568
rect 11704 5584 11756 5636
rect 12164 5584 12216 5636
rect 13176 5652 13228 5704
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 13636 5652 13688 5704
rect 13912 5652 13964 5704
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 15016 5695 15068 5704
rect 15016 5661 15023 5695
rect 15023 5661 15068 5695
rect 15016 5652 15068 5661
rect 15936 5788 15988 5840
rect 15384 5720 15436 5772
rect 18788 5720 18840 5772
rect 19248 5720 19300 5772
rect 19708 5720 19760 5772
rect 21456 5856 21508 5908
rect 22744 5856 22796 5908
rect 25596 5856 25648 5908
rect 22468 5720 22520 5772
rect 24584 5763 24636 5772
rect 24584 5729 24593 5763
rect 24593 5729 24627 5763
rect 24627 5729 24636 5763
rect 24584 5720 24636 5729
rect 15292 5695 15344 5704
rect 15292 5661 15306 5695
rect 15306 5661 15340 5695
rect 15340 5661 15344 5695
rect 15292 5652 15344 5661
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 14004 5584 14056 5636
rect 16580 5627 16632 5636
rect 16580 5593 16589 5627
rect 16589 5593 16623 5627
rect 16623 5593 16632 5627
rect 16580 5584 16632 5593
rect 17592 5627 17644 5636
rect 17592 5593 17601 5627
rect 17601 5593 17635 5627
rect 17635 5593 17644 5627
rect 17592 5584 17644 5593
rect 17684 5627 17736 5636
rect 17684 5593 17693 5627
rect 17693 5593 17727 5627
rect 17727 5593 17736 5627
rect 17684 5584 17736 5593
rect 12716 5516 12768 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 21364 5652 21416 5704
rect 21640 5652 21692 5704
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 18972 5584 19024 5636
rect 21180 5584 21232 5636
rect 16672 5516 16724 5525
rect 19616 5516 19668 5568
rect 20536 5516 20588 5568
rect 21456 5584 21508 5636
rect 26516 5652 26568 5704
rect 24032 5516 24084 5568
rect 24124 5516 24176 5568
rect 25228 5584 25280 5636
rect 26792 5584 26844 5636
rect 26516 5516 26568 5568
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 2780 5312 2832 5364
rect 3056 5312 3108 5364
rect 6276 5312 6328 5364
rect 9036 5312 9088 5364
rect 9496 5312 9548 5364
rect 12348 5312 12400 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 15200 5312 15252 5364
rect 20812 5312 20864 5364
rect 26240 5312 26292 5364
rect 5172 5244 5224 5296
rect 4068 5176 4120 5228
rect 6828 5176 6880 5228
rect 7012 5176 7064 5228
rect 8208 5219 8260 5228
rect 8208 5185 8242 5219
rect 8242 5185 8260 5219
rect 8208 5176 8260 5185
rect 9864 5176 9916 5228
rect 12072 5244 12124 5296
rect 12440 5244 12492 5296
rect 14280 5244 14332 5296
rect 15292 5244 15344 5296
rect 18236 5244 18288 5296
rect 18420 5287 18472 5296
rect 18420 5253 18454 5287
rect 18454 5253 18472 5287
rect 18420 5244 18472 5253
rect 19064 5244 19116 5296
rect 22836 5244 22888 5296
rect 24492 5244 24544 5296
rect 27804 5244 27856 5296
rect 3792 4972 3844 5024
rect 6184 5040 6236 5092
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 12624 5176 12676 5228
rect 12992 5176 13044 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 13820 5176 13872 5228
rect 15752 5176 15804 5228
rect 16672 5176 16724 5228
rect 16764 5176 16816 5228
rect 16304 5108 16356 5160
rect 25228 5219 25280 5228
rect 25228 5185 25237 5219
rect 25237 5185 25271 5219
rect 25271 5185 25280 5219
rect 25228 5176 25280 5185
rect 26424 5176 26476 5228
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 20168 5108 20220 5160
rect 24400 5108 24452 5160
rect 27160 5151 27212 5160
rect 27160 5117 27169 5151
rect 27169 5117 27203 5151
rect 27203 5117 27212 5151
rect 27160 5108 27212 5117
rect 14556 4972 14608 5024
rect 17960 5040 18012 5092
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 16396 4972 16448 5024
rect 22468 5040 22520 5092
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 7104 4768 7156 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 1584 4632 1636 4684
rect 4068 4632 4120 4684
rect 10416 4632 10468 4684
rect 12532 4768 12584 4820
rect 13268 4768 13320 4820
rect 14280 4768 14332 4820
rect 14648 4768 14700 4820
rect 14740 4700 14792 4752
rect 1492 4564 1544 4616
rect 7104 4564 7156 4616
rect 8668 4564 8720 4616
rect 9956 4564 10008 4616
rect 10876 4564 10928 4616
rect 16764 4768 16816 4820
rect 20168 4768 20220 4820
rect 21548 4768 21600 4820
rect 24032 4811 24084 4820
rect 24032 4777 24041 4811
rect 24041 4777 24075 4811
rect 24075 4777 24084 4811
rect 24032 4768 24084 4777
rect 25964 4811 26016 4820
rect 25964 4777 25973 4811
rect 25973 4777 26007 4811
rect 26007 4777 26016 4811
rect 25964 4768 26016 4777
rect 27804 4811 27856 4820
rect 27804 4777 27813 4811
rect 27813 4777 27847 4811
rect 27847 4777 27856 4811
rect 27804 4768 27856 4777
rect 16672 4700 16724 4752
rect 19524 4700 19576 4752
rect 18052 4632 18104 4684
rect 18972 4632 19024 4684
rect 4252 4496 4304 4548
rect 11060 4496 11112 4548
rect 12624 4539 12676 4548
rect 12624 4505 12658 4539
rect 12658 4505 12676 4539
rect 12624 4496 12676 4505
rect 14096 4496 14148 4548
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 15844 4607 15896 4616
rect 15844 4573 15878 4607
rect 15878 4573 15896 4607
rect 15844 4564 15896 4573
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 10508 4428 10560 4480
rect 17408 4496 17460 4548
rect 18052 4539 18104 4548
rect 18052 4505 18061 4539
rect 18061 4505 18095 4539
rect 18095 4505 18104 4539
rect 18052 4496 18104 4505
rect 18144 4496 18196 4548
rect 16764 4428 16816 4480
rect 17776 4428 17828 4480
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 19892 4607 19944 4616
rect 19892 4573 19906 4607
rect 19906 4573 19940 4607
rect 19940 4573 19944 4607
rect 19892 4564 19944 4573
rect 19708 4539 19760 4548
rect 19708 4505 19717 4539
rect 19717 4505 19751 4539
rect 19751 4505 19760 4539
rect 19708 4496 19760 4505
rect 24308 4632 24360 4684
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 22928 4607 22980 4616
rect 22928 4573 22962 4607
rect 22962 4573 22980 4607
rect 20720 4496 20772 4548
rect 22928 4564 22980 4573
rect 26424 4675 26476 4684
rect 26424 4641 26433 4675
rect 26433 4641 26467 4675
rect 26467 4641 26476 4675
rect 26424 4632 26476 4641
rect 22192 4428 22244 4480
rect 22652 4428 22704 4480
rect 26516 4564 26568 4616
rect 25596 4428 25648 4480
rect 25780 4428 25832 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 8300 4224 8352 4276
rect 15844 4224 15896 4276
rect 16948 4224 17000 4276
rect 19892 4224 19944 4276
rect 21364 4224 21416 4276
rect 1584 4088 1636 4140
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 7012 4131 7064 4140
rect 7012 4097 7046 4131
rect 7046 4097 7064 4131
rect 7012 4088 7064 4097
rect 8576 4156 8628 4208
rect 10416 4156 10468 4208
rect 13728 4199 13780 4208
rect 13728 4165 13737 4199
rect 13737 4165 13771 4199
rect 13771 4165 13780 4199
rect 13728 4156 13780 4165
rect 13912 4199 13964 4208
rect 13912 4165 13937 4199
rect 13937 4165 13964 4199
rect 13912 4156 13964 4165
rect 14648 4156 14700 4208
rect 15660 4156 15712 4208
rect 17132 4199 17184 4208
rect 17132 4165 17144 4199
rect 17144 4165 17184 4199
rect 17132 4156 17184 4165
rect 19340 4156 19392 4208
rect 20536 4156 20588 4208
rect 27160 4224 27212 4276
rect 22284 4199 22336 4208
rect 22284 4165 22293 4199
rect 22293 4165 22327 4199
rect 22327 4165 22336 4199
rect 22284 4156 22336 4165
rect 22652 4156 22704 4208
rect 5448 4020 5500 4072
rect 3056 3995 3108 4004
rect 3056 3961 3065 3995
rect 3065 3961 3099 3995
rect 3099 3961 3108 3995
rect 3056 3952 3108 3961
rect 6644 3884 6696 3936
rect 7104 3884 7156 3936
rect 10876 4088 10928 4140
rect 11980 4088 12032 4140
rect 16764 4088 16816 4140
rect 19708 4088 19760 4140
rect 25780 4088 25832 4140
rect 25872 4088 25924 4140
rect 10968 4020 11020 4072
rect 13268 4020 13320 4072
rect 15568 4020 15620 4072
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 9588 3952 9640 4004
rect 11796 3952 11848 4004
rect 11704 3884 11756 3936
rect 12256 3884 12308 3936
rect 13728 3884 13780 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 19524 3884 19576 3936
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 26424 3884 26476 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 4160 3723 4212 3732
rect 4160 3689 4169 3723
rect 4169 3689 4203 3723
rect 4203 3689 4212 3723
rect 4160 3680 4212 3689
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 8576 3680 8628 3732
rect 13084 3680 13136 3732
rect 15384 3680 15436 3732
rect 17132 3680 17184 3732
rect 20536 3680 20588 3732
rect 23020 3680 23072 3732
rect 25044 3680 25096 3732
rect 5264 3612 5316 3664
rect 7012 3612 7064 3664
rect 10508 3612 10560 3664
rect 12072 3612 12124 3664
rect 14464 3612 14516 3664
rect 1584 3544 1636 3596
rect 3792 3544 3844 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 6644 3544 6696 3596
rect 10692 3544 10744 3596
rect 10876 3587 10928 3596
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 1308 3476 1360 3528
rect 5724 3519 5776 3528
rect 5724 3485 5758 3519
rect 5758 3485 5776 3519
rect 5724 3476 5776 3485
rect 14004 3544 14056 3596
rect 19248 3544 19300 3596
rect 22284 3544 22336 3596
rect 26424 3544 26476 3596
rect 26976 3587 27028 3596
rect 26976 3553 26985 3587
rect 26985 3553 27019 3587
rect 27019 3553 27028 3587
rect 26976 3544 27028 3553
rect 1400 3408 1452 3460
rect 9312 3408 9364 3460
rect 13176 3476 13228 3528
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 16856 3476 16908 3528
rect 19340 3476 19392 3528
rect 20812 3519 20864 3528
rect 20812 3485 20846 3519
rect 20846 3485 20864 3519
rect 20812 3476 20864 3485
rect 22468 3476 22520 3528
rect 22652 3519 22704 3528
rect 22652 3485 22675 3519
rect 22675 3485 22704 3519
rect 22652 3476 22704 3485
rect 26884 3476 26936 3528
rect 6184 3340 6236 3392
rect 12900 3451 12952 3460
rect 12900 3417 12909 3451
rect 12909 3417 12943 3451
rect 12943 3417 12952 3451
rect 12900 3408 12952 3417
rect 12624 3340 12676 3392
rect 13360 3408 13412 3460
rect 16212 3408 16264 3460
rect 20904 3408 20956 3460
rect 15200 3340 15252 3392
rect 16028 3340 16080 3392
rect 16304 3340 16356 3392
rect 25596 3408 25648 3460
rect 24216 3340 24268 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 3608 3179 3660 3188
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 11060 3136 11112 3188
rect 12624 3136 12676 3188
rect 13728 3136 13780 3188
rect 14832 3136 14884 3188
rect 15292 3136 15344 3188
rect 16488 3136 16540 3188
rect 11704 3068 11756 3120
rect 15200 3068 15252 3120
rect 17684 3068 17736 3120
rect 17868 3068 17920 3120
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 20720 3136 20772 3188
rect 22928 3136 22980 3188
rect 18880 3068 18932 3120
rect 19524 3068 19576 3120
rect 1584 3000 1636 3052
rect 1952 3000 2004 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 3792 3000 3844 3052
rect 4160 3000 4212 3052
rect 9312 3000 9364 3052
rect 9864 3000 9916 3052
rect 10876 3000 10928 3052
rect 11980 3000 12032 3052
rect 14556 3000 14608 3052
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 14740 2932 14792 2984
rect 11060 2864 11112 2916
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16856 3043 16908 3052
rect 15660 2932 15712 2984
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 20720 3000 20772 3052
rect 20904 3000 20956 3052
rect 22284 3068 22336 3120
rect 24032 3068 24084 3120
rect 24216 3111 24268 3120
rect 24216 3077 24250 3111
rect 24250 3077 24268 3111
rect 24216 3068 24268 3077
rect 22192 3000 22244 3052
rect 23296 3000 23348 3052
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 19340 2932 19392 2984
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 5724 2796 5776 2805
rect 15752 2796 15804 2848
rect 16396 2796 16448 2848
rect 18144 2796 18196 2848
rect 24860 2796 24912 2848
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 5816 2592 5868 2644
rect 9404 2592 9456 2644
rect 12072 2592 12124 2644
rect 12256 2592 12308 2644
rect 12808 2592 12860 2644
rect 13820 2592 13872 2644
rect 17960 2635 18012 2644
rect 17960 2601 17969 2635
rect 17969 2601 18003 2635
rect 18003 2601 18012 2635
rect 17960 2592 18012 2601
rect 18144 2592 18196 2644
rect 18880 2635 18932 2644
rect 18880 2601 18889 2635
rect 18889 2601 18923 2635
rect 18923 2601 18932 2635
rect 18880 2592 18932 2601
rect 18972 2592 19024 2644
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 12256 2456 12308 2508
rect 5448 2388 5500 2440
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6184 2431 6236 2440
rect 6184 2397 6218 2431
rect 6218 2397 6236 2431
rect 6184 2388 6236 2397
rect 10876 2388 10928 2440
rect 11060 2388 11112 2440
rect 12440 2388 12492 2440
rect 16212 2567 16264 2576
rect 16212 2533 16221 2567
rect 16221 2533 16255 2567
rect 16255 2533 16264 2567
rect 16212 2524 16264 2533
rect 14740 2456 14792 2508
rect 17040 2456 17092 2508
rect 13084 2431 13136 2440
rect 13084 2397 13094 2431
rect 13094 2397 13128 2431
rect 13128 2397 13136 2431
rect 13084 2388 13136 2397
rect 13176 2388 13228 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 14648 2388 14700 2440
rect 17316 2431 17368 2440
rect 17316 2397 17325 2431
rect 17325 2397 17359 2431
rect 17359 2397 17368 2431
rect 17316 2388 17368 2397
rect 1676 2320 1728 2372
rect 6460 2320 6512 2372
rect 15292 2320 15344 2372
rect 13084 2252 13136 2304
rect 17316 2252 17368 2304
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 17684 2252 17736 2304
rect 17776 2252 17828 2304
rect 18328 2524 18380 2576
rect 20628 2524 20680 2576
rect 18052 2456 18104 2508
rect 18788 2456 18840 2508
rect 19156 2388 19208 2440
rect 19248 2320 19300 2372
rect 20996 2252 21048 2304
rect 22284 2388 22336 2440
rect 24124 2592 24176 2644
rect 23940 2456 23992 2508
rect 26976 2499 27028 2508
rect 26976 2465 26985 2499
rect 26985 2465 27019 2499
rect 27019 2465 27028 2499
rect 26976 2456 27028 2465
rect 25688 2388 25740 2440
rect 25964 2388 26016 2440
rect 22376 2320 22428 2372
rect 24860 2363 24912 2372
rect 24860 2329 24894 2363
rect 24894 2329 24912 2363
rect 24860 2320 24912 2329
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 1952 1912 2004 1964
rect 4160 1955 4212 1964
rect 4160 1921 4169 1955
rect 4169 1921 4203 1955
rect 4203 1921 4212 1955
rect 4160 1912 4212 1921
rect 7380 2048 7432 2100
rect 9312 2091 9364 2100
rect 9312 2057 9321 2091
rect 9321 2057 9355 2091
rect 9355 2057 9364 2091
rect 9312 2048 9364 2057
rect 9588 1980 9640 2032
rect 11244 1980 11296 2032
rect 13636 2048 13688 2100
rect 14004 2048 14056 2100
rect 15292 2048 15344 2100
rect 12164 1980 12216 2032
rect 3424 1887 3476 1896
rect 3424 1853 3433 1887
rect 3433 1853 3467 1887
rect 3467 1853 3476 1887
rect 3424 1844 3476 1853
rect 9864 1912 9916 1964
rect 12624 1980 12676 2032
rect 12532 1955 12584 1964
rect 12532 1921 12541 1955
rect 12541 1921 12575 1955
rect 12575 1921 12584 1955
rect 12532 1912 12584 1921
rect 13452 1980 13504 2032
rect 15752 1980 15804 2032
rect 16304 1980 16356 2032
rect 17500 1980 17552 2032
rect 17684 1980 17736 2032
rect 19708 1980 19760 2032
rect 21272 2091 21324 2100
rect 21272 2057 21281 2091
rect 21281 2057 21315 2091
rect 21315 2057 21324 2091
rect 21272 2048 21324 2057
rect 22284 2048 22336 2100
rect 23296 2048 23348 2100
rect 21640 1980 21692 2032
rect 5632 1844 5684 1896
rect 5908 1844 5960 1896
rect 8208 1708 8260 1760
rect 11888 1751 11940 1760
rect 11888 1717 11897 1751
rect 11897 1717 11931 1751
rect 11931 1717 11940 1751
rect 11888 1708 11940 1717
rect 14556 1708 14608 1760
rect 17040 1912 17092 1964
rect 15660 1708 15712 1760
rect 20720 1955 20772 1964
rect 20720 1921 20730 1955
rect 20730 1921 20764 1955
rect 20764 1921 20772 1955
rect 20720 1912 20772 1921
rect 20996 1955 21048 1964
rect 20996 1921 21005 1955
rect 21005 1921 21039 1955
rect 21039 1921 21048 1955
rect 20996 1912 21048 1921
rect 21088 1955 21140 1964
rect 22652 1980 22704 2032
rect 23664 1980 23716 2032
rect 24124 2023 24176 2032
rect 24124 1989 24136 2023
rect 24136 1989 24176 2023
rect 24124 1980 24176 1989
rect 24216 1980 24268 2032
rect 24860 1980 24912 2032
rect 21088 1921 21102 1955
rect 21102 1921 21136 1955
rect 21136 1921 21140 1955
rect 21088 1912 21140 1921
rect 23020 1912 23072 1964
rect 23940 1912 23992 1964
rect 21456 1844 21508 1896
rect 25780 1912 25832 1964
rect 25964 1844 26016 1896
rect 4423 1606 4475 1658
rect 4487 1606 4539 1658
rect 4551 1606 4603 1658
rect 4615 1606 4667 1658
rect 4679 1606 4731 1658
rect 11369 1606 11421 1658
rect 11433 1606 11485 1658
rect 11497 1606 11549 1658
rect 11561 1606 11613 1658
rect 11625 1606 11677 1658
rect 18315 1606 18367 1658
rect 18379 1606 18431 1658
rect 18443 1606 18495 1658
rect 18507 1606 18559 1658
rect 18571 1606 18623 1658
rect 25261 1606 25313 1658
rect 25325 1606 25377 1658
rect 25389 1606 25441 1658
rect 25453 1606 25505 1658
rect 25517 1606 25569 1658
rect 5632 1504 5684 1556
rect 11888 1504 11940 1556
rect 14556 1547 14608 1556
rect 14556 1513 14565 1547
rect 14565 1513 14599 1547
rect 14599 1513 14608 1547
rect 14556 1504 14608 1513
rect 16672 1504 16724 1556
rect 17776 1504 17828 1556
rect 14096 1436 14148 1488
rect 1952 1411 2004 1420
rect 1952 1377 1961 1411
rect 1961 1377 1995 1411
rect 1995 1377 2004 1411
rect 1952 1368 2004 1377
rect 13084 1368 13136 1420
rect 8300 1300 8352 1352
rect 9404 1343 9456 1352
rect 9404 1309 9438 1343
rect 9438 1309 9456 1343
rect 9404 1300 9456 1309
rect 11980 1343 12032 1352
rect 11980 1309 11989 1343
rect 11989 1309 12023 1343
rect 12023 1309 12032 1343
rect 11980 1300 12032 1309
rect 2228 1275 2280 1284
rect 2228 1241 2262 1275
rect 2262 1241 2280 1275
rect 2228 1232 2280 1241
rect 3332 1207 3384 1216
rect 3332 1173 3341 1207
rect 3341 1173 3375 1207
rect 3375 1173 3384 1207
rect 3332 1164 3384 1173
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 9496 1232 9548 1284
rect 12348 1232 12400 1284
rect 15476 1300 15528 1352
rect 15752 1343 15804 1352
rect 15752 1309 15761 1343
rect 15761 1309 15795 1343
rect 15795 1309 15804 1343
rect 15752 1300 15804 1309
rect 16028 1343 16080 1352
rect 16028 1309 16037 1343
rect 16037 1309 16071 1343
rect 16071 1309 16080 1343
rect 16028 1300 16080 1309
rect 16120 1343 16172 1352
rect 16120 1309 16129 1343
rect 16129 1309 16163 1343
rect 16163 1309 16172 1343
rect 16120 1300 16172 1309
rect 16396 1300 16448 1352
rect 15936 1275 15988 1284
rect 15936 1241 15945 1275
rect 15945 1241 15979 1275
rect 15979 1241 15988 1275
rect 15936 1232 15988 1241
rect 10324 1164 10376 1216
rect 10508 1207 10560 1216
rect 10508 1173 10517 1207
rect 10517 1173 10551 1207
rect 10551 1173 10560 1207
rect 10508 1164 10560 1173
rect 14740 1164 14792 1216
rect 18052 1300 18104 1352
rect 18420 1232 18472 1284
rect 21456 1368 21508 1420
rect 19524 1300 19576 1352
rect 20536 1300 20588 1352
rect 20904 1343 20956 1352
rect 20904 1309 20913 1343
rect 20913 1309 20947 1343
rect 20947 1309 20956 1343
rect 20904 1300 20956 1309
rect 21088 1343 21140 1352
rect 21088 1309 21097 1343
rect 21097 1309 21131 1343
rect 21131 1309 21140 1343
rect 21088 1300 21140 1309
rect 22560 1504 22612 1556
rect 25964 1504 26016 1556
rect 22284 1300 22336 1352
rect 23388 1300 23440 1352
rect 26976 1300 27028 1352
rect 20168 1275 20220 1284
rect 20168 1241 20177 1275
rect 20177 1241 20211 1275
rect 20211 1241 20220 1275
rect 20168 1232 20220 1241
rect 24032 1232 24084 1284
rect 25044 1232 25096 1284
rect 17868 1164 17920 1216
rect 19248 1164 19300 1216
rect 20628 1164 20680 1216
rect 23756 1207 23808 1216
rect 23756 1173 23765 1207
rect 23765 1173 23799 1207
rect 23799 1173 23808 1207
rect 23756 1164 23808 1173
rect 25780 1164 25832 1216
rect 7896 1062 7948 1114
rect 7960 1062 8012 1114
rect 8024 1062 8076 1114
rect 8088 1062 8140 1114
rect 8152 1062 8204 1114
rect 14842 1062 14894 1114
rect 14906 1062 14958 1114
rect 14970 1062 15022 1114
rect 15034 1062 15086 1114
rect 15098 1062 15150 1114
rect 21788 1062 21840 1114
rect 21852 1062 21904 1114
rect 21916 1062 21968 1114
rect 21980 1062 22032 1114
rect 22044 1062 22096 1114
rect 28734 1062 28786 1114
rect 28798 1062 28850 1114
rect 28862 1062 28914 1114
rect 28926 1062 28978 1114
rect 28990 1062 29042 1114
rect 15936 960 15988 1012
rect 21088 960 21140 1012
rect 19708 892 19760 944
rect 23756 960 23808 1012
rect 20168 824 20220 876
rect 23664 824 23716 876
<< metal2 >>
rect 7896 32668 8204 32677
rect 7896 32666 7902 32668
rect 7958 32666 7982 32668
rect 8038 32666 8062 32668
rect 8118 32666 8142 32668
rect 8198 32666 8204 32668
rect 7958 32614 7960 32666
rect 8140 32614 8142 32666
rect 7896 32612 7902 32614
rect 7958 32612 7982 32614
rect 8038 32612 8062 32614
rect 8118 32612 8142 32614
rect 8198 32612 8204 32614
rect 7896 32603 8204 32612
rect 14842 32668 15150 32677
rect 14842 32666 14848 32668
rect 14904 32666 14928 32668
rect 14984 32666 15008 32668
rect 15064 32666 15088 32668
rect 15144 32666 15150 32668
rect 14904 32614 14906 32666
rect 15086 32614 15088 32666
rect 14842 32612 14848 32614
rect 14904 32612 14928 32614
rect 14984 32612 15008 32614
rect 15064 32612 15088 32614
rect 15144 32612 15150 32614
rect 14842 32603 15150 32612
rect 21788 32668 22096 32677
rect 21788 32666 21794 32668
rect 21850 32666 21874 32668
rect 21930 32666 21954 32668
rect 22010 32666 22034 32668
rect 22090 32666 22096 32668
rect 21850 32614 21852 32666
rect 22032 32614 22034 32666
rect 21788 32612 21794 32614
rect 21850 32612 21874 32614
rect 21930 32612 21954 32614
rect 22010 32612 22034 32614
rect 22090 32612 22096 32614
rect 21788 32603 22096 32612
rect 28734 32668 29042 32677
rect 28734 32666 28740 32668
rect 28796 32666 28820 32668
rect 28876 32666 28900 32668
rect 28956 32666 28980 32668
rect 29036 32666 29042 32668
rect 28796 32614 28798 32666
rect 28978 32614 28980 32666
rect 28734 32612 28740 32614
rect 28796 32612 28820 32614
rect 28876 32612 28900 32614
rect 28956 32612 28980 32614
rect 29036 32612 29042 32614
rect 28734 32603 29042 32612
rect 4344 32564 4396 32570
rect 4344 32506 4396 32512
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 11244 32564 11296 32570
rect 11244 32506 11296 32512
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1492 31340 1544 31346
rect 1492 31282 1544 31288
rect 1504 24206 1532 31282
rect 1596 30054 1624 31758
rect 1584 30048 1636 30054
rect 1584 29990 1636 29996
rect 1584 29504 1636 29510
rect 1688 29492 1716 32370
rect 2778 32328 2834 32337
rect 2778 32263 2834 32272
rect 3332 32292 3384 32298
rect 2792 32026 2820 32263
rect 3332 32234 3384 32240
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 3344 31890 3372 32234
rect 3332 31884 3384 31890
rect 3332 31826 3384 31832
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 1860 30320 1912 30326
rect 1860 30262 1912 30268
rect 1636 29464 1716 29492
rect 1584 29446 1636 29452
rect 1596 26382 1624 29446
rect 1768 29300 1820 29306
rect 1768 29242 1820 29248
rect 1676 28076 1728 28082
rect 1676 28018 1728 28024
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1688 25906 1716 28018
rect 1676 25900 1728 25906
rect 1676 25842 1728 25848
rect 1780 24206 1808 29242
rect 1872 27130 1900 30262
rect 1952 29640 2004 29646
rect 1952 29582 2004 29588
rect 1964 28082 1992 29582
rect 2056 28558 2084 31282
rect 2608 30938 2636 31282
rect 3884 31272 3936 31278
rect 3884 31214 3936 31220
rect 3792 31136 3844 31142
rect 3792 31078 3844 31084
rect 2596 30932 2648 30938
rect 2596 30874 2648 30880
rect 2136 30252 2188 30258
rect 2136 30194 2188 30200
rect 2228 30252 2280 30258
rect 2228 30194 2280 30200
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 2044 28552 2096 28558
rect 2044 28494 2096 28500
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 2044 27464 2096 27470
rect 2044 27406 2096 27412
rect 1860 27124 1912 27130
rect 1912 27084 1992 27112
rect 1860 27066 1912 27072
rect 1860 26920 1912 26926
rect 1860 26862 1912 26868
rect 1872 24750 1900 26862
rect 1964 25498 1992 27084
rect 2056 26450 2084 27406
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 2056 25838 2084 26386
rect 2044 25832 2096 25838
rect 2044 25774 2096 25780
rect 1952 25492 2004 25498
rect 1952 25434 2004 25440
rect 2056 25294 2084 25774
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1492 24200 1544 24206
rect 846 24168 902 24177
rect 1492 24142 1544 24148
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 846 24103 848 24112
rect 900 24103 902 24112
rect 848 24074 900 24080
rect 2056 24070 2084 25230
rect 2148 24410 2176 30194
rect 2240 29782 2268 30194
rect 2228 29776 2280 29782
rect 2228 29718 2280 29724
rect 2424 29646 2452 30194
rect 2504 30048 2556 30054
rect 2504 29990 2556 29996
rect 2412 29640 2464 29646
rect 2412 29582 2464 29588
rect 2412 29232 2464 29238
rect 2412 29174 2464 29180
rect 2424 27962 2452 29174
rect 2516 28082 2544 29990
rect 2884 29306 2912 30194
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2424 27934 2544 27962
rect 2412 26920 2464 26926
rect 2412 26862 2464 26868
rect 2424 26586 2452 26862
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2136 24404 2188 24410
rect 2136 24346 2188 24352
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 664 16584 716 16590
rect 664 16526 716 16532
rect 676 16017 704 16526
rect 662 16008 718 16017
rect 662 15943 718 15952
rect 572 14408 624 14414
rect 572 14350 624 14356
rect 584 13977 612 14350
rect 570 13968 626 13977
rect 570 13903 626 13912
rect 756 12232 808 12238
rect 756 12174 808 12180
rect 768 11937 796 12174
rect 754 11928 810 11937
rect 754 11863 810 11872
rect 848 10056 900 10062
rect 848 9998 900 10004
rect 860 9897 888 9998
rect 846 9888 902 9897
rect 846 9823 902 9832
rect 940 7880 992 7886
rect 938 7848 940 7857
rect 992 7848 994 7857
rect 938 7783 994 7792
rect 1306 3768 1362 3777
rect 1306 3703 1362 3712
rect 1320 3534 1348 3703
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1412 3466 1440 22374
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 4622 1532 20742
rect 1596 16574 1624 23258
rect 1872 22030 1900 24006
rect 1950 22128 2006 22137
rect 1950 22063 1952 22072
rect 2004 22063 2006 22072
rect 1952 22034 2004 22040
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1688 17202 1716 17682
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1688 16794 1716 17138
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 16674 1716 16730
rect 1688 16646 1808 16674
rect 1596 16546 1716 16574
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9586 1624 10406
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1596 9042 1624 9522
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 6866 1624 8978
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6322 1624 6802
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 5778 1624 6258
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1596 4690 1624 5714
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1596 4146 1624 4626
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1596 3602 1624 4082
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1596 3058 1624 3538
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1688 2650 1716 16546
rect 1780 15706 1808 16646
rect 1872 16250 1900 21966
rect 2148 21622 2176 21966
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 2240 19990 2268 24142
rect 2332 24070 2360 24142
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 2332 22030 2360 24006
rect 2516 23610 2544 27934
rect 2608 27674 2636 29106
rect 3436 28558 3464 29446
rect 3424 28552 3476 28558
rect 3424 28494 3476 28500
rect 2688 28484 2740 28490
rect 2688 28426 2740 28432
rect 2596 27668 2648 27674
rect 2596 27610 2648 27616
rect 2608 23798 2636 27610
rect 2700 26994 2728 28426
rect 3516 28416 3568 28422
rect 3516 28358 3568 28364
rect 3424 28144 3476 28150
rect 3424 28086 3476 28092
rect 2688 26988 2740 26994
rect 2688 26930 2740 26936
rect 2700 26450 2728 26930
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2688 26240 2740 26246
rect 2688 26182 2740 26188
rect 2700 24818 2728 26182
rect 3436 25498 3464 28086
rect 3528 28082 3556 28358
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3804 24954 3832 31078
rect 3896 29578 3924 31214
rect 4252 31136 4304 31142
rect 4252 31078 4304 31084
rect 4264 30734 4292 31078
rect 4356 30734 4384 32506
rect 5184 32450 5212 32506
rect 5092 32434 5212 32450
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 5092 32428 5224 32434
rect 5092 32422 5172 32428
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4423 32124 4731 32133
rect 4423 32122 4429 32124
rect 4485 32122 4509 32124
rect 4565 32122 4589 32124
rect 4645 32122 4669 32124
rect 4725 32122 4731 32124
rect 4485 32070 4487 32122
rect 4667 32070 4669 32122
rect 4423 32068 4429 32070
rect 4485 32068 4509 32070
rect 4565 32068 4589 32070
rect 4645 32068 4669 32070
rect 4725 32068 4731 32070
rect 4423 32059 4731 32068
rect 4816 31822 4844 32302
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4436 31816 4488 31822
rect 4436 31758 4488 31764
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4448 31142 4476 31758
rect 4712 31748 4764 31754
rect 4712 31690 4764 31696
rect 4724 31226 4752 31690
rect 4816 31346 4844 31758
rect 4804 31340 4856 31346
rect 4804 31282 4856 31288
rect 4724 31198 4844 31226
rect 4436 31136 4488 31142
rect 4436 31078 4488 31084
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 4252 30728 4304 30734
rect 4252 30670 4304 30676
rect 4344 30728 4396 30734
rect 4344 30670 4396 30676
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3976 30320 4028 30326
rect 3974 30288 3976 30297
rect 4028 30288 4030 30297
rect 3974 30223 4030 30232
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3976 29096 4028 29102
rect 3976 29038 4028 29044
rect 3988 27402 4016 29038
rect 4066 28248 4122 28257
rect 4172 28218 4200 30534
rect 4344 30116 4396 30122
rect 4344 30058 4396 30064
rect 4252 30048 4304 30054
rect 4252 29990 4304 29996
rect 4264 29782 4292 29990
rect 4252 29776 4304 29782
rect 4252 29718 4304 29724
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 4264 28218 4292 29582
rect 4356 28490 4384 30058
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 4344 28484 4396 28490
rect 4344 28426 4396 28432
rect 4066 28183 4122 28192
rect 4160 28212 4212 28218
rect 4080 27674 4108 28183
rect 4160 28154 4212 28160
rect 4252 28212 4304 28218
rect 4252 28154 4304 28160
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 4080 27130 4108 27406
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 4172 27130 4200 27270
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3148 24880 3200 24886
rect 3148 24822 3200 24828
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2700 24206 2728 24754
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2516 23582 2636 23610
rect 2504 22568 2556 22574
rect 2504 22510 2556 22516
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2332 21690 2360 21966
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2228 19984 2280 19990
rect 2228 19926 2280 19932
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1780 15094 1808 15642
rect 1872 15162 1900 16050
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1768 15088 1820 15094
rect 1768 15030 1820 15036
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14618 1808 14758
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1872 14414 1900 15098
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1872 12306 1900 14350
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 1780 10266 1808 11562
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1872 9178 1900 9454
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 8906 1992 16934
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 14822 2268 16526
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 15162 2452 15438
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 13938 2452 14758
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 5817 1808 7346
rect 1766 5808 1822 5817
rect 1766 5743 1822 5752
rect 2516 3058 2544 22510
rect 2608 17610 2636 23582
rect 2976 18426 3004 24754
rect 3160 24274 3188 24822
rect 3884 24812 3936 24818
rect 3884 24754 3936 24760
rect 3896 24410 3924 24754
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18834 3096 19110
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16726 2636 17138
rect 2700 17066 2728 17818
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 17184 2820 17614
rect 3068 17338 3096 18022
rect 3160 17882 3188 21490
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3252 17338 3280 20470
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3344 19378 3372 19654
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3344 17338 3372 18226
rect 3436 18222 3464 19178
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 2872 17196 2924 17202
rect 2792 17156 2872 17184
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2596 16584 2648 16590
rect 2700 16574 2728 17002
rect 2648 16546 2728 16574
rect 2596 16526 2648 16532
rect 2792 16114 2820 17156
rect 2872 17138 2924 17144
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2608 14822 2636 16050
rect 2792 15978 2820 16050
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2976 15366 3004 16594
rect 3344 16590 3372 17274
rect 3436 16590 3464 18158
rect 3528 17202 3556 18634
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3160 15978 3188 16458
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3054 15600 3110 15609
rect 3054 15535 3110 15544
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 10742 2636 14758
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9722 2636 9998
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 2700 6798 2728 6831
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2792 6322 2820 7142
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5370 2820 5510
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1688 2378 1716 2586
rect 1964 2514 1992 2994
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 1964 1970 1992 2450
rect 1952 1964 2004 1970
rect 1952 1906 2004 1912
rect 1964 1426 1992 1906
rect 2884 1737 2912 14962
rect 2976 14618 3004 15302
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6866 3004 7142
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 5352 3004 6802
rect 3068 5914 3096 15535
rect 3160 6662 3188 15914
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3252 13326 3280 14214
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3344 9178 3372 16526
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 10606 3464 11494
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 10062 3464 10542
rect 3528 10266 3556 11018
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3056 5364 3108 5370
rect 2976 5324 3056 5352
rect 3056 5306 3108 5312
rect 3146 5128 3202 5137
rect 3146 5063 3202 5072
rect 3160 4826 3188 5063
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3054 4040 3110 4049
rect 3054 3975 3056 3984
rect 3108 3975 3110 3984
rect 3056 3946 3108 3952
rect 3620 3194 3648 23666
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3712 6390 3740 19450
rect 3896 18057 3924 21898
rect 3988 19446 4016 25638
rect 4080 24682 4108 25842
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 4172 24426 4200 26726
rect 4264 26382 4292 27950
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 4712 26920 4764 26926
rect 4712 26862 4764 26868
rect 4724 26790 4752 26862
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 4816 26314 4844 31198
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 4342 26208 4398 26217
rect 4342 26143 4398 26152
rect 4252 25764 4304 25770
rect 4252 25706 4304 25712
rect 4264 25294 4292 25706
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 4172 24398 4292 24426
rect 4160 24336 4212 24342
rect 4160 24278 4212 24284
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 4080 22030 4108 24074
rect 4172 23526 4200 24278
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4160 23044 4212 23050
rect 4160 22986 4212 22992
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4066 20088 4122 20097
rect 4172 20074 4200 22986
rect 4264 20602 4292 24398
rect 4356 24342 4384 26143
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4528 25220 4580 25226
rect 4528 25162 4580 25168
rect 4540 24954 4568 25162
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4632 24682 4660 24754
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4344 24336 4396 24342
rect 4344 24278 4396 24284
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4540 24070 4568 24142
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4710 23896 4766 23905
rect 4710 23831 4766 23840
rect 4724 23798 4752 23831
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4122 20046 4200 20074
rect 4066 20023 4122 20032
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 4264 18290 4292 20334
rect 4356 18970 4384 21490
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4816 20398 4844 25774
rect 4908 24682 4936 32166
rect 5092 31482 5120 32422
rect 5172 32370 5224 32376
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8208 32360 8260 32366
rect 8208 32302 8260 32308
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5184 31958 5212 32234
rect 5264 32020 5316 32026
rect 5264 31962 5316 31968
rect 5172 31952 5224 31958
rect 5172 31894 5224 31900
rect 5080 31476 5132 31482
rect 5080 31418 5132 31424
rect 5184 31210 5212 31894
rect 5172 31204 5224 31210
rect 5172 31146 5224 31152
rect 5080 30116 5132 30122
rect 5080 30058 5132 30064
rect 4988 28076 5040 28082
rect 4988 28018 5040 28024
rect 5000 25838 5028 28018
rect 4988 25832 5040 25838
rect 4988 25774 5040 25780
rect 5000 25362 5028 25774
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 5000 24750 5028 25298
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4896 24676 4948 24682
rect 4896 24618 4948 24624
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4908 22778 4936 24142
rect 5000 23866 5028 24686
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 4986 23760 5042 23769
rect 4986 23695 4988 23704
rect 5040 23695 5042 23704
rect 4988 23666 5040 23672
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4908 20942 4936 22578
rect 5092 22098 5120 30058
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 5184 28694 5212 29786
rect 5172 28688 5224 28694
rect 5172 28630 5224 28636
rect 5172 28416 5224 28422
rect 5172 28358 5224 28364
rect 5184 26858 5212 28358
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 5184 25838 5212 26794
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 5184 23769 5212 25298
rect 5276 23905 5304 31962
rect 8220 31822 8248 32302
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 5920 31482 5948 31622
rect 5908 31476 5960 31482
rect 5908 31418 5960 31424
rect 6920 31476 6972 31482
rect 6920 31418 6972 31424
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 5908 31204 5960 31210
rect 5908 31146 5960 31152
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5460 29170 5488 30194
rect 5644 30190 5672 30738
rect 5632 30184 5684 30190
rect 5632 30126 5684 30132
rect 5920 29782 5948 31146
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 6000 30660 6052 30666
rect 6000 30602 6052 30608
rect 5908 29776 5960 29782
rect 5908 29718 5960 29724
rect 5540 29640 5592 29646
rect 5540 29582 5592 29588
rect 5448 29164 5500 29170
rect 5368 29124 5448 29152
rect 5368 26602 5396 29124
rect 5448 29106 5500 29112
rect 5552 29034 5580 29582
rect 5816 29572 5868 29578
rect 5816 29514 5868 29520
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5644 29238 5672 29446
rect 5632 29232 5684 29238
rect 5632 29174 5684 29180
rect 5540 29028 5592 29034
rect 5540 28970 5592 28976
rect 5724 28960 5776 28966
rect 5724 28902 5776 28908
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 27062 5488 28358
rect 5736 28082 5764 28902
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5644 26790 5672 27406
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5724 26784 5776 26790
rect 5724 26726 5776 26732
rect 5368 26574 5488 26602
rect 5356 26512 5408 26518
rect 5356 26454 5408 26460
rect 5368 26353 5396 26454
rect 5354 26344 5410 26353
rect 5354 26279 5410 26288
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5368 26042 5396 26182
rect 5460 26042 5488 26574
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 5262 23896 5318 23905
rect 5262 23831 5318 23840
rect 5170 23760 5226 23769
rect 5170 23695 5226 23704
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5276 23118 5304 23666
rect 5368 23254 5396 25230
rect 5460 24818 5488 25978
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5460 23866 5488 24754
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5276 21894 5304 23054
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5276 21418 5304 21830
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5368 21026 5396 21830
rect 5276 20998 5396 21026
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4816 18902 4844 20198
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 4264 17746 4292 18226
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 3804 16998 3832 17138
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 4264 16590 4292 17138
rect 4356 16658 4384 18770
rect 4816 18290 4844 18838
rect 4908 18834 4936 20878
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5000 20058 5028 20402
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 5000 18630 5028 19994
rect 5184 19922 5212 20538
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19378 5212 19654
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18290 5028 18566
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 4816 17746 4844 18226
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4816 17218 4844 17682
rect 5000 17678 5028 18226
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5092 17542 5120 19246
rect 5276 19174 5304 20998
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 19854 5396 20742
rect 5460 20602 5488 23666
rect 5552 23186 5580 26386
rect 5644 25906 5672 26726
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5644 25702 5672 25842
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5644 23186 5672 24890
rect 5736 24206 5764 26726
rect 5828 25498 5856 29514
rect 5920 28150 5948 29718
rect 5908 28144 5960 28150
rect 5908 28086 5960 28092
rect 6012 26382 6040 30602
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 6092 29028 6144 29034
rect 6092 28970 6144 28976
rect 6104 28558 6132 28970
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 27606 6132 28494
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 6104 26994 6132 27542
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 6000 26376 6052 26382
rect 5920 26336 6000 26364
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 5828 24818 5856 25298
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5724 24064 5776 24070
rect 5724 24006 5776 24012
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5736 22030 5764 24006
rect 5828 23798 5856 24754
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5828 21554 5856 23598
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5920 20466 5948 26336
rect 6000 26318 6052 26324
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5460 19334 5488 20334
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5368 19306 5488 19334
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5368 17660 5396 19306
rect 5552 18834 5580 19858
rect 5644 19854 5672 19994
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5644 19417 5672 19654
rect 5630 19408 5686 19417
rect 5630 19343 5686 19352
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18034 5580 18770
rect 5276 17632 5396 17660
rect 5460 18006 5580 18034
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5080 17264 5132 17270
rect 4816 17190 4936 17218
rect 5080 17206 5132 17212
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3988 15434 4016 15642
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3804 5914 3832 15030
rect 3988 14346 4016 15370
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3988 11558 4016 12174
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4080 10198 4108 13874
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13190 4292 13806
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12782 4292 13126
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4264 12442 4292 12718
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4252 12232 4304 12238
rect 4172 12192 4252 12220
rect 4172 11354 4200 12192
rect 4252 12174 4304 12180
rect 4356 11830 4384 16594
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4540 16017 4568 16390
rect 4526 16008 4582 16017
rect 4526 15943 4582 15952
rect 4724 15892 4752 16662
rect 4816 16454 4844 17070
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4724 15864 4844 15892
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4816 14362 4844 15864
rect 4908 15706 4936 17190
rect 5092 16998 5120 17206
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16114 5120 16934
rect 5276 16658 5304 17632
rect 5460 17610 5488 18006
rect 5736 17882 5764 19994
rect 5920 18834 5948 20402
rect 6012 18873 6040 25638
rect 6092 25220 6144 25226
rect 6092 25162 6144 25168
rect 6104 24954 6132 25162
rect 6092 24948 6144 24954
rect 6092 24890 6144 24896
rect 6196 24682 6224 30194
rect 6380 26994 6408 31078
rect 6564 30734 6592 31282
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6564 30258 6592 30670
rect 6932 30394 6960 31418
rect 7576 31278 7604 31758
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 7576 30802 7604 31214
rect 7668 30938 7696 31282
rect 7656 30932 7708 30938
rect 7656 30874 7708 30880
rect 8312 30870 8340 32370
rect 8392 32292 8444 32298
rect 8392 32234 8444 32240
rect 8300 30864 8352 30870
rect 8300 30806 8352 30812
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 6920 30388 6972 30394
rect 6840 30348 6920 30376
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6460 29640 6512 29646
rect 6564 29628 6592 30194
rect 6512 29600 6592 29628
rect 6460 29582 6512 29588
rect 6840 29510 6868 30348
rect 6920 30330 6972 30336
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 6920 30116 6972 30122
rect 6920 30058 6972 30064
rect 6932 29782 6960 30058
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 6920 29776 6972 29782
rect 6920 29718 6972 29724
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6736 29096 6788 29102
rect 6736 29038 6788 29044
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6656 28558 6684 28902
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6748 28082 6776 29038
rect 6932 28150 6960 29106
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6552 27668 6604 27674
rect 6552 27610 6604 27616
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6184 24676 6236 24682
rect 6184 24618 6236 24624
rect 6196 23186 6224 24618
rect 6276 24132 6328 24138
rect 6380 24120 6408 26930
rect 6460 26920 6512 26926
rect 6460 26862 6512 26868
rect 6328 24092 6408 24120
rect 6276 24074 6328 24080
rect 6380 23866 6408 24092
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 6472 23662 6500 26862
rect 6564 25974 6592 27610
rect 6748 26314 6776 28018
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 6736 26308 6788 26314
rect 6736 26250 6788 26256
rect 6552 25968 6604 25974
rect 6552 25910 6604 25916
rect 6644 24132 6696 24138
rect 6748 24120 6776 26250
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6696 24092 6776 24120
rect 6644 24074 6696 24080
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6472 23526 6500 23598
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6656 23186 6684 23462
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6184 23044 6236 23050
rect 6184 22986 6236 22992
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 5998 18864 6054 18873
rect 5908 18828 5960 18834
rect 5998 18799 6054 18808
rect 5908 18770 5960 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5920 18714 5948 18770
rect 5724 17876 5776 17882
rect 5552 17836 5724 17864
rect 5448 17604 5500 17610
rect 5368 17564 5448 17592
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5368 16114 5396 17564
rect 5448 17546 5500 17552
rect 5448 17060 5500 17066
rect 5552 17048 5580 17836
rect 5724 17818 5776 17824
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5500 17020 5580 17048
rect 5448 17002 5500 17008
rect 5552 16574 5580 17020
rect 5736 16998 5764 17682
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16794 5764 16934
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5460 16546 5580 16574
rect 5460 16182 5488 16546
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5080 16108 5132 16114
rect 5356 16108 5408 16114
rect 5132 16068 5212 16096
rect 5080 16050 5132 16056
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 4908 14822 4936 15642
rect 5000 15026 5028 16050
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14550 4936 14758
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4816 14334 4936 14362
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 14006 4568 14214
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12918 4568 13262
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4816 12434 4844 13330
rect 4724 12406 4844 12434
rect 4724 12238 4752 12406
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10266 4200 11086
rect 4264 10674 4292 11630
rect 4724 11626 4752 12174
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4068 10192 4120 10198
rect 4264 10146 4292 10610
rect 4068 10134 4120 10140
rect 4172 10118 4292 10146
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3896 6390 3924 7346
rect 4172 7290 4200 10118
rect 4356 10062 4384 11222
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4816 10266 4844 12310
rect 4908 11694 4936 14334
rect 5000 13734 5028 14418
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 12306 5028 13262
rect 5092 12918 5120 15438
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5184 12730 5212 16068
rect 5356 16050 5408 16056
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14074 5304 14962
rect 5368 14958 5396 16050
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 14414 5396 14894
rect 5460 14618 5488 16118
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5552 14618 5580 15982
rect 5644 15978 5672 16458
rect 5828 16250 5856 18702
rect 5920 18686 6040 18714
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5724 15904 5776 15910
rect 5644 15852 5724 15858
rect 5644 15846 5776 15852
rect 5644 15830 5764 15846
rect 5644 15570 5672 15830
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5736 14890 5764 15506
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5632 14544 5684 14550
rect 5460 14492 5632 14498
rect 5460 14486 5684 14492
rect 5460 14470 5672 14486
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5460 14260 5488 14470
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5368 14232 5488 14260
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13734 5304 13806
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13190 5304 13670
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5184 12702 5304 12730
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12374 5212 12582
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5276 12209 5304 12702
rect 5368 12322 5396 14232
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13326 5488 13738
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12442 5488 13262
rect 5552 12986 5580 14282
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12436 5500 12442
rect 5644 12434 5672 14350
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 13530 5764 13874
rect 5828 13802 5856 15302
rect 5920 14074 5948 18566
rect 6012 18426 6040 18686
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 17270 6132 19994
rect 6196 18426 6224 22986
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6656 22574 6684 22918
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6748 22030 6776 24092
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6274 20904 6330 20913
rect 6274 20839 6276 20848
rect 6328 20839 6330 20848
rect 6276 20810 6328 20816
rect 6288 20602 6316 20810
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6288 17592 6316 20334
rect 6380 19242 6408 21966
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6380 17882 6408 19178
rect 6472 18970 6500 21966
rect 6564 21690 6592 21966
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6564 19689 6592 19722
rect 6550 19680 6606 19689
rect 6550 19615 6606 19624
rect 6550 19408 6606 19417
rect 6550 19343 6552 19352
rect 6604 19343 6606 19352
rect 6552 19314 6604 19320
rect 6656 19310 6684 21490
rect 6748 20330 6776 21966
rect 6840 20602 6868 25978
rect 6932 25906 6960 27814
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 7024 25430 7052 29038
rect 7288 28688 7340 28694
rect 7288 28630 7340 28636
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 7116 26518 7144 26998
rect 7104 26512 7156 26518
rect 7104 26454 7156 26460
rect 7208 25974 7236 27950
rect 7196 25968 7248 25974
rect 7196 25910 7248 25916
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7116 25498 7144 25842
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7012 25424 7064 25430
rect 7300 25378 7328 28630
rect 7392 25498 7420 29786
rect 7484 29646 7512 30262
rect 7576 30258 7604 30738
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 7576 29646 7604 30194
rect 7668 30122 7696 30670
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 7656 30116 7708 30122
rect 7656 30058 7708 30064
rect 8312 29646 8340 30806
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 7484 28506 7512 29582
rect 7576 28762 7604 29582
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 7656 29028 7708 29034
rect 7656 28970 7708 28976
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 7564 28552 7616 28558
rect 7484 28500 7564 28506
rect 7484 28494 7616 28500
rect 7484 28478 7604 28494
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7484 28082 7512 28358
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7576 27130 7604 28478
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 7484 25514 7512 27066
rect 7668 27062 7696 28970
rect 8404 28694 8432 32234
rect 8392 28688 8444 28694
rect 8392 28630 8444 28636
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7760 27402 7788 28426
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7656 27056 7708 27062
rect 7656 26998 7708 27004
rect 7760 26994 7788 27338
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7380 25492 7432 25498
rect 7484 25486 7604 25514
rect 7380 25434 7432 25440
rect 7012 25366 7064 25372
rect 7116 25350 7328 25378
rect 7116 24970 7144 25350
rect 7392 25344 7420 25434
rect 7392 25316 7512 25344
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7024 24942 7144 24970
rect 7024 23866 7052 24942
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 21962 6960 23462
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7024 22234 7052 22578
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 7024 21162 7052 21830
rect 7116 21554 7144 23734
rect 7208 23730 7236 25230
rect 7484 25106 7512 25316
rect 7392 25078 7512 25106
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7208 21978 7236 22578
rect 7392 22574 7420 25078
rect 7576 24970 7604 25486
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7668 25226 7696 25298
rect 7656 25220 7708 25226
rect 7656 25162 7708 25168
rect 7484 24942 7604 24970
rect 7656 24948 7708 24954
rect 7380 22568 7432 22574
rect 7300 22528 7380 22556
rect 7300 22098 7328 22528
rect 7380 22510 7432 22516
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7380 22092 7432 22098
rect 7484 22094 7512 24942
rect 7656 24890 7708 24896
rect 7564 24880 7616 24886
rect 7564 24822 7616 24828
rect 7576 22556 7604 24822
rect 7668 22658 7696 24890
rect 7760 24750 7788 26930
rect 8312 26926 8340 27950
rect 8496 27470 8524 32438
rect 8588 32298 8616 32506
rect 9508 32366 9536 32506
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 11152 32360 11204 32366
rect 11152 32302 11204 32308
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 8588 31822 8616 32234
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 9036 31884 9088 31890
rect 9036 31826 9088 31832
rect 9496 31884 9548 31890
rect 9496 31826 9548 31832
rect 8576 31816 8628 31822
rect 8576 31758 8628 31764
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8588 27538 8616 28358
rect 8852 28212 8904 28218
rect 8852 28154 8904 28160
rect 8864 27674 8892 28154
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8852 27668 8904 27674
rect 8852 27610 8904 27616
rect 8576 27532 8628 27538
rect 8576 27474 8628 27480
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8220 26450 8248 26726
rect 8312 26586 8340 26862
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 8220 25158 8248 25366
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 8312 24206 8340 25230
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 8312 23866 8340 24142
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 7852 23526 7880 23802
rect 8404 23594 8432 27406
rect 8864 26586 8892 27610
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8496 25430 8524 26318
rect 8588 25498 8616 26318
rect 8852 26308 8904 26314
rect 8852 26250 8904 26256
rect 8864 25906 8892 26250
rect 8956 26042 8984 27882
rect 9048 27606 9076 31826
rect 9312 29028 9364 29034
rect 9312 28970 9364 28976
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8484 25424 8536 25430
rect 8484 25366 8536 25372
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 7668 22630 7880 22658
rect 7576 22528 7788 22556
rect 7484 22066 7604 22094
rect 7380 22034 7432 22040
rect 7208 21962 7328 21978
rect 7208 21956 7340 21962
rect 7208 21950 7288 21956
rect 7288 21898 7340 21904
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7116 21350 7144 21490
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6920 21140 6972 21146
rect 7024 21134 7144 21162
rect 7208 21146 7236 21490
rect 6920 21082 6972 21088
rect 6932 20806 6960 21082
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6460 17604 6512 17610
rect 6288 17564 6460 17592
rect 6460 17546 6512 17552
rect 6274 17504 6330 17513
rect 6274 17439 6330 17448
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16522 6040 17138
rect 6288 17134 6316 17439
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6196 16590 6224 16730
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 15366 6040 16458
rect 6196 16182 6224 16526
rect 6184 16176 6236 16182
rect 6288 16153 6316 17070
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6184 16118 6236 16124
rect 6274 16144 6330 16153
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 15609 6132 16050
rect 6196 15978 6224 16118
rect 6274 16079 6276 16088
rect 6328 16079 6330 16088
rect 6276 16050 6328 16056
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6090 15600 6146 15609
rect 6090 15535 6146 15544
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6012 13870 6040 14214
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12782 5764 13330
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5644 12406 5764 12434
rect 5448 12378 5500 12384
rect 5368 12294 5672 12322
rect 5356 12232 5408 12238
rect 5078 12200 5134 12209
rect 5078 12135 5080 12144
rect 5132 12135 5134 12144
rect 5262 12200 5318 12209
rect 5356 12174 5408 12180
rect 5262 12135 5318 12144
rect 5080 12106 5132 12112
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4448 9518 4476 9998
rect 4724 9722 4752 10134
rect 4908 10062 4936 11494
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4724 9518 4752 9658
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4712 9512 4764 9518
rect 4764 9460 4844 9466
rect 4712 9454 4844 9460
rect 4724 9438 4844 9454
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4816 9178 4844 9438
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4080 7262 4200 7290
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3896 5574 3924 6326
rect 3884 5568 3936 5574
rect 4080 5556 4108 7262
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 5710 4200 7142
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4080 5528 4200 5556
rect 3884 5510 3936 5516
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4146 3832 4966
rect 4080 4690 4108 5170
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3804 3602 3832 4082
rect 4172 3738 4200 5528
rect 4264 4554 4292 7686
rect 4356 5914 4384 7822
rect 4816 7206 4844 8910
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4802 7032 4858 7041
rect 4802 6967 4858 6976
rect 4816 6458 4844 6967
rect 4908 6662 4936 8774
rect 5000 8090 5028 11630
rect 5092 9654 5120 11630
rect 5276 11354 5304 11630
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5184 10674 5212 11290
rect 5264 11144 5316 11150
rect 5262 11112 5264 11121
rect 5316 11112 5318 11121
rect 5262 11047 5318 11056
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5184 10130 5212 10610
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5368 9874 5396 12174
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5460 11762 5488 12106
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11286 5488 11698
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5460 11014 5488 11222
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5644 10810 5672 12294
rect 5736 11626 5764 12406
rect 5828 11762 5856 13126
rect 5908 12776 5960 12782
rect 6012 12764 6040 13262
rect 6104 12986 6132 15438
rect 6380 15094 6408 16458
rect 6472 16096 6500 17546
rect 6564 17202 6592 18022
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6552 16108 6604 16114
rect 6472 16068 6552 16096
rect 6552 16050 6604 16056
rect 6564 15910 6592 16050
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5960 12736 6040 12764
rect 5908 12718 5960 12724
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5276 9846 5396 9874
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5092 7886 5120 9454
rect 5184 8906 5212 9522
rect 5276 9042 5304 9846
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 5184 5914 5212 8842
rect 5276 8634 5304 8978
rect 5368 8838 5396 9522
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 5184 4282 5212 5238
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 5276 3670 5304 8434
rect 5368 8022 5396 8774
rect 5460 8634 5488 10746
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5644 8498 5672 9522
rect 5828 9178 5856 11018
rect 5920 10810 5948 12718
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 9994 5948 10406
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 5778 5396 6598
rect 5460 6458 5488 8434
rect 5736 8362 5764 8910
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5552 7750 5580 8298
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5460 5710 5488 6394
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5552 5642 5580 7686
rect 5828 7546 5856 9114
rect 5920 8498 5948 9522
rect 6012 9450 6040 12378
rect 6104 12102 6132 12786
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6196 11898 6224 14894
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6092 11280 6144 11286
rect 6288 11234 6316 12786
rect 6380 12442 6408 14282
rect 6564 13870 6592 15642
rect 6656 15162 6684 18566
rect 6748 16794 6776 19654
rect 6932 19394 6960 20742
rect 7116 20505 7144 21134
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7300 20942 7328 21898
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7196 20868 7248 20874
rect 7196 20810 7248 20816
rect 7102 20496 7158 20505
rect 7102 20431 7158 20440
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19786 7144 20334
rect 7208 20058 7236 20810
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 6840 19378 6960 19394
rect 6828 19372 6960 19378
rect 6880 19366 6960 19372
rect 6828 19314 6880 19320
rect 6932 17746 6960 19366
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6840 16454 6868 17614
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17202 6960 17478
rect 7024 17338 7052 19246
rect 7116 18970 7144 19722
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18760 7156 18766
rect 7102 18728 7104 18737
rect 7156 18728 7158 18737
rect 7102 18663 7158 18672
rect 7208 18408 7236 19654
rect 7300 19258 7328 20742
rect 7392 19446 7420 22034
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7484 20913 7512 21898
rect 7470 20904 7526 20913
rect 7470 20839 7526 20848
rect 7484 20806 7512 20839
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7300 19230 7420 19258
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7116 18380 7236 18408
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7116 16726 7144 18380
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16114 7052 16390
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6932 16017 6960 16050
rect 6918 16008 6974 16017
rect 6918 15943 6974 15952
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15706 6868 15846
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6828 15496 6880 15502
rect 6748 15456 6828 15484
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6748 14822 6776 15456
rect 6828 15438 6880 15444
rect 6920 14952 6972 14958
rect 6840 14900 6920 14906
rect 6840 14894 6972 14900
rect 6840 14878 6960 14894
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14482 6776 14758
rect 6840 14482 6868 14878
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6472 12170 6500 13262
rect 6564 12850 6592 13806
rect 6748 13802 6776 14418
rect 7024 14414 7052 16050
rect 7116 15638 7144 16526
rect 7208 15910 7236 18226
rect 7300 17882 7328 18770
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7116 15094 7144 15574
rect 7300 15162 7328 17070
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7392 14550 7420 19230
rect 7484 18698 7512 20402
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7576 18630 7604 22066
rect 7760 20482 7788 22528
rect 7852 21894 7880 22630
rect 8588 22098 8616 25298
rect 8944 25220 8996 25226
rect 8944 25162 8996 25168
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 8116 20528 8168 20534
rect 7760 20454 7880 20482
rect 8116 20470 8168 20476
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 7668 19514 7696 19926
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7668 18578 7696 19314
rect 7760 18698 7788 20266
rect 7852 19718 7880 20454
rect 8128 19786 8156 20470
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8128 18766 8156 19178
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7472 17672 7524 17678
rect 7470 17640 7472 17649
rect 7524 17640 7526 17649
rect 7470 17575 7526 17584
rect 7576 17270 7604 18566
rect 7668 18550 7788 18578
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16590 7604 17070
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 16182 7604 16390
rect 7564 16176 7616 16182
rect 7564 16118 7616 16124
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7288 14476 7340 14482
rect 7208 14436 7288 14464
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6840 13530 6868 14214
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7208 13326 7236 14436
rect 7288 14418 7340 14424
rect 7392 14414 7420 14486
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7012 13320 7064 13326
rect 6840 13280 7012 13308
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12442 6592 12582
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 11830 6500 12106
rect 6564 11914 6592 12378
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 12050 6684 12174
rect 6840 12050 6868 13280
rect 7012 13262 7064 13268
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6656 12022 6868 12050
rect 6564 11886 6684 11914
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6092 11222 6144 11228
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5736 6798 5764 7414
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5828 6730 5856 7482
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5920 6458 5948 8434
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6012 7886 6040 8366
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6012 6322 6040 7822
rect 6104 7410 6132 11222
rect 6196 11206 6316 11234
rect 6196 11150 6224 11206
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10674 6224 11086
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 10062 6224 10610
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6182 9752 6238 9761
rect 6182 9687 6238 9696
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 6866 6132 7346
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6196 6202 6224 9687
rect 6380 8906 6408 11290
rect 6472 9994 6500 11766
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6564 9586 6592 11562
rect 6656 11121 6684 11886
rect 6748 11830 6776 12022
rect 6932 11898 6960 12650
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 12238 7144 12378
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 7116 11218 7144 12038
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6828 11144 6880 11150
rect 6642 11112 6698 11121
rect 6828 11086 6880 11092
rect 6642 11047 6698 11056
rect 6656 10674 6684 11047
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6656 10266 6684 10610
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6656 10062 6684 10202
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6472 8498 6500 9386
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 7886 6500 8434
rect 6564 8362 6592 9522
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 9042 6684 9454
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 8430 6684 8978
rect 6748 8974 6776 9862
rect 6840 9178 6868 11086
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6748 7954 6776 8910
rect 6840 8634 6868 9114
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6932 8498 6960 11018
rect 7116 10674 7144 11154
rect 7208 11082 7236 12582
rect 7300 12306 7328 13330
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 9110 7052 10474
rect 7116 10062 7144 10610
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 10010 7236 10202
rect 7300 10198 7328 11018
rect 7392 10742 7420 13466
rect 7484 12442 7512 15506
rect 7668 14550 7696 17614
rect 7760 15144 7788 18550
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8312 18408 8340 18770
rect 8220 18380 8340 18408
rect 8220 17678 8248 18380
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8220 16794 8248 17274
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8208 16108 8260 16114
rect 8128 16046 8156 16079
rect 8312 16096 8340 16458
rect 8260 16068 8340 16096
rect 8208 16050 8260 16056
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8128 15366 8156 15982
rect 8312 15502 8340 16068
rect 8404 15706 8432 19246
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8496 18970 8524 19110
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8496 18034 8524 18634
rect 8588 18154 8616 20198
rect 8864 20058 8892 21830
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 18290 8708 19314
rect 8758 18864 8814 18873
rect 8758 18799 8814 18808
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8496 18006 8616 18034
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 17202 8524 17478
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8484 17060 8536 17066
rect 8588 17048 8616 18006
rect 8536 17020 8616 17048
rect 8484 17002 8536 17008
rect 8496 15706 8524 17002
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8668 16584 8720 16590
rect 8772 16572 8800 18799
rect 8864 18698 8892 19994
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8956 18358 8984 25162
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 8720 16544 8800 16572
rect 8668 16526 8720 16532
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8390 15464 8446 15473
rect 8390 15399 8446 15408
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 7760 15116 7880 15144
rect 7852 15026 7880 15116
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 8024 14816 8076 14822
rect 8022 14784 8024 14793
rect 8076 14784 8078 14793
rect 8022 14719 8078 14728
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11218 7512 12174
rect 7576 11762 7604 13262
rect 7668 12986 7696 14350
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8312 14074 8340 14350
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8404 14006 8432 15399
rect 8588 15026 8616 16526
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11642 7604 11698
rect 7576 11614 7696 11642
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11286 7604 11494
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7288 10056 7340 10062
rect 7208 10004 7288 10010
rect 7208 9998 7340 10004
rect 7116 9654 7144 9998
rect 7208 9982 7328 9998
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7208 9382 7236 9982
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 7024 8922 7052 9046
rect 7208 9042 7236 9318
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7024 8894 7236 8922
rect 7300 8906 7328 9862
rect 7392 9722 7420 10066
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7392 8974 7420 9658
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8378 7052 8570
rect 6840 8350 7052 8378
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6840 7886 6868 8350
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 5828 6174 6224 6202
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5460 3602 5488 4014
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3804 3058 3832 3538
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3330 2680 3386 2689
rect 3330 2615 3332 2624
rect 3384 2615 3386 2624
rect 3332 2586 3384 2592
rect 3422 2000 3478 2009
rect 4172 1970 4200 2994
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 5460 2446 5488 3538
rect 5736 3534 5764 5646
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5736 2122 5764 2790
rect 5828 2650 5856 6174
rect 6288 5370 6316 6666
rect 6472 6322 6500 7822
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6196 3398 6224 5034
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6196 2446 6224 3334
rect 6564 2774 6592 7686
rect 6840 6322 6868 7822
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6932 5522 6960 8230
rect 7208 7886 7236 8894
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8634 7328 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7478 7236 7822
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 6798 7052 7278
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7024 6254 7052 6734
rect 7484 6730 7512 10406
rect 7576 10062 7604 11222
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7024 5914 7052 6190
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6840 5494 6960 5522
rect 6840 5234 6868 5494
rect 7024 5234 7052 5850
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3602 6684 3878
rect 6840 3738 6868 5170
rect 7116 4826 7144 5578
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7024 3670 7052 4082
rect 7116 3942 7144 4558
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6472 2746 6592 2774
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5644 2094 5764 2122
rect 3422 1935 3478 1944
rect 4160 1964 4212 1970
rect 3436 1902 3464 1935
rect 4160 1906 4212 1912
rect 5644 1902 5672 2094
rect 5920 1902 5948 2382
rect 6472 2378 6500 2746
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 7392 2106 7420 6326
rect 7576 5642 7604 9658
rect 7668 8480 7696 11614
rect 7760 10810 7788 13874
rect 8312 13841 8340 13874
rect 8298 13832 8354 13841
rect 8298 13767 8354 13776
rect 8496 13326 8524 13874
rect 8484 13320 8536 13326
rect 8404 13268 8484 13274
rect 8404 13262 8536 13268
rect 8404 13246 8524 13262
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 8404 12850 8432 13246
rect 8588 13190 8616 14758
rect 8680 13530 8708 16526
rect 8864 16182 8892 18294
rect 8942 16552 8998 16561
rect 8942 16487 8944 16496
rect 8996 16487 8998 16496
rect 8944 16458 8996 16464
rect 8852 16176 8904 16182
rect 8852 16118 8904 16124
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8496 12782 8524 13126
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8312 12238 8340 12718
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8404 12306 8432 12650
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 8206 11112 8262 11121
rect 8206 11047 8208 11056
rect 8260 11047 8262 11056
rect 8208 11018 8260 11024
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 8496 10742 8524 12582
rect 8588 11014 8616 13126
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8680 12238 8708 12854
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8772 11014 8800 16050
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 9450 7788 10610
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8404 10198 8432 10542
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 8404 9518 8432 10134
rect 8496 9586 8524 10678
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7760 8634 7788 9386
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8492 7800 8498
rect 7668 8452 7748 8480
rect 7748 8434 7800 8440
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8864 7546 8892 15846
rect 8956 15201 8984 16458
rect 9048 16114 9076 23190
rect 9140 21894 9168 28562
rect 9220 25968 9272 25974
rect 9220 25910 9272 25916
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9232 21570 9260 25910
rect 9324 24410 9352 28970
rect 9508 28626 9536 31826
rect 9956 31272 10008 31278
rect 9956 31214 10008 31220
rect 9588 30864 9640 30870
rect 9588 30806 9640 30812
rect 9600 30598 9628 30806
rect 9968 30802 9996 31214
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9968 30258 9996 30738
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 9968 29714 9996 30194
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 10152 29034 10180 32166
rect 10980 31890 11100 31906
rect 10968 31884 11100 31890
rect 11020 31878 11100 31884
rect 10968 31826 11020 31832
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 10244 31482 10272 31622
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 11072 31414 11100 31878
rect 11164 31822 11192 32302
rect 11256 32298 11284 32506
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 11244 32292 11296 32298
rect 11244 32234 11296 32240
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 11256 31498 11284 32234
rect 11369 32124 11677 32133
rect 11369 32122 11375 32124
rect 11431 32122 11455 32124
rect 11511 32122 11535 32124
rect 11591 32122 11615 32124
rect 11671 32122 11677 32124
rect 11431 32070 11433 32122
rect 11613 32070 11615 32122
rect 11369 32068 11375 32070
rect 11431 32068 11455 32070
rect 11511 32068 11535 32070
rect 11591 32068 11615 32070
rect 11671 32068 11677 32070
rect 11369 32059 11677 32068
rect 12544 32026 12572 32370
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 11888 31952 11940 31958
rect 11888 31894 11940 31900
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11164 31482 11284 31498
rect 11152 31476 11284 31482
rect 11204 31470 11284 31476
rect 11152 31418 11204 31424
rect 11060 31408 11112 31414
rect 11060 31350 11112 31356
rect 11072 30802 11100 31350
rect 11164 31346 11192 31418
rect 11152 31340 11204 31346
rect 11152 31282 11204 31288
rect 11532 31278 11560 31758
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 11060 30796 11112 30802
rect 11060 30738 11112 30744
rect 11072 30258 11100 30738
rect 11716 30258 11744 31826
rect 11900 30258 11928 31894
rect 13096 31822 13124 32166
rect 14292 31822 14320 32370
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 13084 31816 13136 31822
rect 13084 31758 13136 31764
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 12164 31680 12216 31686
rect 12164 31622 12216 31628
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11060 30252 11112 30258
rect 11060 30194 11112 30200
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10140 29028 10192 29034
rect 10140 28970 10192 28976
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9404 27396 9456 27402
rect 9404 27338 9456 27344
rect 9416 27130 9444 27338
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9416 24290 9444 27066
rect 9600 26586 9628 28494
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10060 26926 10088 27950
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10048 26920 10100 26926
rect 10048 26862 10100 26868
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9692 25226 9720 26318
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 26042 9812 26182
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9680 25220 9732 25226
rect 9680 25162 9732 25168
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9140 21542 9260 21570
rect 9324 24262 9444 24290
rect 9140 17542 9168 21542
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9126 16824 9182 16833
rect 9126 16759 9182 16768
rect 9140 16726 9168 16759
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9232 15978 9260 21422
rect 9324 20942 9352 24262
rect 9692 22982 9720 24550
rect 9876 23730 9904 26794
rect 9956 26512 10008 26518
rect 9956 26454 10008 26460
rect 9968 24206 9996 26454
rect 10060 26382 10088 26862
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25158 10088 26182
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10152 24818 10180 27270
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 10244 24954 10272 26250
rect 10428 25906 10456 29990
rect 11072 29782 11100 30194
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11060 29776 11112 29782
rect 11060 29718 11112 29724
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10704 29170 10732 29650
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11072 29306 11100 29446
rect 11060 29300 11112 29306
rect 11060 29242 11112 29248
rect 11072 29170 11100 29242
rect 11716 29170 11744 30194
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 10600 27668 10652 27674
rect 10600 27610 10652 27616
rect 10612 27470 10640 27610
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10140 24812 10192 24818
rect 10060 24772 10140 24800
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9784 23186 9812 23666
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 21486 9444 22578
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9324 19378 9352 20402
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18290 9352 18702
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 16697 9352 17546
rect 9416 17184 9444 21422
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9508 20466 9536 21286
rect 9784 20874 9812 22102
rect 9876 21944 9904 23666
rect 9968 23254 9996 24142
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 9968 22098 9996 23054
rect 10060 22166 10088 24772
rect 10140 24754 10192 24760
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10244 24410 10272 24618
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10244 23780 10272 24346
rect 10152 23752 10272 23780
rect 10152 23662 10180 23752
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10428 23186 10456 25366
rect 10980 25158 11008 25842
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10980 24818 11008 25094
rect 11072 24954 11100 28902
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11716 28490 11744 29106
rect 11704 28484 11756 28490
rect 11704 28426 11756 28432
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11716 27130 11744 27950
rect 11808 27674 11836 28358
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11900 27470 11928 29514
rect 11992 27538 12020 31282
rect 12084 31210 12112 31418
rect 12176 31278 12204 31622
rect 12360 31414 12388 31758
rect 13728 31476 13780 31482
rect 13728 31418 13780 31424
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12164 31272 12216 31278
rect 12164 31214 12216 31220
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 12072 31204 12124 31210
rect 12072 31146 12124 31152
rect 12084 30938 12112 31146
rect 12624 31136 12676 31142
rect 12624 31078 12676 31084
rect 12072 30932 12124 30938
rect 12072 30874 12124 30880
rect 12636 30734 12664 31078
rect 13188 30734 13216 31214
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13188 30598 13216 30670
rect 13268 30660 13320 30666
rect 13268 30602 13320 30608
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 12728 30394 12756 30534
rect 12716 30388 12768 30394
rect 12716 30330 12768 30336
rect 12728 29510 12756 30330
rect 13188 30190 13216 30534
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 12900 30116 12952 30122
rect 12900 30058 12952 30064
rect 12912 29782 12940 30058
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 13188 29646 13216 30126
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12360 28558 12388 29038
rect 12728 28966 12756 29446
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12728 28626 12756 28902
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12360 28082 12388 28494
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11704 25220 11756 25226
rect 11704 25162 11756 25168
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10520 24206 10548 24686
rect 10692 24336 10744 24342
rect 10692 24278 10744 24284
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10520 23662 10548 24142
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 10428 22166 10456 23122
rect 10612 23118 10640 23734
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9876 21916 10180 21944
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9600 20262 9628 20810
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9692 20058 9720 20470
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9784 19689 9812 20810
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9876 19922 9904 19994
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9770 19680 9826 19689
rect 9770 19615 9826 19624
rect 9772 19304 9824 19310
rect 9770 19272 9772 19281
rect 9824 19272 9826 19281
rect 9770 19207 9826 19216
rect 9772 19168 9824 19174
rect 9508 19116 9772 19122
rect 9508 19110 9824 19116
rect 9508 19094 9812 19110
rect 9508 18630 9536 19094
rect 9496 18624 9548 18630
rect 9494 18592 9496 18601
rect 9548 18592 9550 18601
rect 9494 18527 9550 18536
rect 9876 18426 9904 19722
rect 9968 19242 9996 20742
rect 10152 19938 10180 21916
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10244 20058 10272 21082
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10230 19952 10286 19961
rect 10152 19910 10230 19938
rect 10230 19887 10286 19896
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10152 19553 10180 19722
rect 10138 19544 10194 19553
rect 10048 19508 10100 19514
rect 10138 19479 10194 19488
rect 10048 19450 10100 19456
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9494 17640 9550 17649
rect 9494 17575 9496 17584
rect 9548 17575 9550 17584
rect 9496 17546 9548 17552
rect 9692 17542 9720 18022
rect 9968 17678 9996 18294
rect 10060 17678 10088 19450
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10152 18630 10180 19382
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 18086 10180 18566
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9496 17196 9548 17202
rect 9416 17156 9496 17184
rect 9496 17138 9548 17144
rect 9600 17082 9628 17478
rect 10060 17338 10088 17614
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9956 17128 10008 17134
rect 9416 17076 9956 17082
rect 9416 17070 10008 17076
rect 9416 17054 9996 17070
rect 9310 16688 9366 16697
rect 9310 16623 9366 16632
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9324 16046 9352 16526
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9416 15892 9444 17054
rect 9586 16824 9642 16833
rect 9586 16759 9642 16768
rect 9600 16726 9628 16759
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9324 15864 9444 15892
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8942 15192 8998 15201
rect 8942 15127 8998 15136
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 13938 8984 14962
rect 9048 14414 9076 15438
rect 9232 14890 9260 15642
rect 9324 15473 9352 15864
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9416 15502 9444 15535
rect 9404 15496 9456 15502
rect 9310 15464 9366 15473
rect 9404 15438 9456 15444
rect 9310 15399 9366 15408
rect 9600 15314 9628 16526
rect 9692 16250 9720 16526
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9692 16153 9720 16186
rect 9678 16144 9734 16153
rect 9784 16114 9812 16662
rect 10060 16114 10088 17274
rect 9678 16079 9734 16088
rect 9772 16108 9824 16114
rect 10048 16108 10100 16114
rect 9824 16068 9996 16096
rect 9772 16050 9824 16056
rect 9416 15286 9628 15314
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9310 14784 9366 14793
rect 9310 14719 9366 14728
rect 9036 14408 9088 14414
rect 9220 14408 9272 14414
rect 9036 14350 9088 14356
rect 9126 14376 9182 14385
rect 9048 13938 9076 14350
rect 9220 14350 9272 14356
rect 9126 14311 9182 14320
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 8974 8984 11086
rect 9048 11082 9076 12786
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 9140 10146 9168 14311
rect 9232 13462 9260 14350
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9324 13258 9352 14719
rect 9416 14396 9444 15286
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9600 14929 9628 14962
rect 9586 14920 9642 14929
rect 9586 14855 9642 14864
rect 9692 14804 9720 14962
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9600 14793 9720 14804
rect 9586 14784 9720 14793
rect 9642 14776 9720 14784
rect 9586 14719 9642 14728
rect 9600 14600 9628 14719
rect 9600 14572 9720 14600
rect 9496 14408 9548 14414
rect 9416 14376 9496 14396
rect 9548 14376 9550 14385
rect 9416 14368 9494 14376
rect 9692 14346 9720 14572
rect 9494 14311 9550 14320
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9232 12646 9260 12922
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 12209 9260 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9218 12200 9274 12209
rect 9218 12135 9274 12144
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 10674 9260 11494
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10266 9260 10406
rect 9324 10266 9352 12242
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9140 10118 9260 10146
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6390 7696 6870
rect 8312 6662 8340 7414
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 8220 5556 8248 6394
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5817 8340 6054
rect 8404 5914 8432 7346
rect 8956 6798 8984 8910
rect 9140 7478 9168 9998
rect 9232 9654 9260 10118
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9232 8430 9260 9590
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9178 9352 9522
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9232 7002 9260 7822
rect 9416 7478 9444 11698
rect 9508 11286 9536 13806
rect 9600 13530 9628 14214
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9680 13320 9732 13326
rect 9678 13288 9680 13297
rect 9772 13320 9824 13326
rect 9732 13288 9734 13297
rect 9772 13262 9824 13268
rect 9678 13223 9734 13232
rect 9634 13184 9686 13190
rect 9784 13172 9812 13262
rect 9686 13144 9812 13172
rect 9634 13126 9686 13132
rect 9678 13016 9734 13025
rect 9678 12951 9734 12960
rect 9586 12880 9642 12889
rect 9586 12815 9588 12824
rect 9640 12815 9642 12824
rect 9588 12786 9640 12792
rect 9692 12434 9720 12951
rect 9876 12782 9904 14826
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9600 12406 9720 12434
rect 9600 11354 9628 12406
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10810 9536 10950
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9600 10674 9628 11290
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 9926 9720 10542
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8956 6322 8984 6734
rect 9232 6322 9260 6938
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8298 5808 8354 5817
rect 8298 5743 8354 5752
rect 8220 5528 8340 5556
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8312 5352 8340 5528
rect 8220 5324 8340 5352
rect 8220 5234 8248 5324
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8220 4536 8248 5170
rect 8680 4622 8708 6054
rect 9128 5772 9180 5778
rect 9232 5760 9260 6258
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9180 5732 9260 5760
rect 9128 5714 9180 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5370 9076 5646
rect 9324 5574 9352 6054
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9402 5536 9458 5545
rect 9402 5471 9458 5480
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8220 4508 8340 4536
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 8312 4282 8340 4508
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8588 4214 8616 4422
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8588 3738 8616 4150
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 9324 3058 9352 3402
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 9324 2106 9352 2994
rect 9416 2650 9444 5471
rect 9508 5370 9536 8026
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9600 5250 9628 8366
rect 9692 7274 9720 9862
rect 9784 9178 9812 12174
rect 9876 12170 9904 12718
rect 9968 12170 9996 16068
rect 10048 16050 10100 16056
rect 10152 16096 10180 17478
rect 10244 16658 10272 19887
rect 10336 17338 10364 20538
rect 10428 20534 10456 22102
rect 10520 20602 10548 22714
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10416 20528 10468 20534
rect 10416 20470 10468 20476
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 20058 10456 20198
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 18970 10456 19654
rect 10520 19514 10548 20334
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10428 18698 10456 18906
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10612 18408 10640 21286
rect 10704 19378 10732 24278
rect 10968 24132 11020 24138
rect 10968 24074 11020 24080
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10888 22234 10916 23054
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10796 19802 10824 19994
rect 10888 19922 10916 20266
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10980 19854 11008 24074
rect 11072 21146 11100 24754
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11716 24274 11744 25162
rect 11808 24818 11836 25978
rect 11900 25498 11928 27406
rect 13004 26994 13032 27814
rect 13188 27470 13216 28018
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 12084 26246 12112 26930
rect 12716 26920 12768 26926
rect 12716 26862 12768 26868
rect 12728 26382 12756 26862
rect 13004 26450 13032 26930
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 12164 26240 12216 26246
rect 12728 26234 12756 26318
rect 12164 26182 12216 26188
rect 12636 26206 12756 26234
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 12084 25226 12112 26182
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11992 24274 12020 24686
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 12084 24206 12112 25162
rect 12176 24886 12204 26182
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12268 25362 12296 25638
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12360 25294 12388 25910
rect 12636 25770 12664 26206
rect 13004 25906 13032 26386
rect 13280 25974 13308 30602
rect 13740 30598 13768 31418
rect 14372 31204 14424 31210
rect 14372 31146 14424 31152
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14016 30734 14044 31078
rect 14384 30802 14412 31146
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13740 30394 13768 30534
rect 13728 30388 13780 30394
rect 13728 30330 13780 30336
rect 14016 30258 14044 30670
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14384 30190 14412 30738
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 13832 29646 13860 30058
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13832 29170 13860 29582
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 14200 29102 14228 29514
rect 14384 29238 14412 30126
rect 14476 29850 14504 32370
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15120 31822 15148 32166
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 15200 31204 15252 31210
rect 15200 31146 15252 31152
rect 15212 30734 15240 31146
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 14464 29844 14516 29850
rect 14464 29786 14516 29792
rect 14844 29714 14872 30194
rect 15212 30122 15240 30670
rect 15200 30116 15252 30122
rect 15200 30058 15252 30064
rect 14832 29708 14884 29714
rect 14832 29650 14884 29656
rect 15212 29646 15240 30058
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 13820 28960 13872 28966
rect 13820 28902 13872 28908
rect 13832 28422 13860 28902
rect 14200 28626 14228 29038
rect 14384 28694 14412 29174
rect 15212 29034 15240 29582
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15764 28762 15792 32370
rect 18315 32124 18623 32133
rect 18315 32122 18321 32124
rect 18377 32122 18401 32124
rect 18457 32122 18481 32124
rect 18537 32122 18561 32124
rect 18617 32122 18623 32124
rect 18377 32070 18379 32122
rect 18559 32070 18561 32122
rect 18315 32068 18321 32070
rect 18377 32068 18401 32070
rect 18457 32068 18481 32070
rect 18537 32068 18561 32070
rect 18617 32068 18623 32070
rect 18315 32059 18623 32068
rect 25261 32124 25569 32133
rect 25261 32122 25267 32124
rect 25323 32122 25347 32124
rect 25403 32122 25427 32124
rect 25483 32122 25507 32124
rect 25563 32122 25569 32124
rect 25323 32070 25325 32122
rect 25505 32070 25507 32122
rect 25261 32068 25267 32070
rect 25323 32068 25347 32070
rect 25403 32068 25427 32070
rect 25483 32068 25507 32070
rect 25563 32068 25569 32070
rect 25261 32059 25569 32068
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16408 29306 16436 31758
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 14372 28688 14424 28694
rect 14372 28630 14424 28636
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13728 27940 13780 27946
rect 13728 27882 13780 27888
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13556 26586 13584 27066
rect 13740 26994 13768 27882
rect 13832 27130 13860 28358
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 13820 27124 13872 27130
rect 13820 27066 13872 27072
rect 14384 26994 14412 27270
rect 14476 27130 14504 27270
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13556 26042 13584 26522
rect 13544 26036 13596 26042
rect 13544 25978 13596 25984
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12268 24206 12296 24754
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11164 21894 11192 23666
rect 12268 23662 12296 24142
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11716 22778 11744 23258
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22438 11744 22578
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10968 19848 11020 19854
rect 10796 19774 10916 19802
rect 10968 19790 11020 19796
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10520 18380 10640 18408
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10428 17814 10456 18226
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10336 16250 10364 16730
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16108 10284 16114
rect 10152 16068 10232 16096
rect 10152 15706 10180 16068
rect 10232 16050 10284 16056
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10060 15026 10088 15642
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10152 12714 10180 15642
rect 10244 15434 10272 15846
rect 10336 15570 10364 16186
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10244 14890 10272 15370
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10230 14512 10286 14521
rect 10230 14447 10286 14456
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11354 9904 11494
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9876 10674 9904 11290
rect 9968 11218 9996 12106
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11898 10180 12038
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9876 10062 9904 10610
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9876 6662 9904 8774
rect 10152 7002 10180 10066
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10046 6896 10102 6905
rect 10046 6831 10102 6840
rect 10060 6798 10088 6831
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9508 5222 9628 5250
rect 9864 5228 9916 5234
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 3424 1896 3476 1902
rect 3424 1838 3476 1844
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 4423 1660 4731 1669
rect 4423 1658 4429 1660
rect 4485 1658 4509 1660
rect 4565 1658 4589 1660
rect 4645 1658 4669 1660
rect 4725 1658 4731 1660
rect 4485 1606 4487 1658
rect 4667 1606 4669 1658
rect 4423 1604 4429 1606
rect 4485 1604 4509 1606
rect 4565 1604 4589 1606
rect 4645 1604 4669 1606
rect 4725 1604 4731 1606
rect 4423 1595 4731 1604
rect 5644 1562 5672 1838
rect 8208 1760 8260 1766
rect 8260 1708 8340 1714
rect 8208 1702 8340 1708
rect 8220 1686 8340 1702
rect 5632 1556 5684 1562
rect 5632 1498 5684 1504
rect 1952 1420 2004 1426
rect 1952 1362 2004 1368
rect 8312 1358 8340 1686
rect 9416 1358 9444 2586
rect 8300 1352 8352 1358
rect 3330 1320 3386 1329
rect 2228 1284 2280 1290
rect 8300 1294 8352 1300
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9508 1290 9536 5222
rect 9916 5188 9996 5216
rect 9864 5170 9916 5176
rect 9968 4622 9996 5188
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 2038 9628 3946
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 2514 9904 2994
rect 10244 2774 10272 14447
rect 10336 12442 10364 15506
rect 10428 15502 10456 15914
rect 10520 15570 10548 18380
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15026 10548 15302
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10428 14618 10456 14962
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10520 14498 10548 14758
rect 10612 14618 10640 18226
rect 10704 16590 10732 18226
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10704 16114 10732 16186
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10796 15162 10824 19450
rect 10888 19378 10916 19774
rect 11072 19553 11100 20334
rect 11058 19544 11114 19553
rect 11164 19530 11192 20878
rect 11256 19854 11284 22170
rect 11716 22094 11744 22374
rect 11716 22066 11928 22094
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11716 20874 11744 21490
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11624 20754 11652 20810
rect 11796 20800 11848 20806
rect 11624 20726 11744 20754
rect 11796 20742 11848 20748
rect 11612 20392 11664 20398
rect 11610 20360 11612 20369
rect 11664 20360 11666 20369
rect 11610 20295 11666 20304
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11244 19848 11296 19854
rect 11242 19816 11244 19825
rect 11296 19816 11298 19825
rect 11440 19786 11468 19887
rect 11242 19751 11298 19760
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11336 19712 11388 19718
rect 11334 19680 11336 19689
rect 11388 19680 11390 19689
rect 11334 19615 11390 19624
rect 11164 19502 11284 19530
rect 11058 19479 11114 19488
rect 11256 19446 11284 19502
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 17882 10916 18566
rect 10980 18290 11008 18838
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15609 10916 15982
rect 10874 15600 10930 15609
rect 10874 15535 10930 15544
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10520 14470 10640 14498
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13258 10548 14214
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 12102 10364 12378
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10428 11778 10456 12174
rect 10336 11762 10456 11778
rect 10324 11756 10456 11762
rect 10376 11750 10456 11756
rect 10324 11698 10376 11704
rect 10428 11218 10456 11750
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 11014 10456 11154
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10336 10810 10364 10950
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10336 10470 10364 10610
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10130 10364 10406
rect 10612 10266 10640 14470
rect 10796 14346 10824 14962
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10796 13938 10824 14282
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13530 10916 15438
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10704 12306 10732 13466
rect 10980 13410 11008 17206
rect 11072 16232 11100 19382
rect 11256 18766 11284 19382
rect 11532 19174 11560 19722
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11164 16794 11192 17614
rect 11256 16998 11284 18702
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11716 17066 11744 20726
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11072 16204 11284 16232
rect 11150 16144 11206 16153
rect 11150 16079 11206 16088
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 14550 11100 15370
rect 11164 15026 11192 16079
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11060 14544 11112 14550
rect 11256 14498 11284 16204
rect 11348 16114 11376 16730
rect 11716 16697 11744 17002
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11808 16590 11836 20742
rect 11900 19378 11928 22066
rect 11992 20398 12020 23258
rect 12084 22642 12112 23462
rect 12360 23322 12388 25230
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12452 24886 12480 25162
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12360 23118 12388 23258
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 20262 12020 20334
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 17270 11928 19178
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11624 15337 11652 15438
rect 11704 15360 11756 15366
rect 11610 15328 11666 15337
rect 11704 15302 11756 15308
rect 11610 15263 11666 15272
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11060 14486 11112 14492
rect 11164 14470 11468 14498
rect 11164 14396 11192 14470
rect 11440 14414 11468 14470
rect 10796 13382 11008 13410
rect 11072 14368 11192 14396
rect 11244 14408 11296 14414
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11354 10732 11630
rect 10796 11558 10824 13382
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12374 10916 13126
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10980 12442 11008 12854
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10336 8294 10364 10066
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9722 10456 9998
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10704 9382 10732 9658
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10336 7206 10364 8230
rect 10428 7410 10456 8230
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 4690 10456 6258
rect 10520 6225 10548 8502
rect 10704 7886 10732 9318
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 6390 10640 7686
rect 10796 7562 10824 8842
rect 10704 7534 10824 7562
rect 11072 7562 11100 14368
rect 11244 14350 11296 14356
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11164 12238 11192 13806
rect 11256 13462 11284 14350
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13938 11652 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11256 12374 11284 13262
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12850 11652 13126
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11354 11192 12038
rect 11244 11552 11296 11558
rect 11624 11540 11652 12378
rect 11716 12238 11744 15302
rect 11808 14521 11836 16390
rect 11900 15162 11928 16458
rect 11992 16250 12020 16934
rect 12084 16454 12112 21898
rect 12176 20602 12204 22578
rect 12452 21894 12480 24822
rect 12636 24138 12664 25706
rect 12728 24614 12756 25842
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13188 24857 13216 25162
rect 13174 24848 13230 24857
rect 13174 24783 13230 24792
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12268 20398 12296 21490
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12176 19689 12204 20334
rect 12162 19680 12218 19689
rect 12162 19615 12218 19624
rect 12268 19446 12296 20334
rect 12360 19786 12388 21082
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 12346 19544 12402 19553
rect 12346 19479 12402 19488
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12268 17202 12296 17682
rect 12360 17610 12388 19479
rect 12452 17882 12480 19926
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 17202 12388 17546
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12268 17082 12296 17138
rect 12268 17054 12388 17082
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15434 12020 16186
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 11888 14544 11940 14550
rect 11794 14512 11850 14521
rect 11888 14486 11940 14492
rect 11794 14447 11850 14456
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11898 11744 12174
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11808 11762 11836 14010
rect 11900 14006 11928 14486
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11900 13274 11928 13942
rect 11900 13246 12112 13274
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11624 11512 11744 11540
rect 11244 11494 11296 11500
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10130 11192 10950
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9586 11192 10066
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11164 8498 11192 9522
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11072 7534 11192 7562
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10506 6216 10562 6225
rect 10506 6151 10562 6160
rect 10520 5914 10548 6151
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10428 4214 10456 4626
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10520 3670 10548 4422
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10244 2746 10364 2774
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9588 2032 9640 2038
rect 9588 1974 9640 1980
rect 9876 1970 9904 2450
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 3330 1255 3386 1264
rect 9496 1284 9548 1290
rect 2228 1226 2280 1232
rect 2240 921 2268 1226
rect 3344 1222 3372 1255
rect 9496 1226 9548 1232
rect 10336 1222 10364 2746
rect 10520 1222 10548 3606
rect 10704 3602 10732 7534
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 4826 10824 7278
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 6934 10916 7142
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10796 2774 10824 4762
rect 11072 4706 11100 6054
rect 10980 4678 11100 4706
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4146 10916 4558
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10888 3602 10916 4082
rect 10980 4078 11008 4678
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10888 3058 10916 3538
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2802 11008 4014
rect 11072 3194 11100 4490
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11072 2922 11100 3130
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10980 2774 11100 2802
rect 10796 2746 10916 2774
rect 10888 2446 10916 2746
rect 11072 2446 11100 2774
rect 11164 2774 11192 7534
rect 11256 5710 11284 11494
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11716 10962 11744 11512
rect 11624 10934 11744 10962
rect 11624 10674 11652 10934
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11716 9466 11744 10746
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11808 9586 11836 9930
rect 11900 9586 11928 12582
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11992 12238 12020 12310
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11716 9438 11836 9466
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11716 5642 11744 9046
rect 11808 9042 11836 9438
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 8378 11836 8978
rect 11900 8974 11928 9522
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11992 8838 12020 12038
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11808 8350 11928 8378
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11808 6798 11836 7958
rect 11900 7721 11928 8350
rect 11886 7712 11942 7721
rect 11886 7647 11942 7656
rect 12084 6934 12112 13246
rect 12176 12986 12204 14962
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12268 12434 12296 16594
rect 12360 16182 12388 17054
rect 12544 16726 12572 23258
rect 12728 20534 12756 24550
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13280 23118 13308 24142
rect 14568 23730 14596 27950
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 25265 15884 25638
rect 15842 25256 15898 25265
rect 15842 25191 15898 25200
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14830 24848 14886 24857
rect 14740 24812 14792 24818
rect 14830 24783 14832 24792
rect 14740 24754 14792 24760
rect 14884 24783 14886 24792
rect 14832 24754 14884 24760
rect 14752 23798 14780 24754
rect 16040 24750 16068 25842
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14740 23792 14792 23798
rect 14740 23734 14792 23740
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22098 12848 22918
rect 12912 22642 12940 22986
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 13004 19378 13032 20878
rect 13280 19718 13308 23054
rect 14568 23050 14596 23666
rect 15580 23526 15608 24686
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13372 22778 13400 22918
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13728 22704 13780 22710
rect 13780 22652 13952 22658
rect 13728 22646 13952 22652
rect 13740 22630 13952 22646
rect 13924 22506 13952 22630
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13648 19378 13676 21626
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 12992 19372 13044 19378
rect 13636 19372 13688 19378
rect 13044 19332 13124 19360
rect 12992 19314 13044 19320
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12636 17678 12664 18362
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12728 17338 12756 18158
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14074 12388 15506
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12452 13433 12480 13874
rect 12636 13716 12664 15846
rect 12716 14272 12768 14278
rect 12714 14240 12716 14249
rect 12768 14240 12770 14249
rect 12714 14175 12770 14184
rect 12820 14074 12848 18702
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12912 17678 12940 18634
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12898 17504 12954 17513
rect 12898 17439 12954 17448
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12636 13688 12756 13716
rect 12438 13424 12494 13433
rect 12438 13359 12494 13368
rect 12176 12406 12296 12434
rect 12176 8906 12204 12406
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12268 9518 12296 11222
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11900 4026 11928 6666
rect 12176 6662 12204 8502
rect 12268 7546 12296 9454
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12268 6390 12296 6802
rect 12360 6662 12388 11290
rect 12452 8634 12480 13359
rect 12728 12918 12756 13688
rect 12912 13462 12940 17439
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12544 8945 12572 9590
rect 12636 8974 12664 12650
rect 12728 8974 12756 12854
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12209 12848 12786
rect 12806 12200 12862 12209
rect 12806 12135 12862 12144
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12624 8968 12676 8974
rect 12530 8936 12586 8945
rect 12624 8910 12676 8916
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12530 8871 12586 8880
rect 12440 8628 12492 8634
rect 12544 8616 12572 8871
rect 12544 8588 12664 8616
rect 12440 8570 12492 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 7954 12572 8434
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12438 7712 12494 7721
rect 12438 7647 12494 7656
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5302 12112 5646
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12176 4593 12204 5578
rect 12360 5370 12388 6258
rect 12452 5778 12480 7647
rect 12636 7410 12664 8588
rect 12820 7886 12848 11494
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 9994 12940 10610
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12912 9586 12940 9930
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8022 12940 8774
rect 13004 8498 13032 19178
rect 13096 18426 13124 19332
rect 13636 19314 13688 19320
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13464 17746 13492 18022
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13188 17202 13216 17546
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13648 15994 13676 19314
rect 13726 19272 13782 19281
rect 13726 19207 13782 19216
rect 13740 16182 13768 19207
rect 13832 18358 13860 20742
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13924 18630 13952 20470
rect 14016 19514 14044 21286
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14016 18698 14044 18906
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13648 15966 13768 15994
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13096 11558 13124 15030
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13280 13394 13308 13738
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13372 13190 13400 15574
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14074 13676 14826
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12850 13400 13126
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13464 12714 13492 14010
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13556 13870 13584 13942
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13266 12200 13322 12209
rect 13266 12135 13322 12144
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5370 12572 6666
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12162 4584 12218 4593
rect 12162 4519 12218 4528
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11808 4010 11928 4026
rect 11796 4004 11928 4010
rect 11848 3998 11928 4004
rect 11796 3946 11848 3952
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11716 3126 11744 3878
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11992 3058 12020 4082
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11164 2746 11284 2774
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11256 2038 11284 2746
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 12084 2650 12112 3606
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12176 2038 12204 4519
rect 12268 3942 12296 5170
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12268 2514 12296 2586
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 11244 2032 11296 2038
rect 11244 1974 11296 1980
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11369 1660 11677 1669
rect 11369 1658 11375 1660
rect 11431 1658 11455 1660
rect 11511 1658 11535 1660
rect 11591 1658 11615 1660
rect 11671 1658 11677 1660
rect 11431 1606 11433 1658
rect 11613 1606 11615 1658
rect 11369 1604 11375 1606
rect 11431 1604 11455 1606
rect 11511 1604 11535 1606
rect 11591 1604 11615 1606
rect 11671 1604 11677 1606
rect 11369 1595 11677 1604
rect 11900 1562 11928 1702
rect 11888 1556 11940 1562
rect 11888 1498 11940 1504
rect 11980 1352 12032 1358
rect 11978 1320 11980 1329
rect 12032 1320 12034 1329
rect 12360 1290 12388 5306
rect 12440 5296 12492 5302
rect 12438 5264 12440 5273
rect 12492 5264 12494 5273
rect 12636 5234 12664 7346
rect 12820 6882 12848 7346
rect 12728 6854 12848 6882
rect 12728 6730 12756 6854
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12820 5846 12848 6734
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12438 5199 12494 5208
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12728 5114 12756 5510
rect 12452 5086 12756 5114
rect 12452 2446 12480 5086
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12452 1465 12480 2382
rect 12544 1970 12572 4762
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12636 3398 12664 4490
rect 12820 3448 12848 5782
rect 12912 5273 12940 7958
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 5681 13032 7822
rect 13280 7478 13308 12135
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 8022 13400 9522
rect 13464 9110 13492 11290
rect 13556 9110 13584 13806
rect 13740 13734 13768 15966
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 14550 13860 15846
rect 13924 14822 13952 18566
rect 14016 17542 14044 18634
rect 14108 18358 14136 22374
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21554 14228 21830
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14200 21010 14228 21490
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 17270 14044 17478
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14016 15366 14044 17206
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13832 13546 13860 14214
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13740 13518 13860 13546
rect 13740 13462 13768 13518
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13832 12986 13860 13398
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12646 13768 12786
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13818 12608 13874 12617
rect 13648 9217 13676 12582
rect 13818 12543 13874 12552
rect 13726 10568 13782 10577
rect 13726 10503 13782 10512
rect 13740 10198 13768 10503
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13634 9208 13690 9217
rect 13634 9143 13690 9152
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8362 13492 8774
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13464 7800 13492 8298
rect 13372 7772 13492 7800
rect 13084 7472 13136 7478
rect 13082 7440 13084 7449
rect 13268 7472 13320 7478
rect 13136 7440 13138 7449
rect 13082 7375 13138 7384
rect 13188 7432 13268 7460
rect 13188 5710 13216 7432
rect 13268 7414 13320 7420
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13176 5704 13228 5710
rect 12990 5672 13046 5681
rect 13176 5646 13228 5652
rect 12990 5607 13046 5616
rect 12898 5264 12954 5273
rect 13082 5264 13138 5273
rect 12898 5199 12954 5208
rect 12992 5228 13044 5234
rect 13280 5234 13308 5782
rect 13372 5710 13400 7772
rect 13556 7410 13584 9046
rect 13740 8634 13768 9998
rect 13832 9654 13860 12543
rect 13924 12434 13952 13670
rect 14108 13530 14136 18294
rect 14200 17882 14228 20402
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14200 17338 14228 17546
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14200 15502 14228 17274
rect 14292 16998 14320 18702
rect 14568 18290 14596 22986
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15580 21554 15608 23462
rect 16040 22778 16068 23462
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15672 21418 15700 21966
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14660 18086 14688 18838
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14372 17536 14424 17542
rect 14370 17504 14372 17513
rect 14424 17504 14426 17513
rect 14370 17439 14426 17448
rect 14476 17134 14504 17614
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14200 14346 14228 15438
rect 14292 15434 14320 16934
rect 14384 15638 14412 17002
rect 14476 16114 14504 17070
rect 14568 16980 14596 17614
rect 14660 17134 14688 18022
rect 14752 17338 14780 18566
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 15304 17649 15332 21354
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20754 15608 20810
rect 15488 20726 15608 20754
rect 15488 20262 15516 20726
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 18272 15424 18702
rect 15488 18426 15516 20198
rect 15580 19786 15608 20402
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15580 19446 15608 19722
rect 15672 19718 15700 20334
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15672 19514 15700 19654
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15476 18284 15528 18290
rect 15396 18244 15476 18272
rect 15290 17640 15346 17649
rect 15290 17575 15346 17584
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14752 16980 14780 17138
rect 14568 16952 14780 16980
rect 14568 16182 14596 16952
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14752 16250 14780 16594
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14292 14482 14320 15370
rect 14384 14482 14412 15574
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14200 13326 14228 14282
rect 14292 13938 14320 14418
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14292 13802 14320 13874
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14384 13172 14412 14282
rect 14568 14278 14596 15302
rect 14556 14272 14608 14278
rect 14476 14232 14556 14260
rect 14476 13870 14504 14232
rect 14556 14214 14608 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14462 13560 14518 13569
rect 14462 13495 14518 13504
rect 14476 13190 14504 13495
rect 14200 13144 14412 13172
rect 14464 13184 14516 13190
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12442 14136 12718
rect 14096 12436 14148 12442
rect 13924 12406 14044 12434
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 10810 13952 11630
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 9722 13952 10610
rect 14016 10606 14044 12406
rect 14096 12378 14148 12384
rect 14200 11898 14228 13144
rect 14464 13126 14516 13132
rect 14476 13002 14504 13126
rect 14384 12974 14504 13002
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14096 11756 14148 11762
rect 14148 11716 14228 11744
rect 14096 11698 14148 11704
rect 14094 11656 14150 11665
rect 14094 11591 14150 11600
rect 14108 11150 14136 11591
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 14016 9058 14044 10367
rect 13832 9030 14044 9058
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8288 13688 8294
rect 13832 8242 13860 9030
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14016 8498 14044 8910
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13688 8236 13860 8242
rect 13636 8230 13860 8236
rect 13648 8214 13860 8230
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13082 5199 13138 5208
rect 13268 5228 13320 5234
rect 12992 5170 13044 5176
rect 12900 3460 12952 3466
rect 12820 3420 12900 3448
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12636 2038 12664 3130
rect 12820 2650 12848 3420
rect 12900 3402 12952 3408
rect 13004 3097 13032 5170
rect 13096 3890 13124 5199
rect 13268 5170 13320 5176
rect 13280 4826 13308 5170
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13280 4078 13308 4762
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13096 3862 13216 3890
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12990 3088 13046 3097
rect 12990 3023 13046 3032
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13096 2446 13124 3674
rect 13188 3534 13216 3862
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 2446 13216 3470
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13372 2446 13400 3402
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12532 1964 12584 1970
rect 12532 1906 12584 1912
rect 12438 1456 12494 1465
rect 13096 1426 13124 2246
rect 13464 2038 13492 6938
rect 13726 6896 13782 6905
rect 13726 6831 13782 6840
rect 13740 6662 13768 6831
rect 13544 6656 13596 6662
rect 13728 6656 13780 6662
rect 13596 6616 13676 6644
rect 13544 6598 13596 6604
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5914 13584 6258
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5710 13676 6616
rect 13728 6598 13780 6604
rect 13924 5846 13952 7822
rect 14016 7154 14044 8434
rect 14108 7274 14136 10474
rect 14200 10470 14228 11716
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14292 10130 14320 12174
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14384 9466 14412 12974
rect 14480 9988 14532 9994
rect 14292 9450 14412 9466
rect 14280 9444 14412 9450
rect 14332 9438 14412 9444
rect 14476 9936 14480 9976
rect 14476 9930 14532 9936
rect 14280 9386 14332 9392
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14292 7410 14320 8191
rect 14384 7886 14412 9318
rect 14476 8906 14504 9930
rect 14568 8974 14596 14010
rect 14660 13462 14688 16050
rect 14752 15026 14780 16186
rect 15396 16114 15424 18244
rect 15476 18226 15528 18232
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14752 13988 14780 14418
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 14832 14000 14884 14006
rect 14752 13960 14832 13988
rect 14832 13942 14884 13948
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14752 13258 14780 13806
rect 14844 13326 14872 13806
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 15028 13190 15056 13738
rect 15396 13569 15424 16050
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15580 15026 15608 15438
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15474 13832 15530 13841
rect 15474 13767 15530 13776
rect 15382 13560 15438 13569
rect 15382 13495 15438 13504
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15488 13138 15516 13767
rect 15580 13734 15608 14962
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15580 13258 15608 13670
rect 15672 13569 15700 16390
rect 15764 15910 15792 22374
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 20777 15884 21422
rect 15842 20768 15898 20777
rect 15842 20703 15898 20712
rect 15948 20330 15976 21490
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 16040 18970 16068 22714
rect 16132 20602 16160 24074
rect 16316 23730 16344 27814
rect 17604 26586 17632 28018
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 18340 26994 18368 27406
rect 20260 27396 20312 27402
rect 20260 27338 20312 27344
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 16488 24812 16540 24818
rect 16488 24754 16540 24760
rect 16500 24206 16528 24754
rect 16592 24410 16620 25910
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17236 24818 17264 25842
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 17052 24206 17080 24754
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16224 20806 16252 21490
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16132 19174 16160 20538
rect 16224 19514 16252 20742
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 16120 18828 16172 18834
rect 16040 18788 16120 18816
rect 16040 18358 16068 18788
rect 16120 18770 16172 18776
rect 16316 18698 16344 23666
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 19786 16436 20198
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15856 15706 15884 16458
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15764 14006 15792 15030
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15658 13560 15714 13569
rect 15658 13495 15714 13504
rect 15764 13326 15792 13942
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 14660 9110 14688 13126
rect 15488 13110 15608 13138
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 10554 14780 11834
rect 15200 11824 15252 11830
rect 15014 11792 15070 11801
rect 14832 11756 14884 11762
rect 15200 11766 15252 11772
rect 15014 11727 15016 11736
rect 14832 11698 14884 11704
rect 15068 11727 15070 11736
rect 15016 11698 15068 11704
rect 14844 11150 14872 11698
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14936 11014 14964 11562
rect 15212 11354 15240 11766
rect 15304 11762 15332 12038
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15304 11665 15332 11698
rect 15290 11656 15346 11665
rect 15290 11591 15346 11600
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 14752 10526 14872 10554
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9602 14780 10406
rect 14844 9994 14872 10526
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 14752 9574 15148 9602
rect 15120 9110 15148 9574
rect 15212 9178 15240 9658
rect 15304 9382 15332 11154
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14372 7880 14424 7886
rect 14424 7840 14504 7868
rect 14372 7822 14424 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14016 7126 14136 7154
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5846 14044 6054
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13740 4214 13768 5714
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13728 4208 13780 4214
rect 13648 4168 13728 4196
rect 13648 2106 13676 4168
rect 13728 4150 13780 4156
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3194 13768 3878
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13832 2650 13860 5170
rect 13924 4214 13952 5646
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 14016 3602 14044 5578
rect 14108 4554 14136 7126
rect 14200 6118 14228 7278
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14292 7002 14320 7142
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 6934 14412 7142
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14476 6390 14504 7840
rect 14554 7168 14610 7177
rect 14554 7103 14610 7112
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14568 6322 14596 7103
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14660 6202 14688 8842
rect 14476 6174 14688 6202
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14292 5302 14320 5850
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14292 4826 14320 5238
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14016 2106 14044 3538
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 14004 2100 14056 2106
rect 14004 2042 14056 2048
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 14108 1494 14136 3878
rect 14476 3670 14504 6174
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14568 3058 14596 4966
rect 14660 4826 14688 5782
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14660 4214 14688 4762
rect 14752 4758 14780 8978
rect 15292 8968 15344 8974
rect 15290 8936 15292 8945
rect 15344 8936 15346 8945
rect 15290 8871 15346 8880
rect 15396 8838 15424 11086
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15488 10810 15516 11018
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15488 9450 15516 9522
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 15580 7886 15608 13110
rect 15658 12880 15714 12889
rect 15856 12850 15884 15642
rect 15948 14346 15976 18022
rect 16040 17542 16068 18294
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16132 17134 16160 18634
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16132 16658 16160 17070
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 15162 16160 15302
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16132 14906 16160 15098
rect 16040 14878 16160 14906
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 13297 15976 14282
rect 15934 13288 15990 13297
rect 15934 13223 15990 13232
rect 16040 13190 16068 14878
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16132 13433 16160 13466
rect 16118 13424 16174 13433
rect 16118 13359 16174 13368
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15658 12815 15660 12824
rect 15712 12815 15714 12824
rect 15844 12844 15896 12850
rect 15660 12786 15712 12792
rect 15844 12786 15896 12792
rect 15934 11792 15990 11801
rect 15660 11756 15712 11762
rect 15934 11727 15990 11736
rect 15660 11698 15712 11704
rect 15672 10674 15700 11698
rect 15948 11694 15976 11727
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 10674 15976 11630
rect 16040 10674 16068 13126
rect 16224 12918 16252 18090
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16316 16454 16344 16487
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 13938 16344 15438
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 10810 16160 12786
rect 16224 12306 16252 12854
rect 16316 12850 16344 13874
rect 16408 13734 16436 19722
rect 16500 18986 16528 21082
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20398 16804 20878
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16776 19922 16804 20334
rect 17420 20058 17448 26250
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16776 19666 16804 19858
rect 16776 19638 16896 19666
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16500 18958 16620 18986
rect 16592 18834 16620 18958
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16592 18154 16620 18634
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16684 18034 16712 18634
rect 16592 18006 16712 18034
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 14634 16528 17546
rect 16592 15094 16620 18006
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 15638 16712 17478
rect 16776 15706 16804 19450
rect 16868 17678 16896 19638
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16960 17542 16988 19314
rect 17052 17814 17080 19314
rect 17144 18290 17172 19994
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17236 19310 17264 19382
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18698 17264 19246
rect 17604 18698 17632 26522
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18340 26246 18368 26318
rect 19168 26246 19196 26930
rect 20272 26790 20300 27338
rect 20732 27062 20760 27406
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 17684 26240 17736 26246
rect 17684 26182 17736 26188
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 19156 26240 19208 26246
rect 19156 26182 19208 26188
rect 17696 25498 17724 26182
rect 18340 25906 18368 26182
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18340 25786 18368 25842
rect 18248 25758 18368 25786
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 18248 23118 18276 25758
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17972 22778 18000 22986
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 18156 21962 18184 22918
rect 18248 22030 18276 23054
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17788 21690 17816 21830
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 17052 17202 17080 17750
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16672 15632 16724 15638
rect 16868 15586 16896 16526
rect 16672 15574 16724 15580
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16684 15026 16712 15574
rect 16776 15558 16896 15586
rect 16776 15094 16804 15558
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16776 14958 16804 15030
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16500 14618 16620 14634
rect 16500 14612 16632 14618
rect 16500 14606 16580 14612
rect 16580 14554 16632 14560
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16394 13560 16450 13569
rect 16394 13495 16450 13504
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16224 11830 16252 12242
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16224 11150 16252 11766
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15658 9072 15714 9081
rect 15658 9007 15714 9016
rect 15672 8498 15700 9007
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15292 7336 15344 7342
rect 15014 7304 15070 7313
rect 15292 7278 15344 7284
rect 15014 7239 15070 7248
rect 15200 7268 15252 7274
rect 15028 6798 15056 7239
rect 15200 7210 15252 7216
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14830 6352 14886 6361
rect 14830 6287 14886 6296
rect 14924 6316 14976 6322
rect 14844 5710 14872 6287
rect 14924 6258 14976 6264
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14936 6225 14964 6258
rect 14922 6216 14978 6225
rect 14922 6151 14978 6160
rect 15028 6089 15056 6258
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15014 6080 15070 6089
rect 15014 6015 15070 6024
rect 15120 5914 15148 6122
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15014 5808 15070 5817
rect 15014 5743 15070 5752
rect 15028 5710 15056 5743
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 15212 5370 15240 7210
rect 15304 6458 15332 7278
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15304 5710 15332 6258
rect 15396 5914 15424 7414
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15304 5302 15332 5646
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14752 2990 14780 3470
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14844 3058 14872 3130
rect 15212 3126 15240 3334
rect 15304 3194 15332 5238
rect 15396 3738 15424 5714
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3120 15252 3126
rect 15014 3088 15070 3097
rect 14832 3052 14884 3058
rect 15200 3062 15252 3068
rect 15014 3023 15016 3032
rect 14832 2994 14884 3000
rect 15068 3023 15070 3032
rect 15016 2994 15068 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14752 2514 14780 2926
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14648 2440 14700 2446
rect 14844 2394 14872 2994
rect 14700 2388 14872 2394
rect 14648 2382 14872 2388
rect 14660 2366 14872 2382
rect 15292 2372 15344 2378
rect 14556 1760 14608 1766
rect 14556 1702 14608 1708
rect 14568 1562 14596 1702
rect 14556 1556 14608 1562
rect 14556 1498 14608 1504
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 12438 1391 12494 1400
rect 13084 1420 13136 1426
rect 13084 1362 13136 1368
rect 11978 1255 12034 1264
rect 12348 1284 12400 1290
rect 12348 1226 12400 1232
rect 14752 1222 14780 2366
rect 15292 2314 15344 2320
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 15304 2106 15332 2314
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15488 1358 15516 7346
rect 15580 7002 15608 7686
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15672 6458 15700 8230
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15580 4078 15608 4558
rect 15672 4214 15700 6190
rect 15764 5234 15792 7686
rect 15856 7449 15884 10610
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16040 7546 16068 9590
rect 16132 8634 16160 9998
rect 16224 9110 16252 10950
rect 16316 9450 16344 12582
rect 16408 12442 16436 13495
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11694 16528 12106
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16486 11248 16542 11257
rect 16486 11183 16542 11192
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15842 7440 15898 7449
rect 15842 7375 15898 7384
rect 16132 6934 16160 7822
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16224 6866 16252 8298
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 15844 6792 15896 6798
rect 15842 6760 15844 6769
rect 15896 6760 15898 6769
rect 15842 6695 15898 6704
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 5846 15976 6598
rect 16224 6322 16252 6802
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15856 4282 15884 4558
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15672 1766 15700 2926
rect 15764 2854 15792 2994
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15764 1358 15792 1974
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 15752 1352 15804 1358
rect 15752 1294 15804 1300
rect 15948 1290 15976 5782
rect 16224 5030 16252 6122
rect 16316 5166 16344 9046
rect 16408 7886 16436 10746
rect 16500 8974 16528 11183
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 6458 16436 7822
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 1358 16068 3334
rect 16224 2582 16252 3402
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16316 2038 16344 3334
rect 16408 2854 16436 4966
rect 16500 3194 16528 8774
rect 16592 8022 16620 14554
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 13977 16712 14350
rect 16776 14278 16804 14418
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16670 13968 16726 13977
rect 16670 13903 16726 13912
rect 16684 12374 16712 13903
rect 16868 13530 16896 15438
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 14074 16988 14758
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12782 16896 13262
rect 16946 13152 17002 13161
rect 16946 13087 17002 13096
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16960 12442 16988 13087
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 10441 16712 12038
rect 16776 11150 16804 12378
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11144 16816 11150
rect 16868 11121 16896 11698
rect 16960 11558 16988 12106
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16948 11144 17000 11150
rect 16764 11086 16816 11092
rect 16854 11112 16910 11121
rect 16948 11086 17000 11092
rect 16854 11047 16910 11056
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10674 16896 10950
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16670 10432 16726 10441
rect 16670 10367 16726 10376
rect 16670 10024 16726 10033
rect 16670 9959 16726 9968
rect 16764 9988 16816 9994
rect 16684 9586 16712 9959
rect 16764 9930 16816 9936
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16684 6866 16712 9318
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16776 6798 16804 9930
rect 16960 9178 16988 11086
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16868 8634 16896 9114
rect 16946 9072 17002 9081
rect 16946 9007 17002 9016
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16960 6798 16988 9007
rect 17052 7546 17080 14214
rect 17144 12442 17172 16730
rect 17236 16726 17264 16934
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17328 16454 17356 18226
rect 17420 18154 17448 18634
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17236 13802 17264 15982
rect 17328 15502 17356 16390
rect 17420 15570 17448 17478
rect 17512 15706 17540 18566
rect 17972 18290 18000 18838
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17684 18080 17736 18086
rect 17960 18080 18012 18086
rect 17684 18022 17736 18028
rect 17958 18048 17960 18057
rect 18012 18048 18014 18057
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 13841 17356 15438
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17314 13832 17370 13841
rect 17224 13796 17276 13802
rect 17314 13767 17370 13776
rect 17224 13738 17276 13744
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11626 17172 12174
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17144 11150 17172 11562
rect 17236 11286 17264 13126
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17328 11218 17356 13670
rect 17420 12238 17448 14350
rect 17604 13530 17632 17274
rect 17696 15502 17724 18022
rect 17958 17983 18014 17992
rect 18064 17954 18092 20742
rect 18156 18290 18184 21898
rect 18248 21554 18276 21966
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18248 19961 18276 20402
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18234 19952 18290 19961
rect 18234 19887 18290 19896
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18248 18290 18276 18566
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18064 17926 18184 17954
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16590 17816 17138
rect 17866 16688 17922 16697
rect 17866 16623 17868 16632
rect 17920 16623 17922 16632
rect 17868 16594 17920 16600
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 16114 17816 16526
rect 17972 16250 18000 17206
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17512 13025 17540 13262
rect 17498 13016 17554 13025
rect 17604 12986 17632 13262
rect 17498 12951 17554 12960
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17696 12714 17724 14894
rect 17788 14618 17816 15846
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17788 12918 17816 13738
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17880 12782 17908 15302
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14006 18000 14758
rect 18064 14550 18092 17002
rect 18156 16425 18184 17926
rect 18142 16416 18198 16425
rect 18142 16351 18198 16360
rect 18156 16182 18184 16351
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17868 12776 17920 12782
rect 17774 12744 17830 12753
rect 17684 12708 17736 12714
rect 17868 12718 17920 12724
rect 17774 12679 17830 12688
rect 17684 12650 17736 12656
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12434 17632 12582
rect 17604 12406 17724 12434
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 8362 17172 11086
rect 17420 11082 17448 12038
rect 17512 11762 17540 12310
rect 17696 12238 17724 12406
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 11558 17540 11698
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11218 17540 11494
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17328 10266 17356 11018
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 8974 17264 9454
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17144 7478 17172 7754
rect 17420 7750 17448 11018
rect 17512 11014 17540 11154
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17604 9654 17632 12106
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17604 9058 17632 9590
rect 17696 9586 17724 12174
rect 17788 10742 17816 12679
rect 17972 12646 18000 13398
rect 18064 12753 18092 14214
rect 18156 13326 18184 15846
rect 18248 15570 18276 18226
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18708 17882 18736 21558
rect 18800 18834 18828 22714
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18892 17746 18920 18702
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18616 15892 18644 16186
rect 18708 16114 18736 17206
rect 18786 16824 18842 16833
rect 18786 16759 18788 16768
rect 18840 16759 18842 16768
rect 18880 16788 18932 16794
rect 18788 16730 18840 16736
rect 18880 16730 18932 16736
rect 18892 16522 18920 16730
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18786 16008 18842 16017
rect 18786 15943 18842 15952
rect 18616 15864 18736 15892
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18236 15360 18288 15366
rect 18328 15360 18380 15366
rect 18236 15302 18288 15308
rect 18326 15328 18328 15337
rect 18380 15328 18382 15337
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18050 12744 18106 12753
rect 18050 12679 18106 12688
rect 17960 12640 18012 12646
rect 17958 12608 17960 12617
rect 18052 12640 18104 12646
rect 18012 12608 18014 12617
rect 18052 12582 18104 12588
rect 17958 12543 18014 12552
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17880 11801 17908 12310
rect 17866 11792 17922 11801
rect 17866 11727 17922 11736
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17788 9722 17816 9930
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17512 9030 17632 9058
rect 17512 8838 17540 9030
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17512 7546 17540 8366
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17132 7472 17184 7478
rect 17130 7440 17132 7449
rect 17184 7440 17186 7449
rect 17130 7375 17186 7384
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17328 7177 17356 7346
rect 17408 7200 17460 7206
rect 17314 7168 17370 7177
rect 17408 7142 17460 7148
rect 17314 7103 17370 7112
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16578 5672 16634 5681
rect 16578 5607 16580 5616
rect 16632 5607 16634 5616
rect 16580 5578 16632 5584
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5234 16712 5510
rect 16776 5234 16804 6734
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16776 4826 16804 5170
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16304 2032 16356 2038
rect 16304 1974 16356 1980
rect 16118 1456 16174 1465
rect 16118 1391 16174 1400
rect 16132 1358 16160 1391
rect 16408 1358 16436 2790
rect 16684 1562 16712 4694
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16776 4146 16804 4422
rect 16948 4276 17000 4282
rect 17000 4236 17080 4264
rect 16948 4218 17000 4224
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16868 3534 16896 4014
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 3058 16896 3470
rect 17052 3097 17080 4236
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17144 3738 17172 4150
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17038 3088 17094 3097
rect 16856 3052 16908 3058
rect 17038 3023 17094 3032
rect 16856 2994 16908 3000
rect 17052 2514 17080 3023
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17236 2122 17264 6802
rect 17420 6338 17448 7142
rect 17604 6458 17632 8842
rect 17696 7410 17724 9522
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17880 7342 17908 11494
rect 17972 9450 18000 11698
rect 18064 10112 18092 12582
rect 18142 12336 18198 12345
rect 18142 12271 18198 12280
rect 18156 12238 18184 12271
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18248 11506 18276 15302
rect 18326 15263 18382 15272
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 14074 18368 14214
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18512 14068 18564 14074
rect 18708 14056 18736 15864
rect 18512 14010 18564 14016
rect 18616 14028 18736 14056
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18340 13841 18368 13874
rect 18326 13832 18382 13841
rect 18524 13802 18552 14010
rect 18326 13767 18382 13776
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18616 13716 18644 14028
rect 18694 13968 18750 13977
rect 18694 13903 18696 13912
rect 18748 13903 18750 13912
rect 18696 13874 18748 13880
rect 18616 13688 18736 13716
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18524 13190 18552 13466
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18708 12986 18736 13688
rect 18800 13161 18828 15943
rect 18984 15570 19012 17614
rect 19076 16182 19104 19722
rect 19168 16998 19196 24074
rect 19260 21350 19288 25910
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19720 22094 19748 25638
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19720 22066 19932 22094
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19260 19242 19288 21286
rect 19352 20942 19380 21422
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20534 19380 20878
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19352 18290 19380 19450
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 19168 16114 19196 16662
rect 19260 16164 19288 18226
rect 19352 17270 19380 18226
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16833 19380 16934
rect 19338 16824 19394 16833
rect 19338 16759 19394 16768
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19432 16448 19484 16454
rect 19430 16416 19432 16425
rect 19484 16416 19486 16425
rect 19430 16351 19486 16360
rect 19430 16280 19486 16289
rect 19536 16250 19564 16526
rect 19430 16215 19486 16224
rect 19524 16244 19576 16250
rect 19340 16176 19392 16182
rect 19260 16136 19340 16164
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19168 15881 19196 16050
rect 19154 15872 19210 15881
rect 19154 15807 19210 15816
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18984 15008 19012 15506
rect 18892 14980 19012 15008
rect 18892 14550 18920 14980
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18786 13152 18842 13161
rect 18786 13087 18842 13096
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18340 12646 18368 12854
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18708 12186 18736 12922
rect 18616 12170 18828 12186
rect 18604 12164 18828 12170
rect 18656 12158 18828 12164
rect 18604 12106 18656 12112
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18156 11478 18276 11506
rect 18156 11082 18184 11478
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18142 10976 18198 10985
rect 18142 10911 18198 10920
rect 18156 10266 18184 10911
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18064 10084 18184 10112
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 18064 9654 18092 9930
rect 18156 9654 18184 10084
rect 18248 10062 18276 11290
rect 18708 11234 18736 12038
rect 18524 11206 18736 11234
rect 18524 10470 18552 11206
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18512 10464 18564 10470
rect 18708 10441 18736 11018
rect 18512 10406 18564 10412
rect 18694 10432 18750 10441
rect 18315 10364 18623 10373
rect 18694 10367 18750 10376
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17958 9208 18014 9217
rect 17958 9143 18014 9152
rect 17972 8634 18000 9143
rect 18064 8809 18092 9590
rect 18708 9568 18736 10367
rect 18800 10266 18828 12158
rect 18892 11082 18920 13874
rect 18984 11830 19012 14826
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 11830 19104 13262
rect 19168 12918 19196 15807
rect 19260 15745 19288 16136
rect 19340 16118 19392 16124
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19246 15736 19302 15745
rect 19246 15671 19302 15680
rect 19260 15094 19288 15671
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19260 13190 19288 15030
rect 19352 14074 19380 15914
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12986 19288 13126
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19444 12918 19472 16215
rect 19524 16186 19576 16192
rect 19628 16114 19656 17818
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19720 16522 19748 16730
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19706 16144 19762 16153
rect 19616 16108 19668 16114
rect 19706 16079 19762 16088
rect 19616 16050 19668 16056
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19536 14006 19564 14894
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19536 12730 19564 13670
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19352 12702 19564 12730
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18616 9540 18736 9568
rect 18512 9512 18564 9518
rect 18142 9480 18198 9489
rect 18616 9500 18644 9540
rect 18564 9472 18644 9500
rect 18512 9454 18564 9460
rect 18142 9415 18198 9424
rect 18696 9444 18748 9450
rect 18050 8800 18106 8809
rect 18050 8735 18106 8744
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17958 8528 18014 8537
rect 18156 8498 18184 9415
rect 18696 9386 18748 9392
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18326 9072 18382 9081
rect 18326 9007 18382 9016
rect 18340 8974 18368 9007
rect 18524 8974 18552 9114
rect 18708 9058 18736 9386
rect 18616 9030 18736 9058
rect 18616 8974 18644 9030
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18432 8820 18460 8910
rect 18248 8792 18460 8820
rect 17958 8463 18014 8472
rect 18052 8492 18104 8498
rect 17972 8362 18000 8463
rect 18052 8434 18104 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18064 8401 18092 8434
rect 18050 8392 18106 8401
rect 17960 8356 18012 8362
rect 18050 8327 18106 8336
rect 17960 8298 18012 8304
rect 18248 7818 18276 8792
rect 18800 8616 18828 10202
rect 18892 8974 18920 10610
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18708 8588 18828 8616
rect 18326 8528 18382 8537
rect 18326 8463 18328 8472
rect 18380 8463 18382 8472
rect 18328 8434 18380 8440
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17972 7274 18000 7686
rect 18524 7410 18552 7822
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18708 6769 18736 8588
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18694 6760 18750 6769
rect 18694 6695 18696 6704
rect 18748 6695 18750 6704
rect 18696 6666 18748 6672
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17328 6310 17448 6338
rect 17604 6322 17632 6394
rect 17592 6316 17644 6322
rect 17328 6225 17356 6310
rect 17592 6258 17644 6264
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 17314 6216 17370 6225
rect 17314 6151 17370 6160
rect 17774 6216 17830 6225
rect 17774 6151 17830 6160
rect 17328 2689 17356 6151
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 4554 17448 5646
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17314 2680 17370 2689
rect 17314 2615 17370 2624
rect 17314 2544 17370 2553
rect 17314 2479 17370 2488
rect 17328 2446 17356 2479
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17316 2304 17368 2310
rect 17314 2272 17316 2281
rect 17368 2272 17370 2281
rect 17314 2207 17370 2216
rect 17052 2094 17264 2122
rect 17052 1970 17080 2094
rect 17512 2038 17540 6054
rect 17788 5710 17816 6151
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17604 5273 17632 5578
rect 17590 5264 17646 5273
rect 17590 5199 17646 5208
rect 17696 3126 17724 5578
rect 18156 5166 18184 6258
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18418 5808 18474 5817
rect 18418 5743 18474 5752
rect 18432 5302 18460 5743
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17788 2774 17816 4422
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17696 2746 17816 2774
rect 17696 2446 17724 2746
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17788 2310 17816 2615
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17696 2038 17724 2246
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17684 2032 17736 2038
rect 17684 1974 17736 1980
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 17788 1562 17816 2246
rect 16672 1556 16724 1562
rect 16672 1498 16724 1504
rect 17776 1556 17828 1562
rect 17776 1498 17828 1504
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 15936 1284 15988 1290
rect 15936 1226 15988 1232
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10508 1216 10560 1222
rect 10508 1158 10560 1164
rect 14740 1216 14792 1222
rect 14740 1158 14792 1164
rect 2226 912 2282 921
rect 2226 847 2282 856
rect 5368 785 5396 1158
rect 7896 1116 8204 1125
rect 7896 1114 7902 1116
rect 7958 1114 7982 1116
rect 8038 1114 8062 1116
rect 8118 1114 8142 1116
rect 8198 1114 8204 1116
rect 7958 1062 7960 1114
rect 8140 1062 8142 1114
rect 7896 1060 7902 1062
rect 7958 1060 7982 1062
rect 8038 1060 8062 1062
rect 8118 1060 8142 1062
rect 8198 1060 8204 1062
rect 7896 1051 8204 1060
rect 14842 1116 15150 1125
rect 14842 1114 14848 1116
rect 14904 1114 14928 1116
rect 14984 1114 15008 1116
rect 15064 1114 15088 1116
rect 15144 1114 15150 1116
rect 14904 1062 14906 1114
rect 15086 1062 15088 1114
rect 14842 1060 14848 1062
rect 14904 1060 14928 1062
rect 14984 1060 15008 1062
rect 15064 1060 15088 1062
rect 15144 1060 15150 1062
rect 14842 1051 15150 1060
rect 15948 1018 15976 1226
rect 17880 1222 17908 3062
rect 17972 2650 18000 5034
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4554 18092 4626
rect 18142 4584 18198 4593
rect 18052 4548 18104 4554
rect 18142 4519 18144 4528
rect 18052 4490 18104 4496
rect 18196 4519 18198 4528
rect 18144 4490 18196 4496
rect 18248 3194 18276 5238
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18156 2650 18184 2790
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18328 2576 18380 2582
rect 18326 2544 18328 2553
rect 18380 2544 18382 2553
rect 18052 2508 18104 2514
rect 18326 2479 18382 2488
rect 18708 2530 18736 5850
rect 18800 5778 18828 8434
rect 18878 8392 18934 8401
rect 18878 8327 18880 8336
rect 18932 8327 18934 8336
rect 18880 8298 18932 8304
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18892 5914 18920 7890
rect 18984 7478 19012 11222
rect 19076 8022 19104 11766
rect 19168 10742 19196 12650
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19168 9926 19196 10542
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18984 6882 19012 7278
rect 19076 7206 19104 7686
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18984 6854 19104 6882
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18984 5642 19012 6666
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18984 4690 19012 5578
rect 19076 5302 19104 6854
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18892 2650 18920 3062
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18708 2514 18828 2530
rect 18708 2508 18840 2514
rect 18708 2502 18788 2508
rect 18052 2450 18104 2456
rect 18064 1358 18092 2450
rect 18315 1660 18623 1669
rect 18315 1658 18321 1660
rect 18377 1658 18401 1660
rect 18457 1658 18481 1660
rect 18537 1658 18561 1660
rect 18617 1658 18623 1660
rect 18377 1606 18379 1658
rect 18559 1606 18561 1658
rect 18315 1604 18321 1606
rect 18377 1604 18401 1606
rect 18457 1604 18481 1606
rect 18537 1604 18561 1606
rect 18617 1604 18623 1606
rect 18315 1595 18623 1604
rect 18708 1442 18736 2502
rect 18788 2450 18840 2456
rect 18984 2281 19012 2586
rect 19168 2446 19196 9318
rect 19260 9178 19288 12242
rect 19352 10810 19380 12702
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12050 19472 12582
rect 19522 12336 19578 12345
rect 19522 12271 19578 12280
rect 19536 12170 19564 12271
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19444 12022 19564 12050
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19340 10192 19392 10198
rect 19338 10160 19340 10169
rect 19392 10160 19394 10169
rect 19338 10095 19394 10104
rect 19340 10056 19392 10062
rect 19444 10044 19472 11834
rect 19536 11218 19564 12022
rect 19628 11762 19656 15302
rect 19720 14550 19748 16079
rect 19812 15434 19840 21286
rect 19904 20466 19932 22066
rect 20088 21350 20116 22578
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19904 17066 19932 20402
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19996 19922 20024 20334
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20180 18986 20208 21830
rect 20272 19174 20300 26726
rect 20640 22438 20668 26930
rect 20732 24274 20760 26998
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 21836 26450 21864 26862
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20732 23118 20760 24210
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22710 20760 23054
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20180 18958 20300 18986
rect 20272 18766 20300 18958
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19904 15314 19932 16662
rect 19996 16289 20024 18566
rect 20088 18426 20116 18702
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 17202 20208 17546
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 19982 16280 20038 16289
rect 19982 16215 20038 16224
rect 20180 16182 20208 17138
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 20168 16176 20220 16182
rect 20220 16136 20300 16164
rect 20168 16118 20220 16124
rect 19812 15286 19932 15314
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19720 14414 19748 14486
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19706 13288 19762 13297
rect 19706 13223 19762 13232
rect 19720 11830 19748 13223
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19628 10606 19656 11698
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19536 10062 19564 10474
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10305 19656 10406
rect 19614 10296 19670 10305
rect 19614 10231 19670 10240
rect 19616 10192 19668 10198
rect 19614 10160 19616 10169
rect 19668 10160 19670 10169
rect 19614 10095 19670 10104
rect 19392 10016 19472 10044
rect 19524 10056 19576 10062
rect 19340 9998 19392 10004
rect 19524 9998 19576 10004
rect 19522 9888 19578 9897
rect 19522 9823 19578 9832
rect 19338 9752 19394 9761
rect 19536 9722 19564 9823
rect 19338 9687 19394 9696
rect 19524 9716 19576 9722
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19352 9042 19380 9687
rect 19524 9658 19576 9664
rect 19522 9616 19578 9625
rect 19522 9551 19578 9560
rect 19536 9450 19564 9551
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19614 9344 19670 9353
rect 19614 9279 19670 9288
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8294 19288 8910
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19338 8664 19394 8673
rect 19338 8599 19340 8608
rect 19392 8599 19394 8608
rect 19340 8570 19392 8576
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19260 7342 19288 8230
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19260 5778 19288 6258
rect 19352 6118 19380 8434
rect 19444 8265 19472 8842
rect 19430 8256 19486 8265
rect 19430 8191 19486 8200
rect 19430 8120 19486 8129
rect 19430 8055 19486 8064
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19260 3602 19288 5714
rect 19444 4622 19472 8055
rect 19536 4758 19564 9114
rect 19628 8498 19656 9279
rect 19720 8974 19748 11494
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19706 8800 19762 8809
rect 19706 8735 19762 8744
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 19628 6798 19656 8327
rect 19720 7970 19748 8735
rect 19812 8498 19840 15286
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19904 13870 19932 15030
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19904 12753 19932 12786
rect 19890 12744 19946 12753
rect 19890 12679 19946 12688
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 11257 19932 12582
rect 19996 12345 20024 16118
rect 20168 15904 20220 15910
rect 20272 15881 20300 16136
rect 20364 15910 20392 21490
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18970 20484 19110
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17202 20484 18022
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16794 20484 17138
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20442 16688 20498 16697
rect 20442 16623 20498 16632
rect 20456 16590 20484 16623
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20352 15904 20404 15910
rect 20168 15846 20220 15852
rect 20258 15872 20314 15881
rect 20076 15088 20128 15094
rect 20074 15056 20076 15065
rect 20128 15056 20130 15065
rect 20074 14991 20130 15000
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20088 13462 20116 13670
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19982 12336 20038 12345
rect 19982 12271 20038 12280
rect 19996 11268 20024 12271
rect 20180 12170 20208 15846
rect 20352 15846 20404 15852
rect 20258 15807 20314 15816
rect 20272 15502 20300 15807
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20456 14226 20484 16526
rect 20548 14346 20576 21558
rect 20640 18358 20668 22374
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 19854 20760 20878
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20732 18766 20760 19790
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20628 17672 20680 17678
rect 20732 17660 20760 18566
rect 20680 17632 20760 17660
rect 20628 17614 20680 17620
rect 20628 17060 20680 17066
rect 20732 17048 20760 17632
rect 20680 17020 20760 17048
rect 20628 17002 20680 17008
rect 20732 16674 20760 17020
rect 20824 16794 20852 18838
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20916 17134 20944 17478
rect 21008 17202 21036 17478
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20732 16646 20852 16674
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20640 15706 20668 15846
rect 20732 15706 20760 16458
rect 20824 15994 20852 16646
rect 20916 16182 20944 17070
rect 21008 16182 21036 17138
rect 21100 16590 21128 18226
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20824 15966 20944 15994
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20732 15570 20760 15642
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20718 15464 20774 15473
rect 20718 15399 20720 15408
rect 20772 15399 20774 15408
rect 20720 15370 20772 15376
rect 20916 15366 20944 15966
rect 21008 15910 21036 16118
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21100 15586 21128 15982
rect 21192 15910 21220 23598
rect 21468 21622 21496 26386
rect 22572 26314 22600 27270
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22848 26586 22876 26930
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21560 21894 21588 24006
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21652 22642 21680 22918
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21652 22030 21680 22578
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 21284 16561 21312 18634
rect 21364 18352 21416 18358
rect 21364 18294 21416 18300
rect 21270 16552 21326 16561
rect 21270 16487 21326 16496
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 16017 21312 16390
rect 21376 16114 21404 18294
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21270 16008 21326 16017
rect 21270 15943 21326 15952
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21008 15558 21128 15586
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20456 14198 20576 14226
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20258 13968 20314 13977
rect 20258 13903 20260 13912
rect 20312 13903 20314 13912
rect 20260 13874 20312 13880
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20272 13297 20300 13330
rect 20364 13326 20392 14010
rect 20352 13320 20404 13326
rect 20258 13288 20314 13297
rect 20352 13262 20404 13268
rect 20258 13223 20314 13232
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20272 12345 20300 12378
rect 20258 12336 20314 12345
rect 20258 12271 20314 12280
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20548 11830 20576 14198
rect 20640 13938 20668 15030
rect 20916 14822 20944 15302
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20640 12918 20668 13874
rect 20916 13734 20944 14758
rect 21008 14278 21036 15558
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 14346 21128 15438
rect 21180 14816 21232 14822
rect 21178 14784 21180 14793
rect 21232 14784 21234 14793
rect 21178 14719 21234 14728
rect 21284 14618 21312 15846
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20824 13138 20852 13194
rect 20732 13110 20852 13138
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20076 11280 20128 11286
rect 19890 11248 19946 11257
rect 19996 11240 20076 11268
rect 20076 11222 20128 11228
rect 19890 11183 19946 11192
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10713 19932 11086
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19996 10742 20024 11018
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19984 10736 20036 10742
rect 19890 10704 19946 10713
rect 19984 10678 20036 10684
rect 19890 10639 19946 10648
rect 19890 10432 19946 10441
rect 19890 10367 19946 10376
rect 19904 10062 19932 10367
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 9761 19932 9862
rect 19890 9752 19946 9761
rect 19890 9687 19946 9696
rect 19892 9648 19944 9654
rect 19890 9616 19892 9625
rect 19944 9616 19946 9625
rect 19890 9551 19946 9560
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19904 9110 19932 9454
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19904 8634 19932 8774
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19720 7942 19840 7970
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19628 5574 19656 6734
rect 19720 5778 19748 7822
rect 19812 7188 19840 7942
rect 19904 7886 19932 8230
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19904 7290 19932 7414
rect 19996 7410 20024 10678
rect 20088 8974 20116 10950
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 20088 7936 20116 8774
rect 20180 8362 20208 11630
rect 20272 9722 20300 11698
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 10062 20392 11630
rect 20626 11384 20682 11393
rect 20626 11319 20628 11328
rect 20680 11319 20682 11328
rect 20628 11290 20680 11296
rect 20444 11280 20496 11286
rect 20732 11234 20760 13110
rect 21008 12238 21036 13738
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21100 12306 21128 12922
rect 21192 12442 21220 14350
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21100 11898 21128 12242
rect 21180 12232 21232 12238
rect 21178 12200 21180 12209
rect 21232 12200 21234 12209
rect 21178 12135 21234 12144
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21284 11778 21312 14418
rect 21376 13818 21404 15098
rect 21468 14618 21496 18702
rect 21560 15502 21588 21830
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20534 21680 20742
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 22296 20466 22324 21830
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22204 19417 22232 19654
rect 22190 19408 22246 19417
rect 22190 19343 22246 19352
rect 22192 18624 22244 18630
rect 22190 18592 22192 18601
rect 22244 18592 22246 18601
rect 21788 18524 22096 18533
rect 22190 18527 22246 18536
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22112 17610 22140 18294
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22296 17338 22324 20402
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21652 16114 21680 17070
rect 22388 16674 22416 20810
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22480 17610 22508 19382
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22296 16646 22416 16674
rect 22112 16522 22232 16538
rect 22100 16516 22232 16522
rect 22152 16510 22232 16516
rect 22100 16458 22152 16464
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21914 15600 21970 15609
rect 21914 15535 21916 15544
rect 21968 15535 21970 15544
rect 21916 15506 21968 15512
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21730 15464 21786 15473
rect 21652 15408 21730 15416
rect 21652 15388 21732 15408
rect 21652 15008 21680 15388
rect 21784 15399 21786 15408
rect 21732 15370 21784 15376
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 21560 14980 21680 15008
rect 22008 15020 22060 15026
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21456 13864 21508 13870
rect 21376 13812 21456 13818
rect 21376 13806 21508 13812
rect 21376 13790 21496 13806
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 20444 11222 20496 11228
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20272 8838 20300 9658
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20364 8566 20392 9998
rect 20456 9518 20484 11222
rect 20640 11206 20760 11234
rect 21100 11750 21312 11778
rect 20640 10674 20668 11206
rect 21100 11150 21128 11750
rect 21376 11218 21404 13670
rect 21468 11762 21496 13790
rect 21560 12442 21588 14980
rect 22008 14962 22060 14968
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21456 11552 21508 11558
rect 21454 11520 21456 11529
rect 21508 11520 21510 11529
rect 21510 11478 21588 11506
rect 21454 11455 21510 11464
rect 21454 11384 21510 11393
rect 21454 11319 21510 11328
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20640 10577 20668 10610
rect 20626 10568 20682 10577
rect 20626 10503 20682 10512
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20548 9994 20576 10202
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20732 9874 20760 11086
rect 21468 11082 21496 11319
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 20994 10976 21050 10985
rect 20994 10911 21050 10920
rect 21008 10266 21036 10911
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21180 10464 21232 10470
rect 21086 10432 21142 10441
rect 21180 10406 21232 10412
rect 21086 10367 21142 10376
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21100 10062 21128 10367
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20640 9846 20760 9874
rect 20640 9625 20668 9846
rect 20824 9738 20852 9930
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20994 9888 21050 9897
rect 20732 9710 20852 9738
rect 20626 9616 20682 9625
rect 20626 9551 20682 9560
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 9042 20484 9454
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20364 8294 20392 8502
rect 20456 8498 20484 8978
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20272 8266 20392 8294
rect 20088 7908 20208 7936
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 20088 7290 20116 7754
rect 19904 7262 20116 7290
rect 19812 7160 19932 7188
rect 19904 6662 19932 7160
rect 20074 6896 20130 6905
rect 20180 6866 20208 7908
rect 20272 7410 20300 8266
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20074 6831 20130 6840
rect 20168 6860 20220 6866
rect 20088 6730 20116 6831
rect 20168 6802 20220 6808
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19812 6225 19840 6598
rect 19798 6216 19854 6225
rect 19798 6151 19854 6160
rect 19904 6100 19932 6598
rect 20272 6186 20300 6734
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 19812 6072 19932 6100
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19708 4548 19760 4554
rect 19812 4536 19840 6072
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 20180 4826 20208 5102
rect 20364 5030 20392 7686
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20548 7426 20576 9318
rect 20732 9110 20760 9710
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20626 8936 20682 8945
rect 20626 8871 20628 8880
rect 20680 8871 20682 8880
rect 20628 8842 20680 8848
rect 20626 8664 20682 8673
rect 20626 8599 20682 8608
rect 20640 8498 20668 8599
rect 20824 8566 20852 9386
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20824 8090 20852 8502
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20916 8022 20944 9862
rect 20994 9823 21050 9832
rect 21008 9586 21036 9823
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 8838 21036 9522
rect 21100 8906 21128 9998
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7546 20668 7754
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20456 6322 20484 7414
rect 20548 7398 20668 7426
rect 20640 6798 20668 7398
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20628 6792 20680 6798
rect 20534 6760 20590 6769
rect 20628 6734 20680 6740
rect 20534 6695 20536 6704
rect 20588 6695 20590 6704
rect 20536 6666 20588 6672
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5574 20576 6258
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 19760 4508 19840 4536
rect 19708 4490 19760 4496
rect 19904 4282 19932 4558
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 20548 4214 20576 4558
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19352 3534 19380 4150
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 2990 19380 3470
rect 19536 3126 19564 3878
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 18970 2272 19026 2281
rect 18970 2207 19026 2216
rect 18432 1414 18736 1442
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 18432 1290 18460 1414
rect 18420 1284 18472 1290
rect 18420 1226 18472 1232
rect 19260 1222 19288 2314
rect 19536 1358 19564 3062
rect 19720 2038 19748 4082
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3738 20576 3878
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20640 3618 20668 6734
rect 20732 4554 20760 7278
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 6390 20944 6598
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20548 3590 20668 3618
rect 19708 2032 19760 2038
rect 19708 1974 19760 1980
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 17868 1216 17920 1222
rect 17868 1158 17920 1164
rect 19248 1216 19300 1222
rect 19248 1158 19300 1164
rect 15936 1012 15988 1018
rect 15936 954 15988 960
rect 19720 950 19748 1974
rect 20548 1358 20576 3590
rect 20732 3194 20760 4490
rect 20824 3534 20852 5306
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20536 1352 20588 1358
rect 20536 1294 20588 1300
rect 20168 1284 20220 1290
rect 20168 1226 20220 1232
rect 19708 944 19760 950
rect 19708 886 19760 892
rect 20180 882 20208 1226
rect 20640 1222 20668 2518
rect 20732 1970 20760 2994
rect 20824 2774 20852 3470
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 3058 20944 3402
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20824 2746 20944 2774
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20916 1358 20944 2746
rect 21008 2394 21036 8570
rect 21192 8514 21220 10406
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21100 8486 21220 8514
rect 21100 7313 21128 8486
rect 21086 7304 21142 7313
rect 21086 7239 21142 7248
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21192 5642 21220 6734
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21008 2366 21128 2394
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21008 1970 21036 2246
rect 21100 1970 21128 2366
rect 21284 2106 21312 10202
rect 21376 10169 21404 10746
rect 21560 10674 21588 11478
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21362 10160 21418 10169
rect 21362 10095 21418 10104
rect 21362 9752 21418 9761
rect 21362 9687 21364 9696
rect 21416 9687 21418 9696
rect 21364 9658 21416 9664
rect 21468 5914 21496 10474
rect 21560 7954 21588 10610
rect 21652 10130 21680 14826
rect 22020 14260 22048 14962
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22112 14414 22140 14894
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22204 14362 22232 16510
rect 22296 15366 22324 16646
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22480 16538 22508 17546
rect 22572 16726 22600 26250
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22756 21146 22784 21286
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22664 19718 22692 19790
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22388 16402 22416 16526
rect 22480 16510 22600 16538
rect 22388 16374 22508 16402
rect 22480 16250 22508 16374
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22388 15706 22416 16186
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22572 15586 22600 16510
rect 22664 16153 22692 19654
rect 22650 16144 22706 16153
rect 22650 16079 22706 16088
rect 22756 15994 22784 21082
rect 22848 17882 22876 26522
rect 23204 26240 23256 26246
rect 23204 26182 23256 26188
rect 23216 24138 23244 26182
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 22710 24164 24006
rect 24412 23798 24440 26726
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24400 23792 24452 23798
rect 24400 23734 24452 23740
rect 24596 23662 24624 24142
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24596 23186 24624 23598
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22480 15558 22600 15586
rect 22664 15966 22784 15994
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22388 14770 22416 15438
rect 22296 14742 22416 14770
rect 22296 14482 22324 14742
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22204 14334 22324 14362
rect 22020 14232 22232 14260
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22204 14056 22232 14232
rect 22020 14028 22232 14056
rect 22020 13326 22048 14028
rect 22190 13696 22246 13705
rect 22190 13631 22246 13640
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 22204 11762 22232 13631
rect 22296 12646 22324 14334
rect 22388 14074 22416 14554
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22480 14006 22508 15558
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22572 15162 22600 15438
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22572 13818 22600 14894
rect 22664 14822 22692 15966
rect 22742 15736 22798 15745
rect 22742 15671 22798 15680
rect 22756 15434 22784 15671
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22848 15337 22876 16390
rect 22940 15570 22968 18702
rect 23124 18601 23152 21558
rect 23308 21554 23336 21830
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23204 21480 23256 21486
rect 23400 21434 23428 22578
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23204 21422 23256 21428
rect 23216 20942 23244 21422
rect 23308 21406 23428 21434
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23216 20534 23244 20878
rect 23204 20528 23256 20534
rect 23204 20470 23256 20476
rect 23216 20058 23244 20470
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23216 19378 23244 19994
rect 23308 19514 23336 21406
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 19786 23428 20198
rect 23492 20058 23520 21490
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23664 20324 23716 20330
rect 23664 20266 23716 20272
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23110 18592 23166 18601
rect 23110 18527 23166 18536
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23032 17678 23060 18158
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23308 17270 23336 19450
rect 23388 19440 23440 19446
rect 23386 19408 23388 19417
rect 23440 19408 23442 19417
rect 23386 19343 23442 19352
rect 23492 18766 23520 19994
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23032 16046 23060 16934
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22834 15328 22890 15337
rect 22834 15263 22890 15272
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22480 13790 22600 13818
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12850 22416 13126
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22480 12730 22508 13790
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22388 12702 22508 12730
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22112 11506 22140 11630
rect 22112 11478 22232 11506
rect 22204 11286 22232 11478
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22190 10840 22246 10849
rect 22190 10775 22246 10784
rect 22204 10742 22232 10775
rect 22008 10736 22060 10742
rect 22192 10736 22244 10742
rect 22060 10696 22140 10724
rect 22008 10678 22060 10684
rect 22008 10600 22060 10606
rect 22112 10577 22140 10696
rect 22192 10678 22244 10684
rect 22008 10542 22060 10548
rect 22098 10568 22154 10577
rect 21730 10296 21786 10305
rect 22020 10266 22048 10542
rect 22098 10503 22154 10512
rect 21730 10231 21786 10240
rect 22008 10260 22060 10266
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21744 10010 21772 10231
rect 22008 10202 22060 10208
rect 22296 10062 22324 12038
rect 22388 11082 22416 12702
rect 22572 12594 22600 12786
rect 22664 12594 22692 14282
rect 22756 13462 22784 14758
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22848 13308 22876 14010
rect 22756 13280 22876 13308
rect 22756 13190 22784 13280
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22480 12566 22600 12594
rect 22655 12566 22692 12594
rect 22480 12374 22508 12566
rect 22655 12458 22683 12566
rect 22572 12430 22683 12458
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22480 12238 22508 12310
rect 22572 12238 22600 12430
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22652 12232 22704 12238
rect 22756 12220 22784 12786
rect 22848 12753 22876 13126
rect 22834 12744 22890 12753
rect 22834 12679 22890 12688
rect 23032 12322 23060 15846
rect 22704 12192 22784 12220
rect 22848 12294 23060 12322
rect 22652 12174 22704 12180
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22376 10736 22428 10742
rect 22374 10704 22376 10713
rect 22428 10704 22430 10713
rect 22374 10639 22430 10648
rect 22376 10600 22428 10606
rect 22480 10577 22508 12174
rect 22664 12084 22692 12174
rect 22572 12056 22692 12084
rect 22742 12064 22798 12073
rect 22572 11830 22600 12056
rect 22742 11999 22798 12008
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22664 11642 22692 11834
rect 22756 11830 22784 11999
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22664 11614 22784 11642
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22376 10542 22428 10548
rect 22466 10568 22522 10577
rect 21652 9982 21772 10010
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21652 7528 21680 9982
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22020 8498 22048 8570
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22112 7886 22140 7958
rect 21824 7880 21876 7886
rect 21822 7848 21824 7857
rect 22100 7880 22152 7886
rect 21876 7848 21878 7857
rect 22100 7822 22152 7828
rect 21822 7783 21878 7792
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 21560 7500 21680 7528
rect 21560 6254 21588 7500
rect 22204 7478 22232 8774
rect 22282 8256 22338 8265
rect 22282 8191 22338 8200
rect 22296 8090 22324 8191
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22282 7984 22338 7993
rect 22282 7919 22338 7928
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 4282 21404 5646
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21272 2100 21324 2106
rect 21272 2042 21324 2048
rect 20996 1964 21048 1970
rect 20996 1906 21048 1912
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 21100 1465 21128 1906
rect 21468 1902 21496 5578
rect 21560 4826 21588 6190
rect 21652 5710 21680 7346
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21744 6866 21772 6938
rect 21916 6928 21968 6934
rect 21822 6896 21878 6905
rect 21732 6860 21784 6866
rect 21916 6870 21968 6876
rect 21822 6831 21878 6840
rect 21732 6802 21784 6808
rect 21836 6798 21864 6831
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21928 6730 21956 6870
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 22296 6225 22324 7919
rect 22388 7546 22416 10542
rect 22466 10503 22522 10512
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22480 9897 22508 9930
rect 22466 9888 22522 9897
rect 22466 9823 22522 9832
rect 22572 9761 22600 11222
rect 22664 11150 22692 11494
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 10033 22692 10406
rect 22650 10024 22706 10033
rect 22650 9959 22706 9968
rect 22558 9752 22614 9761
rect 22756 9738 22784 11614
rect 22848 11150 22876 12294
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 23032 12050 23060 12106
rect 22940 12022 23060 12050
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22834 10704 22890 10713
rect 22834 10639 22836 10648
rect 22888 10639 22890 10648
rect 22836 10610 22888 10616
rect 22558 9687 22614 9696
rect 22664 9710 22784 9738
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22282 6216 22338 6225
rect 22282 6151 22338 6160
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21652 2038 21680 5646
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22296 4434 22324 6054
rect 22388 5710 22416 6870
rect 22480 5778 22508 9522
rect 22572 9382 22600 9687
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22572 8616 22600 9318
rect 22664 8786 22692 9710
rect 22742 9616 22798 9625
rect 22742 9551 22744 9560
rect 22796 9551 22798 9560
rect 22744 9522 22796 9528
rect 22836 8832 22888 8838
rect 22664 8758 22784 8786
rect 22836 8774 22888 8780
rect 22940 8786 22968 12022
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23032 11762 23060 11834
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23124 11506 23152 16934
rect 23202 16688 23258 16697
rect 23202 16623 23204 16632
rect 23256 16623 23258 16632
rect 23204 16594 23256 16600
rect 23308 16590 23336 17002
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23216 14958 23244 15370
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23032 11478 23152 11506
rect 23032 11354 23060 11478
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23032 11218 23060 11290
rect 23110 11248 23166 11257
rect 23020 11212 23072 11218
rect 23110 11183 23166 11192
rect 23020 11154 23072 11160
rect 23124 11098 23152 11183
rect 23032 11070 23152 11098
rect 23032 9450 23060 11070
rect 23216 10441 23244 14350
rect 23308 14346 23336 16390
rect 23400 15434 23428 16526
rect 23492 16289 23520 18294
rect 23478 16280 23534 16289
rect 23478 16215 23534 16224
rect 23478 16144 23534 16153
rect 23478 16079 23480 16088
rect 23532 16079 23534 16088
rect 23480 16050 23532 16056
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23492 15026 23520 15370
rect 23584 15026 23612 18838
rect 23676 17202 23704 20266
rect 23860 18358 23888 20742
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23952 18086 23980 22646
rect 24596 22642 24624 23122
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24596 22098 24624 22578
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24492 21956 24544 21962
rect 24492 21898 24544 21904
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 23940 17604 23992 17610
rect 23940 17546 23992 17552
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23676 14906 23704 17138
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 23768 16538 23796 16662
rect 23768 16510 23888 16538
rect 23754 16280 23810 16289
rect 23754 16215 23810 16224
rect 23768 15026 23796 16215
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23584 14878 23704 14906
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 23308 13274 23336 13942
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 13410 23428 13670
rect 23584 13530 23612 14878
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 13938 23704 14214
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23676 13530 23704 13670
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23400 13382 23704 13410
rect 23676 13326 23704 13382
rect 23572 13320 23624 13326
rect 23308 13246 23428 13274
rect 23572 13262 23624 13268
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23400 12730 23428 13246
rect 23308 12702 23428 12730
rect 23308 12170 23336 12702
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23492 12442 23520 12582
rect 23584 12442 23612 13262
rect 23768 12968 23796 13670
rect 23676 12940 23796 12968
rect 23676 12782 23704 12940
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23400 12322 23428 12378
rect 23400 12294 23520 12322
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23308 11121 23336 11154
rect 23294 11112 23350 11121
rect 23294 11047 23350 11056
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23202 10432 23258 10441
rect 23202 10367 23258 10376
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23216 10062 23244 10202
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 23124 9382 23152 9998
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 8906 23152 9318
rect 23112 8900 23164 8906
rect 23112 8842 23164 8848
rect 22572 8588 22692 8616
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22572 8294 22600 8434
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22572 7342 22600 8230
rect 22664 7818 22692 8588
rect 22756 7993 22784 8758
rect 22742 7984 22798 7993
rect 22742 7919 22798 7928
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22558 6216 22614 6225
rect 22558 6151 22614 6160
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 22204 3058 22232 4422
rect 22296 4406 22416 4434
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22296 3602 22324 4150
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22296 3126 22324 3538
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22296 2446 22324 3062
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 22296 2106 22324 2382
rect 22388 2378 22416 4406
rect 22480 3534 22508 5034
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22376 2372 22428 2378
rect 22376 2314 22428 2320
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 21640 2032 21692 2038
rect 21640 1974 21692 1980
rect 21456 1896 21508 1902
rect 21456 1838 21508 1844
rect 21086 1456 21142 1465
rect 21468 1426 21496 1838
rect 21086 1391 21142 1400
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 22296 1358 22324 2042
rect 22572 1562 22600 6151
rect 22756 5914 22784 7822
rect 22848 6798 22876 8774
rect 22940 8758 23152 8786
rect 22928 7880 22980 7886
rect 22980 7840 23060 7868
rect 22928 7822 22980 7828
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22848 5302 22876 6734
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 22836 5296 22888 5302
rect 22836 5238 22888 5244
rect 22940 4622 22968 6122
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 4214 22692 4422
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22664 2038 22692 3470
rect 22940 3194 22968 4558
rect 23032 3738 23060 7840
rect 23124 6390 23152 8758
rect 23216 8090 23244 9862
rect 23308 9178 23336 10950
rect 23400 10849 23428 11494
rect 23386 10840 23442 10849
rect 23386 10775 23442 10784
rect 23492 10674 23520 12294
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23584 11762 23612 11834
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23572 11620 23624 11626
rect 23572 11562 23624 11568
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23400 10266 23428 10610
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23584 10198 23612 11562
rect 23676 11286 23704 11630
rect 23664 11280 23716 11286
rect 23664 11222 23716 11228
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23400 8974 23428 9522
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23308 6934 23336 7958
rect 23400 7857 23428 8230
rect 23386 7848 23442 7857
rect 23386 7783 23442 7792
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 22652 2032 22704 2038
rect 22652 1974 22704 1980
rect 23032 1970 23060 3674
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23308 2106 23336 2994
rect 23296 2100 23348 2106
rect 23296 2042 23348 2048
rect 23020 1964 23072 1970
rect 23020 1906 23072 1912
rect 22560 1556 22612 1562
rect 22560 1498 22612 1504
rect 23400 1358 23428 7783
rect 23492 6662 23520 9998
rect 23676 9722 23704 10610
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23584 7342 23612 8570
rect 23768 7818 23796 11766
rect 23860 10810 23888 16510
rect 23952 15910 23980 17546
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 24044 13734 24072 17478
rect 24136 15473 24164 18158
rect 24412 18086 24440 20402
rect 24400 18080 24452 18086
rect 24398 18048 24400 18057
rect 24452 18048 24454 18057
rect 24398 17983 24454 17992
rect 24504 17066 24532 21898
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24780 18358 24808 18634
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24122 15464 24178 15473
rect 24122 15399 24178 15408
rect 24136 15026 24164 15399
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24136 13938 24164 14350
rect 24228 14056 24256 16730
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24320 15162 24348 16526
rect 24596 16114 24624 16526
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15910 24624 16050
rect 24780 16046 24808 18294
rect 24872 18290 24900 21286
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 24872 16522 24900 17750
rect 24964 17354 24992 19314
rect 25056 18834 25084 26250
rect 25148 25838 25176 26318
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26160 26042 26188 26250
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 26148 26036 26200 26042
rect 26148 25978 26200 25984
rect 25596 25968 25648 25974
rect 25596 25910 25648 25916
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 24206 25176 25774
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 21962 25176 22374
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25608 21350 25636 25910
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25976 25401 26004 25434
rect 25962 25392 26018 25401
rect 25962 25327 26018 25336
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25148 20262 25176 20810
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24964 17326 25084 17354
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24596 15570 24624 15846
rect 24584 15564 24636 15570
rect 24872 15552 24900 16458
rect 24584 15506 24636 15512
rect 24688 15524 24900 15552
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24320 14346 24348 15098
rect 24412 15026 24440 15370
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24412 14414 24440 14962
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24228 14028 24348 14056
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24136 13258 24164 13874
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24032 12844 24084 12850
rect 24084 12804 24164 12832
rect 24032 12786 24084 12792
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9654 23888 10406
rect 24044 10198 24072 11018
rect 24136 10810 24164 12804
rect 24228 11898 24256 13874
rect 24320 12850 24348 14028
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24124 10804 24176 10810
rect 24124 10746 24176 10752
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 24122 9752 24178 9761
rect 24122 9687 24178 9696
rect 24136 9654 24164 9687
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24044 9081 24072 9114
rect 24030 9072 24086 9081
rect 24030 9007 24086 9016
rect 23938 8936 23994 8945
rect 23938 8871 23994 8880
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23952 7002 23980 8871
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24136 7274 24164 8298
rect 24228 7546 24256 11834
rect 24320 11801 24348 12786
rect 24306 11792 24362 11801
rect 24306 11727 24362 11736
rect 24320 11393 24348 11727
rect 24306 11384 24362 11393
rect 24306 11319 24362 11328
rect 24412 11257 24440 14214
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24398 11248 24454 11257
rect 24398 11183 24454 11192
rect 24504 11014 24532 13262
rect 24688 12918 24716 15524
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 14074 24900 15370
rect 24964 15094 24992 17206
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 25056 13410 25084 17326
rect 25148 16590 25176 20198
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19310 25268 19654
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 24872 13382 25084 13410
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24780 12782 24808 13194
rect 24872 12850 24900 13382
rect 25056 13258 25084 13382
rect 25148 14396 25176 15982
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25608 15366 25636 16118
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25228 14408 25280 14414
rect 25148 14368 25228 14396
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24584 12708 24636 12714
rect 24584 12650 24636 12656
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24320 8022 24348 10950
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24412 8906 24440 10678
rect 24490 10160 24546 10169
rect 24490 10095 24546 10104
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24398 8800 24454 8809
rect 24398 8735 24454 8744
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23480 6656 23532 6662
rect 23676 6610 23704 6666
rect 23532 6604 23704 6610
rect 23480 6598 23704 6604
rect 23492 6582 23704 6598
rect 23676 4706 23704 6582
rect 24136 5574 24164 7210
rect 24306 6760 24362 6769
rect 24306 6695 24362 6704
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24044 4826 24072 5510
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 23676 4678 24164 4706
rect 24320 4690 24348 6695
rect 24412 5166 24440 8735
rect 24504 5302 24532 10095
rect 24596 6458 24624 12650
rect 24780 12238 24808 12718
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24964 11778 24992 13194
rect 25148 13138 25176 14368
rect 25228 14350 25280 14356
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25056 13110 25176 13138
rect 25056 12073 25084 13110
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25042 12064 25098 12073
rect 25042 11999 25098 12008
rect 25042 11928 25098 11937
rect 25042 11863 25044 11872
rect 25096 11863 25098 11872
rect 25044 11834 25096 11840
rect 24688 11750 24992 11778
rect 24688 11150 24716 11750
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 11529 24808 11630
rect 24766 11520 24822 11529
rect 24766 11455 24822 11464
rect 24780 11150 24808 11455
rect 24964 11286 24992 11750
rect 25148 11354 25176 12922
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25424 12170 25452 12378
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25516 11762 25544 12106
rect 25608 12102 25636 15302
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 25056 11234 25084 11290
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24780 10418 24808 10746
rect 24872 10674 24900 11222
rect 25056 11218 25268 11234
rect 25056 11212 25280 11218
rect 25056 11206 25228 11212
rect 25228 11154 25280 11160
rect 24952 11144 25004 11150
rect 25608 11098 25636 11766
rect 24952 11086 25004 11092
rect 24964 11014 24992 11086
rect 25516 11070 25636 11098
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25332 10674 25360 10746
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24780 10390 24900 10418
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24766 10160 24822 10169
rect 24688 6458 24716 10134
rect 24766 10095 24822 10104
rect 24780 10062 24808 10095
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24872 8634 24900 10390
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24964 8566 24992 10542
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24768 8424 24820 8430
rect 24820 8372 24900 8378
rect 24768 8366 24900 8372
rect 24780 8350 24900 8366
rect 24872 7886 24900 8350
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24872 6798 24900 7822
rect 25056 7410 25084 10406
rect 25148 10130 25176 10610
rect 25226 10568 25282 10577
rect 25226 10503 25282 10512
rect 25240 10470 25268 10503
rect 25228 10464 25280 10470
rect 25516 10452 25544 11070
rect 25516 10424 25636 10452
rect 25228 10406 25280 10412
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25148 8974 25176 10066
rect 25502 9888 25558 9897
rect 25502 9823 25558 9832
rect 25516 9722 25544 9823
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25410 9480 25466 9489
rect 25516 9450 25544 9522
rect 25410 9415 25412 9424
rect 25464 9415 25466 9424
rect 25504 9444 25556 9450
rect 25412 9386 25464 9392
rect 25504 9386 25556 9392
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25332 8809 25360 8842
rect 25318 8800 25374 8809
rect 25318 8735 25374 8744
rect 25608 8634 25636 10424
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25148 7002 25176 8570
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 24780 6458 24808 6734
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24872 6254 24900 6734
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24596 6118 24624 6190
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24596 5778 24624 6054
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 24492 5296 24544 5302
rect 24492 5238 24544 5244
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23952 2514 23980 2994
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23664 2032 23716 2038
rect 23664 1974 23716 1980
rect 20904 1352 20956 1358
rect 20904 1294 20956 1300
rect 21088 1352 21140 1358
rect 21088 1294 21140 1300
rect 22284 1352 22336 1358
rect 22284 1294 22336 1300
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 20628 1216 20680 1222
rect 20628 1158 20680 1164
rect 21100 1018 21128 1294
rect 21788 1116 22096 1125
rect 21788 1114 21794 1116
rect 21850 1114 21874 1116
rect 21930 1114 21954 1116
rect 22010 1114 22034 1116
rect 22090 1114 22096 1116
rect 21850 1062 21852 1114
rect 22032 1062 22034 1114
rect 21788 1060 21794 1062
rect 21850 1060 21874 1062
rect 21930 1060 21954 1062
rect 22010 1060 22034 1062
rect 22090 1060 22096 1062
rect 21788 1051 22096 1060
rect 21088 1012 21140 1018
rect 21088 954 21140 960
rect 23676 882 23704 1974
rect 23952 1970 23980 2450
rect 23940 1964 23992 1970
rect 23940 1906 23992 1912
rect 24044 1290 24072 3062
rect 24136 2774 24164 4678
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 25056 3738 25084 6598
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25148 5624 25176 6190
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25608 5914 25636 8434
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 25228 5636 25280 5642
rect 25148 5596 25228 5624
rect 25228 5578 25280 5584
rect 25240 5234 25268 5578
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24228 3126 24256 3334
rect 24216 3120 24268 3126
rect 24216 3062 24268 3068
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24136 2746 24256 2774
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 24136 2038 24164 2586
rect 24228 2038 24256 2746
rect 24872 2378 24900 2790
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24872 2038 24900 2314
rect 24124 2032 24176 2038
rect 24124 1974 24176 1980
rect 24216 2032 24268 2038
rect 24216 1974 24268 1980
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 25056 1290 25084 3674
rect 25608 3466 25636 4422
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25700 2446 25728 25162
rect 26988 24206 27016 25230
rect 27252 25220 27304 25226
rect 27252 25162 27304 25168
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 26068 22982 26096 23462
rect 27264 22982 27292 25162
rect 27528 25152 27580 25158
rect 27528 25094 27580 25100
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25976 21622 26004 21966
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 25976 20942 26004 21558
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25976 20534 26004 20878
rect 25964 20528 26016 20534
rect 25964 20470 26016 20476
rect 25976 19854 26004 20470
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25780 19780 25832 19786
rect 25780 19722 25832 19728
rect 25792 15502 25820 19722
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25976 18834 26004 19110
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25884 17202 25912 17614
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25884 16114 25912 17138
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25780 15496 25832 15502
rect 25780 15438 25832 15444
rect 25792 14074 25820 15438
rect 26068 14346 26096 22918
rect 27264 22681 27292 22918
rect 27250 22672 27306 22681
rect 27250 22607 27306 22616
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26160 17270 26188 21830
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26344 18698 26372 19110
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 26056 14340 26108 14346
rect 26056 14282 26108 14288
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 26160 14006 26188 15370
rect 26252 14006 26280 16458
rect 26344 16250 26372 18634
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26436 15706 26464 17478
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26344 15026 26372 15438
rect 26528 15094 26556 20742
rect 26896 18358 26924 21898
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26884 18352 26936 18358
rect 26884 18294 26936 18300
rect 26988 17746 27016 19790
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26620 15434 26648 15846
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 26516 15088 26568 15094
rect 26516 15030 26568 15036
rect 26332 15020 26384 15026
rect 26384 14980 26464 15008
rect 26332 14962 26384 14968
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26252 13530 26280 13942
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25884 10810 25912 13126
rect 26148 12640 26200 12646
rect 26146 12608 26148 12617
rect 26200 12608 26202 12617
rect 26146 12543 26202 12552
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25792 9178 25820 10202
rect 25884 9994 25912 10746
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25976 9602 26004 11222
rect 26056 11076 26108 11082
rect 26056 11018 26108 11024
rect 26068 9674 26096 11018
rect 26160 11014 26188 11698
rect 26344 11694 26372 13874
rect 26436 13394 26464 14980
rect 26528 14482 26556 15030
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26620 13258 26648 15370
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26608 13252 26660 13258
rect 26608 13194 26660 13200
rect 26514 12200 26570 12209
rect 26514 12135 26570 12144
rect 26528 12102 26556 12135
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26422 11792 26478 11801
rect 26422 11727 26478 11736
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26252 10169 26280 10542
rect 26238 10160 26294 10169
rect 26238 10095 26294 10104
rect 26436 9674 26464 11727
rect 26068 9646 26280 9674
rect 25976 9574 26188 9602
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25792 7886 25820 9114
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25884 7528 25912 8570
rect 25792 7500 25912 7528
rect 25792 4486 25820 7500
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25780 4480 25832 4486
rect 25780 4422 25832 4428
rect 25884 4146 25912 7346
rect 25976 4826 26004 9454
rect 26068 6458 26096 9454
rect 26160 6610 26188 9574
rect 26252 7002 26280 9646
rect 26344 9646 26464 9674
rect 26344 9586 26372 9646
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26528 9382 26556 12038
rect 26620 11898 26648 12038
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26712 9489 26740 14010
rect 26804 12434 26832 14758
rect 26896 12850 26924 16934
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26988 16114 27016 16594
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26988 14482 27016 16050
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 27080 14346 27108 16390
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 13802 27108 14282
rect 27068 13796 27120 13802
rect 27068 13738 27120 13744
rect 26884 12844 26936 12850
rect 26884 12786 26936 12792
rect 26804 12406 27016 12434
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26884 11824 26936 11830
rect 26884 11766 26936 11772
rect 26804 10266 26832 11766
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 26698 9480 26754 9489
rect 26698 9415 26754 9424
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26516 7812 26568 7818
rect 26516 7754 26568 7760
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26252 6730 26280 6938
rect 26344 6866 26372 7686
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26528 6798 26556 7754
rect 26620 7546 26648 8842
rect 26712 7886 26740 8910
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26712 6866 26740 7822
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26516 6792 26568 6798
rect 26422 6760 26478 6769
rect 26240 6724 26292 6730
rect 26516 6734 26568 6740
rect 26422 6695 26478 6704
rect 26240 6666 26292 6672
rect 26160 6582 26280 6610
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 26252 5370 26280 6582
rect 26436 6458 26464 6695
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26516 5704 26568 5710
rect 26516 5646 26568 5652
rect 26528 5574 26556 5646
rect 26804 5642 26832 10202
rect 26896 10062 26924 11766
rect 26988 10146 27016 12406
rect 27172 11898 27200 18566
rect 27356 17898 27384 24074
rect 27540 21962 27568 25094
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 27356 17870 27568 17898
rect 27540 17542 27568 17870
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27344 12436 27396 12442
rect 27448 12434 27476 15302
rect 27540 13870 27568 17478
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28356 14272 28408 14278
rect 28356 14214 28408 14220
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27396 12406 27476 12434
rect 27816 12434 27844 13194
rect 27816 12406 27936 12434
rect 27344 12378 27396 12384
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27068 11688 27120 11694
rect 27068 11630 27120 11636
rect 27080 10606 27108 11630
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27068 10600 27120 10606
rect 27068 10542 27120 10548
rect 26988 10118 27108 10146
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26884 9920 26936 9926
rect 26884 9862 26936 9868
rect 26792 5636 26844 5642
rect 26792 5578 26844 5584
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25792 1970 25820 4082
rect 25976 2446 26004 4762
rect 26436 4690 26464 5170
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26436 3942 26464 4626
rect 26528 4622 26556 5510
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26436 3602 26464 3878
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26896 3534 26924 9862
rect 26988 8974 27016 9998
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27080 8294 27108 10118
rect 27172 8906 27200 10610
rect 27264 9178 27292 11698
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27252 9172 27304 9178
rect 27252 9114 27304 9120
rect 27160 8900 27212 8906
rect 27160 8842 27212 8848
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27356 7818 27384 11222
rect 27448 10674 27476 12406
rect 27526 11792 27582 11801
rect 27526 11727 27528 11736
rect 27580 11727 27582 11736
rect 27528 11698 27580 11704
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27528 10804 27580 10810
rect 27528 10746 27580 10752
rect 27540 10713 27568 10746
rect 27526 10704 27582 10713
rect 27436 10668 27488 10674
rect 27526 10639 27582 10648
rect 27436 10610 27488 10616
rect 27724 9625 27752 11494
rect 27710 9616 27766 9625
rect 27710 9551 27766 9560
rect 27908 9450 27936 12406
rect 28368 12238 28396 14214
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 27896 9444 27948 9450
rect 27896 9386 27948 9392
rect 27908 8090 27936 9386
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27344 7812 27396 7818
rect 27344 7754 27396 7760
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27172 5166 27200 7142
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 27804 5296 27856 5302
rect 27804 5238 27856 5244
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27172 4282 27200 5102
rect 27816 4826 27844 5238
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 26976 3596 27028 3602
rect 26976 3538 27028 3544
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 26988 2514 27016 3538
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 26976 2508 27028 2514
rect 26976 2450 27028 2456
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25780 1964 25832 1970
rect 25780 1906 25832 1912
rect 25261 1660 25569 1669
rect 25261 1658 25267 1660
rect 25323 1658 25347 1660
rect 25403 1658 25427 1660
rect 25483 1658 25507 1660
rect 25563 1658 25569 1660
rect 25323 1606 25325 1658
rect 25505 1606 25507 1658
rect 25261 1604 25267 1606
rect 25323 1604 25347 1606
rect 25403 1604 25427 1606
rect 25483 1604 25507 1606
rect 25563 1604 25569 1606
rect 25261 1595 25569 1604
rect 24032 1284 24084 1290
rect 24032 1226 24084 1232
rect 25044 1284 25096 1290
rect 25044 1226 25096 1232
rect 25792 1222 25820 1906
rect 25964 1896 26016 1902
rect 25964 1838 26016 1844
rect 25976 1562 26004 1838
rect 25964 1556 26016 1562
rect 25964 1498 26016 1504
rect 26988 1358 27016 2450
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 26976 1352 27028 1358
rect 26976 1294 27028 1300
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 25780 1216 25832 1222
rect 25780 1158 25832 1164
rect 23768 1018 23796 1158
rect 28734 1116 29042 1125
rect 28734 1114 28740 1116
rect 28796 1114 28820 1116
rect 28876 1114 28900 1116
rect 28956 1114 28980 1116
rect 29036 1114 29042 1116
rect 28796 1062 28798 1114
rect 28978 1062 28980 1114
rect 28734 1060 28740 1062
rect 28796 1060 28820 1062
rect 28876 1060 28900 1062
rect 28956 1060 28980 1062
rect 29036 1060 29042 1062
rect 28734 1051 29042 1060
rect 23756 1012 23808 1018
rect 23756 954 23808 960
rect 20168 876 20220 882
rect 20168 818 20220 824
rect 23664 876 23716 882
rect 23664 818 23716 824
rect 5354 776 5410 785
rect 5354 711 5410 720
<< via2 >>
rect 7902 32666 7958 32668
rect 7982 32666 8038 32668
rect 8062 32666 8118 32668
rect 8142 32666 8198 32668
rect 7902 32614 7948 32666
rect 7948 32614 7958 32666
rect 7982 32614 8012 32666
rect 8012 32614 8024 32666
rect 8024 32614 8038 32666
rect 8062 32614 8076 32666
rect 8076 32614 8088 32666
rect 8088 32614 8118 32666
rect 8142 32614 8152 32666
rect 8152 32614 8198 32666
rect 7902 32612 7958 32614
rect 7982 32612 8038 32614
rect 8062 32612 8118 32614
rect 8142 32612 8198 32614
rect 14848 32666 14904 32668
rect 14928 32666 14984 32668
rect 15008 32666 15064 32668
rect 15088 32666 15144 32668
rect 14848 32614 14894 32666
rect 14894 32614 14904 32666
rect 14928 32614 14958 32666
rect 14958 32614 14970 32666
rect 14970 32614 14984 32666
rect 15008 32614 15022 32666
rect 15022 32614 15034 32666
rect 15034 32614 15064 32666
rect 15088 32614 15098 32666
rect 15098 32614 15144 32666
rect 14848 32612 14904 32614
rect 14928 32612 14984 32614
rect 15008 32612 15064 32614
rect 15088 32612 15144 32614
rect 21794 32666 21850 32668
rect 21874 32666 21930 32668
rect 21954 32666 22010 32668
rect 22034 32666 22090 32668
rect 21794 32614 21840 32666
rect 21840 32614 21850 32666
rect 21874 32614 21904 32666
rect 21904 32614 21916 32666
rect 21916 32614 21930 32666
rect 21954 32614 21968 32666
rect 21968 32614 21980 32666
rect 21980 32614 22010 32666
rect 22034 32614 22044 32666
rect 22044 32614 22090 32666
rect 21794 32612 21850 32614
rect 21874 32612 21930 32614
rect 21954 32612 22010 32614
rect 22034 32612 22090 32614
rect 28740 32666 28796 32668
rect 28820 32666 28876 32668
rect 28900 32666 28956 32668
rect 28980 32666 29036 32668
rect 28740 32614 28786 32666
rect 28786 32614 28796 32666
rect 28820 32614 28850 32666
rect 28850 32614 28862 32666
rect 28862 32614 28876 32666
rect 28900 32614 28914 32666
rect 28914 32614 28926 32666
rect 28926 32614 28956 32666
rect 28980 32614 28990 32666
rect 28990 32614 29036 32666
rect 28740 32612 28796 32614
rect 28820 32612 28876 32614
rect 28900 32612 28956 32614
rect 28980 32612 29036 32614
rect 2778 32272 2834 32328
rect 846 24132 902 24168
rect 846 24112 848 24132
rect 848 24112 900 24132
rect 900 24112 902 24132
rect 662 15952 718 16008
rect 570 13912 626 13968
rect 754 11872 810 11928
rect 846 9832 902 9888
rect 938 7828 940 7848
rect 940 7828 992 7848
rect 992 7828 994 7848
rect 938 7792 994 7828
rect 1306 3712 1362 3768
rect 1950 22092 2006 22128
rect 1950 22072 1952 22092
rect 1952 22072 2004 22092
rect 2004 22072 2006 22092
rect 4429 32122 4485 32124
rect 4509 32122 4565 32124
rect 4589 32122 4645 32124
rect 4669 32122 4725 32124
rect 4429 32070 4475 32122
rect 4475 32070 4485 32122
rect 4509 32070 4539 32122
rect 4539 32070 4551 32122
rect 4551 32070 4565 32122
rect 4589 32070 4603 32122
rect 4603 32070 4615 32122
rect 4615 32070 4645 32122
rect 4669 32070 4679 32122
rect 4679 32070 4725 32122
rect 4429 32068 4485 32070
rect 4509 32068 4565 32070
rect 4589 32068 4645 32070
rect 4669 32068 4725 32070
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 3974 30268 3976 30288
rect 3976 30268 4028 30288
rect 4028 30268 4030 30288
rect 3974 30232 4030 30268
rect 4066 28192 4122 28248
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 1766 5752 1822 5808
rect 3054 15544 3110 15600
rect 2686 6840 2742 6896
rect 3146 5072 3202 5128
rect 3054 4004 3110 4040
rect 3054 3984 3056 4004
rect 3056 3984 3108 4004
rect 3108 3984 3110 4004
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4342 26152 4398 26208
rect 4066 20032 4122 20088
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4710 23840 4766 23896
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4986 23724 5042 23760
rect 4986 23704 4988 23724
rect 4988 23704 5040 23724
rect 5040 23704 5042 23724
rect 5354 26288 5410 26344
rect 5262 23840 5318 23896
rect 5170 23704 5226 23760
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 3882 17992 3938 18048
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 5630 19352 5686 19408
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4526 15952 4582 16008
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 5998 18808 6054 18864
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 6274 20868 6330 20904
rect 6274 20848 6276 20868
rect 6276 20848 6328 20868
rect 6328 20848 6330 20868
rect 6550 19624 6606 19680
rect 6550 19372 6606 19408
rect 6550 19352 6552 19372
rect 6552 19352 6604 19372
rect 6604 19352 6606 19372
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 6274 17448 6330 17504
rect 6274 16108 6330 16144
rect 6274 16088 6276 16108
rect 6276 16088 6328 16108
rect 6328 16088 6330 16108
rect 6090 15544 6146 15600
rect 5078 12164 5134 12200
rect 5078 12144 5080 12164
rect 5080 12144 5132 12164
rect 5132 12144 5134 12164
rect 5262 12144 5318 12200
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 4802 6976 4858 7032
rect 5262 11092 5264 11112
rect 5264 11092 5316 11112
rect 5316 11092 5318 11112
rect 5262 11056 5318 11092
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7102 20440 7158 20496
rect 7102 18708 7104 18728
rect 7104 18708 7156 18728
rect 7156 18708 7158 18728
rect 7102 18672 7158 18708
rect 7470 20848 7526 20904
rect 6918 15952 6974 16008
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7470 17620 7472 17640
rect 7472 17620 7524 17640
rect 7524 17620 7526 17640
rect 7470 17584 7526 17620
rect 6182 9696 6238 9752
rect 6642 11056 6698 11112
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 8114 16088 8170 16144
rect 8758 18808 8814 18864
rect 8390 15408 8446 15464
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 8022 14764 8024 14784
rect 8024 14764 8076 14784
rect 8076 14764 8078 14784
rect 8022 14728 8078 14764
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 3330 2644 3386 2680
rect 3330 2624 3332 2644
rect 3332 2624 3384 2644
rect 3384 2624 3386 2644
rect 3422 1944 3478 2000
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 8298 13776 8354 13832
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 8942 16516 8998 16552
rect 8942 16496 8944 16516
rect 8944 16496 8996 16516
rect 8996 16496 8998 16516
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 8206 11076 8262 11112
rect 8206 11056 8208 11076
rect 8208 11056 8260 11076
rect 8260 11056 8262 11076
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 11375 32122 11431 32124
rect 11455 32122 11511 32124
rect 11535 32122 11591 32124
rect 11615 32122 11671 32124
rect 11375 32070 11421 32122
rect 11421 32070 11431 32122
rect 11455 32070 11485 32122
rect 11485 32070 11497 32122
rect 11497 32070 11511 32122
rect 11535 32070 11549 32122
rect 11549 32070 11561 32122
rect 11561 32070 11591 32122
rect 11615 32070 11625 32122
rect 11625 32070 11671 32122
rect 11375 32068 11431 32070
rect 11455 32068 11511 32070
rect 11535 32068 11591 32070
rect 11615 32068 11671 32070
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 9126 16768 9182 16824
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 9770 19624 9826 19680
rect 9770 19252 9772 19272
rect 9772 19252 9824 19272
rect 9824 19252 9826 19272
rect 9770 19216 9826 19252
rect 9494 18572 9496 18592
rect 9496 18572 9548 18592
rect 9548 18572 9550 18592
rect 9494 18536 9550 18572
rect 10230 19896 10286 19952
rect 10138 19488 10194 19544
rect 9494 17604 9550 17640
rect 9494 17584 9496 17604
rect 9496 17584 9548 17604
rect 9548 17584 9550 17604
rect 9310 16632 9366 16688
rect 9586 16768 9642 16824
rect 8942 15136 8998 15192
rect 9402 15544 9458 15600
rect 9310 15408 9366 15464
rect 9678 16088 9734 16144
rect 9310 14728 9366 14784
rect 9126 14320 9182 14376
rect 9586 14864 9642 14920
rect 9586 14728 9642 14784
rect 9494 14356 9496 14376
rect 9496 14356 9548 14376
rect 9548 14356 9550 14376
rect 9494 14320 9550 14356
rect 9218 12144 9274 12200
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 9678 13268 9680 13288
rect 9680 13268 9732 13288
rect 9732 13268 9734 13288
rect 9678 13232 9734 13268
rect 9678 12960 9734 13016
rect 9586 12844 9642 12880
rect 9586 12824 9588 12844
rect 9588 12824 9640 12844
rect 9640 12824 9642 12844
rect 8298 5752 8354 5808
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 9402 5480 9458 5536
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 18321 32122 18377 32124
rect 18401 32122 18457 32124
rect 18481 32122 18537 32124
rect 18561 32122 18617 32124
rect 18321 32070 18367 32122
rect 18367 32070 18377 32122
rect 18401 32070 18431 32122
rect 18431 32070 18443 32122
rect 18443 32070 18457 32122
rect 18481 32070 18495 32122
rect 18495 32070 18507 32122
rect 18507 32070 18537 32122
rect 18561 32070 18571 32122
rect 18571 32070 18617 32122
rect 18321 32068 18377 32070
rect 18401 32068 18457 32070
rect 18481 32068 18537 32070
rect 18561 32068 18617 32070
rect 25267 32122 25323 32124
rect 25347 32122 25403 32124
rect 25427 32122 25483 32124
rect 25507 32122 25563 32124
rect 25267 32070 25313 32122
rect 25313 32070 25323 32122
rect 25347 32070 25377 32122
rect 25377 32070 25389 32122
rect 25389 32070 25403 32122
rect 25427 32070 25441 32122
rect 25441 32070 25453 32122
rect 25453 32070 25483 32122
rect 25507 32070 25517 32122
rect 25517 32070 25563 32122
rect 25267 32068 25323 32070
rect 25347 32068 25403 32070
rect 25427 32068 25483 32070
rect 25507 32068 25563 32070
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 10230 14456 10286 14512
rect 10046 6840 10102 6896
rect 2870 1672 2926 1728
rect 4429 1658 4485 1660
rect 4509 1658 4565 1660
rect 4589 1658 4645 1660
rect 4669 1658 4725 1660
rect 4429 1606 4475 1658
rect 4475 1606 4485 1658
rect 4509 1606 4539 1658
rect 4539 1606 4551 1658
rect 4551 1606 4565 1658
rect 4589 1606 4603 1658
rect 4603 1606 4615 1658
rect 4615 1606 4645 1658
rect 4669 1606 4679 1658
rect 4679 1606 4725 1658
rect 4429 1604 4485 1606
rect 4509 1604 4565 1606
rect 4589 1604 4645 1606
rect 4669 1604 4725 1606
rect 3330 1264 3386 1320
rect 11058 19488 11114 19544
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11610 20340 11612 20360
rect 11612 20340 11664 20360
rect 11664 20340 11666 20360
rect 11610 20304 11666 20340
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11426 19896 11482 19952
rect 11242 19796 11244 19816
rect 11244 19796 11296 19816
rect 11296 19796 11298 19816
rect 11242 19760 11298 19796
rect 11334 19660 11336 19680
rect 11336 19660 11388 19680
rect 11388 19660 11390 19680
rect 11334 19624 11390 19660
rect 10874 15544 10930 15600
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11150 16088 11206 16144
rect 11702 16632 11758 16688
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11610 15272 11666 15328
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 13174 24792 13230 24848
rect 12162 19624 12218 19680
rect 12346 19488 12402 19544
rect 11794 14456 11850 14512
rect 10506 6160 10562 6216
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11886 7656 11942 7712
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 15842 25200 15898 25256
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14830 24812 14886 24848
rect 14830 24792 14832 24812
rect 14832 24792 14884 24812
rect 14884 24792 14886 24812
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 12714 14220 12716 14240
rect 12716 14220 12768 14240
rect 12768 14220 12770 14240
rect 12714 14184 12770 14220
rect 12898 17448 12954 17504
rect 12438 13368 12494 13424
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 12806 12144 12862 12200
rect 12530 8880 12586 8936
rect 12438 7656 12494 7712
rect 13726 19216 13782 19272
rect 13266 12144 13322 12200
rect 12162 4528 12218 4584
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 11375 1658 11431 1660
rect 11455 1658 11511 1660
rect 11535 1658 11591 1660
rect 11615 1658 11671 1660
rect 11375 1606 11421 1658
rect 11421 1606 11431 1658
rect 11455 1606 11485 1658
rect 11485 1606 11497 1658
rect 11497 1606 11511 1658
rect 11535 1606 11549 1658
rect 11549 1606 11561 1658
rect 11561 1606 11591 1658
rect 11615 1606 11625 1658
rect 11625 1606 11671 1658
rect 11375 1604 11431 1606
rect 11455 1604 11511 1606
rect 11535 1604 11591 1606
rect 11615 1604 11671 1606
rect 11978 1300 11980 1320
rect 11980 1300 12032 1320
rect 12032 1300 12034 1320
rect 11978 1264 12034 1300
rect 12438 5244 12440 5264
rect 12440 5244 12492 5264
rect 12492 5244 12494 5264
rect 12438 5208 12494 5244
rect 13818 12552 13874 12608
rect 13726 10512 13782 10568
rect 13634 9152 13690 9208
rect 13082 7420 13084 7440
rect 13084 7420 13136 7440
rect 13136 7420 13138 7440
rect 13082 7384 13138 7420
rect 12990 5616 13046 5672
rect 12898 5208 12954 5264
rect 13082 5208 13138 5264
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14370 17484 14372 17504
rect 14372 17484 14424 17504
rect 14424 17484 14426 17504
rect 14370 17448 14426 17484
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 15290 17584 15346 17640
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14462 13504 14518 13560
rect 14094 11600 14150 11656
rect 14002 10376 14058 10432
rect 12990 3032 13046 3088
rect 12438 1400 12494 1456
rect 13726 6840 13782 6896
rect 14278 8200 14334 8256
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 15474 13776 15530 13832
rect 15382 13504 15438 13560
rect 15842 20712 15898 20768
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 15658 13504 15714 13560
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 15014 11756 15070 11792
rect 15014 11736 15016 11756
rect 15016 11736 15068 11756
rect 15068 11736 15070 11756
rect 15290 11600 15346 11656
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14554 7112 14610 7168
rect 15290 8916 15292 8936
rect 15292 8916 15344 8936
rect 15344 8916 15346 8936
rect 15290 8880 15346 8916
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 15658 12844 15714 12880
rect 15934 13232 15990 13288
rect 16118 13368 16174 13424
rect 15658 12824 15660 12844
rect 15660 12824 15712 12844
rect 15712 12824 15714 12844
rect 15934 11736 15990 11792
rect 16302 16496 16358 16552
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 16394 13504 16450 13560
rect 15658 9016 15714 9072
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 15014 7248 15070 7304
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14830 6296 14886 6352
rect 14922 6160 14978 6216
rect 15014 6024 15070 6080
rect 15014 5752 15070 5808
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 15014 3052 15070 3088
rect 15014 3032 15016 3052
rect 15016 3032 15068 3052
rect 15068 3032 15070 3052
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 16486 11192 16542 11248
rect 15842 7384 15898 7440
rect 15842 6740 15844 6760
rect 15844 6740 15896 6760
rect 15896 6740 15898 6760
rect 15842 6704 15898 6740
rect 16670 13912 16726 13968
rect 16946 13096 17002 13152
rect 16854 11056 16910 11112
rect 16670 10376 16726 10432
rect 16670 9968 16726 10024
rect 16946 9016 17002 9072
rect 17958 18028 17960 18048
rect 17960 18028 18012 18048
rect 18012 18028 18014 18048
rect 17314 13776 17370 13832
rect 17958 17992 18014 18028
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18234 19896 18290 19952
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 17866 16652 17922 16688
rect 17866 16632 17868 16652
rect 17868 16632 17920 16652
rect 17920 16632 17922 16652
rect 17498 12960 17554 13016
rect 18142 16360 18198 16416
rect 17774 12688 17830 12744
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18786 16788 18842 16824
rect 18786 16768 18788 16788
rect 18788 16768 18840 16788
rect 18840 16768 18842 16788
rect 18786 15952 18842 16008
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18326 15308 18328 15328
rect 18328 15308 18380 15328
rect 18380 15308 18382 15328
rect 18050 12688 18106 12744
rect 17958 12588 17960 12608
rect 17960 12588 18012 12608
rect 18012 12588 18014 12608
rect 17958 12552 18014 12588
rect 17866 11736 17922 11792
rect 17130 7420 17132 7440
rect 17132 7420 17184 7440
rect 17184 7420 17186 7440
rect 17130 7384 17186 7420
rect 17314 7112 17370 7168
rect 16578 5636 16634 5672
rect 16578 5616 16580 5636
rect 16580 5616 16632 5636
rect 16632 5616 16634 5636
rect 16118 1400 16174 1456
rect 17038 3032 17094 3088
rect 18142 12280 18198 12336
rect 18326 15272 18382 15308
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18326 13776 18382 13832
rect 18694 13932 18750 13968
rect 18694 13912 18696 13932
rect 18696 13912 18748 13932
rect 18748 13912 18750 13932
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 19338 16768 19394 16824
rect 19430 16396 19432 16416
rect 19432 16396 19484 16416
rect 19484 16396 19486 16416
rect 19430 16360 19486 16396
rect 19430 16224 19486 16280
rect 19154 15816 19210 15872
rect 18786 13096 18842 13152
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18142 10920 18198 10976
rect 18694 10376 18750 10432
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 17958 9152 18014 9208
rect 19246 15680 19302 15736
rect 19706 16088 19762 16144
rect 18142 9424 18198 9480
rect 18050 8744 18106 8800
rect 17958 8472 18014 8528
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18326 9016 18382 9072
rect 18050 8336 18106 8392
rect 18326 8492 18382 8528
rect 18326 8472 18328 8492
rect 18328 8472 18380 8492
rect 18380 8472 18382 8492
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18694 6724 18750 6760
rect 18694 6704 18696 6724
rect 18696 6704 18748 6724
rect 18748 6704 18750 6724
rect 17314 6160 17370 6216
rect 17774 6160 17830 6216
rect 17314 2624 17370 2680
rect 17314 2488 17370 2544
rect 17314 2252 17316 2272
rect 17316 2252 17368 2272
rect 17368 2252 17370 2272
rect 17314 2216 17370 2252
rect 17590 5208 17646 5264
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18418 5752 18474 5808
rect 17774 2624 17830 2680
rect 2226 856 2282 912
rect 7902 1114 7958 1116
rect 7982 1114 8038 1116
rect 8062 1114 8118 1116
rect 8142 1114 8198 1116
rect 7902 1062 7948 1114
rect 7948 1062 7958 1114
rect 7982 1062 8012 1114
rect 8012 1062 8024 1114
rect 8024 1062 8038 1114
rect 8062 1062 8076 1114
rect 8076 1062 8088 1114
rect 8088 1062 8118 1114
rect 8142 1062 8152 1114
rect 8152 1062 8198 1114
rect 7902 1060 7958 1062
rect 7982 1060 8038 1062
rect 8062 1060 8118 1062
rect 8142 1060 8198 1062
rect 14848 1114 14904 1116
rect 14928 1114 14984 1116
rect 15008 1114 15064 1116
rect 15088 1114 15144 1116
rect 14848 1062 14894 1114
rect 14894 1062 14904 1114
rect 14928 1062 14958 1114
rect 14958 1062 14970 1114
rect 14970 1062 14984 1114
rect 15008 1062 15022 1114
rect 15022 1062 15034 1114
rect 15034 1062 15064 1114
rect 15088 1062 15098 1114
rect 15098 1062 15144 1114
rect 14848 1060 14904 1062
rect 14928 1060 14984 1062
rect 15008 1060 15064 1062
rect 15088 1060 15144 1062
rect 18142 4548 18198 4584
rect 18142 4528 18144 4548
rect 18144 4528 18196 4548
rect 18196 4528 18198 4548
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 18326 2524 18328 2544
rect 18328 2524 18380 2544
rect 18380 2524 18382 2544
rect 18326 2488 18382 2524
rect 18878 8356 18934 8392
rect 18878 8336 18880 8356
rect 18880 8336 18932 8356
rect 18932 8336 18934 8356
rect 18321 1658 18377 1660
rect 18401 1658 18457 1660
rect 18481 1658 18537 1660
rect 18561 1658 18617 1660
rect 18321 1606 18367 1658
rect 18367 1606 18377 1658
rect 18401 1606 18431 1658
rect 18431 1606 18443 1658
rect 18443 1606 18457 1658
rect 18481 1606 18495 1658
rect 18495 1606 18507 1658
rect 18507 1606 18537 1658
rect 18561 1606 18571 1658
rect 18571 1606 18617 1658
rect 18321 1604 18377 1606
rect 18401 1604 18457 1606
rect 18481 1604 18537 1606
rect 18561 1604 18617 1606
rect 19522 12280 19578 12336
rect 19338 10140 19340 10160
rect 19340 10140 19392 10160
rect 19392 10140 19394 10160
rect 19338 10104 19394 10140
rect 19982 16224 20038 16280
rect 19706 13232 19762 13288
rect 19614 10240 19670 10296
rect 19614 10140 19616 10160
rect 19616 10140 19668 10160
rect 19668 10140 19670 10160
rect 19614 10104 19670 10140
rect 19522 9832 19578 9888
rect 19338 9696 19394 9752
rect 19522 9560 19578 9616
rect 19614 9288 19670 9344
rect 19338 8628 19394 8664
rect 19338 8608 19340 8628
rect 19340 8608 19392 8628
rect 19392 8608 19394 8628
rect 19430 8200 19486 8256
rect 19430 8064 19486 8120
rect 19706 8744 19762 8800
rect 19614 8336 19670 8392
rect 19890 12688 19946 12744
rect 20442 16632 20498 16688
rect 20074 15036 20076 15056
rect 20076 15036 20128 15056
rect 20128 15036 20130 15056
rect 20074 15000 20130 15036
rect 19982 12280 20038 12336
rect 20258 15816 20314 15872
rect 20718 15428 20774 15464
rect 20718 15408 20720 15428
rect 20720 15408 20772 15428
rect 20772 15408 20774 15428
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21270 16496 21326 16552
rect 21270 15952 21326 16008
rect 20258 13932 20314 13968
rect 20258 13912 20260 13932
rect 20260 13912 20312 13932
rect 20312 13912 20314 13932
rect 20258 13232 20314 13288
rect 20258 12280 20314 12336
rect 21178 14764 21180 14784
rect 21180 14764 21232 14784
rect 21232 14764 21234 14784
rect 21178 14728 21234 14764
rect 19890 11192 19946 11248
rect 19890 10648 19946 10704
rect 19890 10376 19946 10432
rect 19890 9696 19946 9752
rect 19890 9596 19892 9616
rect 19892 9596 19944 9616
rect 19944 9596 19946 9616
rect 19890 9560 19946 9596
rect 20626 11348 20682 11384
rect 20626 11328 20628 11348
rect 20628 11328 20680 11348
rect 20680 11328 20682 11348
rect 21178 12180 21180 12200
rect 21180 12180 21232 12200
rect 21232 12180 21234 12200
rect 21178 12144 21234 12180
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 22190 19352 22246 19408
rect 22190 18572 22192 18592
rect 22192 18572 22244 18592
rect 22244 18572 22246 18592
rect 22190 18536 22246 18572
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21914 15564 21970 15600
rect 21914 15544 21916 15564
rect 21916 15544 21968 15564
rect 21968 15544 21970 15564
rect 21730 15428 21786 15464
rect 21730 15408 21732 15428
rect 21732 15408 21784 15428
rect 21784 15408 21786 15428
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21454 11500 21456 11520
rect 21456 11500 21508 11520
rect 21508 11500 21510 11520
rect 21454 11464 21510 11500
rect 21454 11328 21510 11384
rect 20626 10512 20682 10568
rect 20994 10920 21050 10976
rect 21086 10376 21142 10432
rect 20626 9560 20682 9616
rect 20074 6840 20130 6896
rect 19798 6160 19854 6216
rect 20626 8900 20682 8936
rect 20626 8880 20628 8900
rect 20628 8880 20680 8900
rect 20680 8880 20682 8900
rect 20626 8608 20682 8664
rect 20994 9832 21050 9888
rect 20534 6724 20590 6760
rect 20534 6704 20536 6724
rect 20536 6704 20588 6724
rect 20588 6704 20590 6724
rect 18970 2216 19026 2272
rect 21086 7248 21142 7304
rect 21362 10104 21418 10160
rect 21362 9716 21418 9752
rect 21362 9696 21364 9716
rect 21364 9696 21416 9716
rect 21416 9696 21418 9716
rect 22650 16088 22706 16144
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 22190 13640 22246 13696
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 22742 15680 22798 15736
rect 23110 18536 23166 18592
rect 23386 19388 23388 19408
rect 23388 19388 23440 19408
rect 23440 19388 23442 19408
rect 23386 19352 23442 19388
rect 22834 15272 22890 15328
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 22190 10784 22246 10840
rect 21730 10240 21786 10296
rect 22098 10512 22154 10568
rect 22834 12688 22890 12744
rect 22374 10684 22376 10704
rect 22376 10684 22428 10704
rect 22428 10684 22430 10704
rect 22374 10648 22430 10684
rect 22742 12008 22798 12064
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21822 7828 21824 7848
rect 21824 7828 21876 7848
rect 21876 7828 21878 7848
rect 21822 7792 21878 7828
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 22282 8200 22338 8256
rect 22282 7928 22338 7984
rect 21822 6840 21878 6896
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 22466 10512 22522 10568
rect 22466 9832 22522 9888
rect 22650 9968 22706 10024
rect 22558 9696 22614 9752
rect 22834 10668 22890 10704
rect 22834 10648 22836 10668
rect 22836 10648 22888 10668
rect 22888 10648 22890 10668
rect 22282 6160 22338 6216
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 22742 9580 22798 9616
rect 22742 9560 22744 9580
rect 22744 9560 22796 9580
rect 22796 9560 22798 9580
rect 23202 16652 23258 16688
rect 23202 16632 23204 16652
rect 23204 16632 23256 16652
rect 23256 16632 23258 16652
rect 23110 11192 23166 11248
rect 23478 16224 23534 16280
rect 23478 16108 23534 16144
rect 23478 16088 23480 16108
rect 23480 16088 23532 16108
rect 23532 16088 23534 16108
rect 23754 16224 23810 16280
rect 23294 11056 23350 11112
rect 23202 10376 23258 10432
rect 22742 7928 22798 7984
rect 22558 6160 22614 6216
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 21086 1400 21142 1456
rect 23386 10784 23442 10840
rect 23386 7792 23442 7848
rect 24398 18028 24400 18048
rect 24400 18028 24452 18048
rect 24452 18028 24454 18048
rect 24398 17992 24454 18028
rect 24122 15408 24178 15464
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25962 25336 26018 25392
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 24122 9696 24178 9752
rect 24030 9016 24086 9072
rect 23938 8880 23994 8936
rect 24306 11736 24362 11792
rect 24306 11328 24362 11384
rect 24398 11192 24454 11248
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 24490 10104 24546 10160
rect 24398 8744 24454 8800
rect 24306 6704 24362 6760
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25042 12008 25098 12064
rect 25042 11892 25098 11928
rect 25042 11872 25044 11892
rect 25044 11872 25096 11892
rect 25096 11872 25098 11892
rect 24766 11464 24822 11520
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 24766 10104 24822 10160
rect 25226 10512 25282 10568
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 25502 9832 25558 9888
rect 25410 9444 25466 9480
rect 25410 9424 25412 9444
rect 25412 9424 25464 9444
rect 25464 9424 25466 9444
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25318 8744 25374 8800
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 21794 1114 21850 1116
rect 21874 1114 21930 1116
rect 21954 1114 22010 1116
rect 22034 1114 22090 1116
rect 21794 1062 21840 1114
rect 21840 1062 21850 1114
rect 21874 1062 21904 1114
rect 21904 1062 21916 1114
rect 21916 1062 21930 1114
rect 21954 1062 21968 1114
rect 21968 1062 21980 1114
rect 21980 1062 22010 1114
rect 22034 1062 22044 1114
rect 22044 1062 22090 1114
rect 21794 1060 21850 1062
rect 21874 1060 21930 1062
rect 21954 1060 22010 1062
rect 22034 1060 22090 1062
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 27250 22616 27306 22672
rect 26146 12588 26148 12608
rect 26148 12588 26200 12608
rect 26200 12588 26202 12608
rect 26146 12552 26202 12588
rect 26514 12144 26570 12200
rect 26422 11736 26478 11792
rect 26238 10104 26294 10160
rect 26698 9424 26754 9480
rect 26422 6704 26478 6760
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 27526 11756 27582 11792
rect 27526 11736 27528 11756
rect 27528 11736 27580 11756
rect 27580 11736 27582 11756
rect 27526 10648 27582 10704
rect 27710 9560 27766 9616
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 25267 1658 25323 1660
rect 25347 1658 25403 1660
rect 25427 1658 25483 1660
rect 25507 1658 25563 1660
rect 25267 1606 25313 1658
rect 25313 1606 25323 1658
rect 25347 1606 25377 1658
rect 25377 1606 25389 1658
rect 25389 1606 25403 1658
rect 25427 1606 25441 1658
rect 25441 1606 25453 1658
rect 25453 1606 25483 1658
rect 25507 1606 25517 1658
rect 25517 1606 25563 1658
rect 25267 1604 25323 1606
rect 25347 1604 25403 1606
rect 25427 1604 25483 1606
rect 25507 1604 25563 1606
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 28740 1114 28796 1116
rect 28820 1114 28876 1116
rect 28900 1114 28956 1116
rect 28980 1114 29036 1116
rect 28740 1062 28786 1114
rect 28786 1062 28796 1114
rect 28820 1062 28850 1114
rect 28850 1062 28862 1114
rect 28862 1062 28876 1114
rect 28900 1062 28914 1114
rect 28914 1062 28926 1114
rect 28926 1062 28956 1114
rect 28980 1062 28990 1114
rect 28990 1062 29036 1114
rect 28740 1060 28796 1062
rect 28820 1060 28876 1062
rect 28900 1060 28956 1062
rect 28980 1060 29036 1062
rect 5354 720 5410 776
<< metal3 >>
rect 7892 32672 8208 32673
rect 7892 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8208 32672
rect 7892 32607 8208 32608
rect 14838 32672 15154 32673
rect 14838 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15154 32672
rect 14838 32607 15154 32608
rect 21784 32672 22100 32673
rect 21784 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22100 32672
rect 21784 32607 22100 32608
rect 28730 32672 29046 32673
rect 28730 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29046 32672
rect 28730 32607 29046 32608
rect 0 32330 400 32360
rect 2773 32330 2839 32333
rect 0 32328 2839 32330
rect 0 32272 2778 32328
rect 2834 32272 2839 32328
rect 0 32270 2839 32272
rect 0 32240 400 32270
rect 2773 32267 2839 32270
rect 4419 32128 4735 32129
rect 4419 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4735 32128
rect 4419 32063 4735 32064
rect 11365 32128 11681 32129
rect 11365 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11681 32128
rect 11365 32063 11681 32064
rect 18311 32128 18627 32129
rect 18311 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18627 32128
rect 18311 32063 18627 32064
rect 25257 32128 25573 32129
rect 25257 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25573 32128
rect 25257 32063 25573 32064
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 4419 31040 4735 31041
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 28730 30431 29046 30432
rect 0 30290 400 30320
rect 3969 30290 4035 30293
rect 0 30288 4035 30290
rect 0 30232 3974 30288
rect 4030 30232 4035 30288
rect 0 30230 4035 30232
rect 0 30200 400 30230
rect 3969 30227 4035 30230
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 7892 28320 8208 28321
rect 0 28250 400 28280
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 4061 28250 4127 28253
rect 0 28248 4127 28250
rect 0 28192 4066 28248
rect 4122 28192 4127 28248
rect 0 28190 4127 28192
rect 0 28160 400 28190
rect 4061 28187 4127 28190
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 5349 26346 5415 26349
rect 7414 26346 7420 26348
rect 5349 26344 7420 26346
rect 5349 26288 5354 26344
rect 5410 26288 7420 26344
rect 5349 26286 7420 26288
rect 5349 26283 5415 26286
rect 7414 26284 7420 26286
rect 7484 26284 7490 26348
rect 0 26210 400 26240
rect 4337 26210 4403 26213
rect 0 26208 4403 26210
rect 0 26152 4342 26208
rect 4398 26152 4403 26208
rect 0 26150 4403 26152
rect 0 26120 400 26150
rect 4337 26147 4403 26150
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 10174 25332 10180 25396
rect 10244 25394 10250 25396
rect 25957 25394 26023 25397
rect 10244 25392 26023 25394
rect 10244 25336 25962 25392
rect 26018 25336 26023 25392
rect 10244 25334 26023 25336
rect 10244 25332 10250 25334
rect 25957 25331 26023 25334
rect 13118 25196 13124 25260
rect 13188 25258 13194 25260
rect 15837 25258 15903 25261
rect 13188 25256 15903 25258
rect 13188 25200 15842 25256
rect 15898 25200 15903 25256
rect 13188 25198 15903 25200
rect 13188 25196 13194 25198
rect 15837 25195 15903 25198
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 12934 24788 12940 24852
rect 13004 24850 13010 24852
rect 13169 24850 13235 24853
rect 14825 24850 14891 24853
rect 13004 24848 14891 24850
rect 13004 24792 13174 24848
rect 13230 24792 14830 24848
rect 14886 24792 14891 24848
rect 13004 24790 14891 24792
rect 13004 24788 13010 24790
rect 13169 24787 13235 24790
rect 14825 24787 14891 24790
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 0 24170 400 24200
rect 841 24170 907 24173
rect 0 24168 907 24170
rect 0 24112 846 24168
rect 902 24112 907 24168
rect 0 24110 907 24112
rect 0 24080 400 24110
rect 841 24107 907 24110
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 4705 23898 4771 23901
rect 5257 23898 5323 23901
rect 4705 23896 5323 23898
rect 4705 23840 4710 23896
rect 4766 23840 5262 23896
rect 5318 23840 5323 23896
rect 4705 23838 5323 23840
rect 4705 23835 4771 23838
rect 5257 23835 5323 23838
rect 4981 23762 5047 23765
rect 5165 23762 5231 23765
rect 4981 23760 5231 23762
rect 4981 23704 4986 23760
rect 5042 23704 5170 23760
rect 5226 23704 5231 23760
rect 4981 23702 5231 23704
rect 4981 23699 5047 23702
rect 5165 23699 5231 23702
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 21398 22612 21404 22676
rect 21468 22674 21474 22676
rect 27245 22674 27311 22677
rect 21468 22672 27311 22674
rect 21468 22616 27250 22672
rect 27306 22616 27311 22672
rect 21468 22614 27311 22616
rect 21468 22612 21474 22614
rect 27245 22611 27311 22614
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 0 22130 400 22160
rect 1945 22130 2011 22133
rect 0 22128 2011 22130
rect 0 22072 1950 22128
rect 2006 22072 2011 22128
rect 0 22070 2011 22072
rect 0 22040 400 22070
rect 1945 22067 2011 22070
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 6269 20906 6335 20909
rect 7465 20906 7531 20909
rect 6269 20904 7531 20906
rect 6269 20848 6274 20904
rect 6330 20848 7470 20904
rect 7526 20848 7531 20904
rect 6269 20846 7531 20848
rect 6269 20843 6335 20846
rect 7465 20843 7531 20846
rect 15837 20772 15903 20773
rect 15837 20768 15884 20772
rect 15948 20770 15954 20772
rect 15837 20712 15842 20768
rect 15837 20708 15884 20712
rect 15948 20710 15994 20770
rect 15948 20708 15954 20710
rect 15837 20707 15903 20708
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 7097 20498 7163 20501
rect 7230 20498 7236 20500
rect 7097 20496 7236 20498
rect 7097 20440 7102 20496
rect 7158 20440 7236 20496
rect 7097 20438 7236 20440
rect 7097 20435 7163 20438
rect 7230 20436 7236 20438
rect 7300 20436 7306 20500
rect 11605 20362 11671 20365
rect 11240 20360 11671 20362
rect 11240 20304 11610 20360
rect 11666 20304 11671 20360
rect 11240 20302 11671 20304
rect 4419 20160 4735 20161
rect 0 20090 400 20120
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 4061 20090 4127 20093
rect 0 20088 4127 20090
rect 0 20032 4066 20088
rect 4122 20032 4127 20088
rect 0 20030 4127 20032
rect 0 20000 400 20030
rect 4061 20027 4127 20030
rect 10225 19954 10291 19957
rect 11240 19954 11300 20302
rect 11605 20299 11671 20302
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 11421 19954 11487 19957
rect 10225 19952 11487 19954
rect 10225 19896 10230 19952
rect 10286 19896 11426 19952
rect 11482 19896 11487 19952
rect 10225 19894 11487 19896
rect 10225 19891 10291 19894
rect 11421 19891 11487 19894
rect 16430 19892 16436 19956
rect 16500 19954 16506 19956
rect 18229 19954 18295 19957
rect 16500 19952 18295 19954
rect 16500 19896 18234 19952
rect 18290 19896 18295 19952
rect 16500 19894 18295 19896
rect 16500 19892 16506 19894
rect 18229 19891 18295 19894
rect 11094 19756 11100 19820
rect 11164 19818 11170 19820
rect 11237 19818 11303 19821
rect 11164 19816 11303 19818
rect 11164 19760 11242 19816
rect 11298 19760 11303 19816
rect 11164 19758 11303 19760
rect 11164 19756 11170 19758
rect 11237 19755 11303 19758
rect 6545 19684 6611 19685
rect 6494 19620 6500 19684
rect 6564 19682 6611 19684
rect 9765 19684 9831 19685
rect 9765 19682 9812 19684
rect 6564 19680 6656 19682
rect 6606 19624 6656 19680
rect 6564 19622 6656 19624
rect 9724 19680 9812 19682
rect 9876 19682 9882 19684
rect 11329 19682 11395 19685
rect 12157 19682 12223 19685
rect 9876 19680 12223 19682
rect 9724 19624 9770 19680
rect 9876 19624 11334 19680
rect 11390 19624 12162 19680
rect 12218 19624 12223 19680
rect 9724 19622 9812 19624
rect 6564 19620 6611 19622
rect 6545 19619 6611 19620
rect 9765 19620 9812 19622
rect 9876 19622 12223 19624
rect 9876 19620 9882 19622
rect 9765 19619 9831 19620
rect 11329 19619 11395 19622
rect 12157 19619 12223 19622
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 10133 19546 10199 19549
rect 11053 19546 11119 19549
rect 12341 19546 12407 19549
rect 10133 19544 12407 19546
rect 10133 19488 10138 19544
rect 10194 19488 11058 19544
rect 11114 19488 12346 19544
rect 12402 19488 12407 19544
rect 10133 19486 12407 19488
rect 10133 19483 10199 19486
rect 11053 19483 11119 19486
rect 12341 19483 12407 19486
rect 5625 19410 5691 19413
rect 6126 19410 6132 19412
rect 5625 19408 6132 19410
rect 5625 19352 5630 19408
rect 5686 19352 6132 19408
rect 5625 19350 6132 19352
rect 5625 19347 5691 19350
rect 6126 19348 6132 19350
rect 6196 19410 6202 19412
rect 6545 19410 6611 19413
rect 6196 19408 6611 19410
rect 6196 19352 6550 19408
rect 6606 19352 6611 19408
rect 6196 19350 6611 19352
rect 6196 19348 6202 19350
rect 6545 19347 6611 19350
rect 20110 19348 20116 19412
rect 20180 19410 20186 19412
rect 22185 19410 22251 19413
rect 20180 19408 22251 19410
rect 20180 19352 22190 19408
rect 22246 19352 22251 19408
rect 20180 19350 22251 19352
rect 20180 19348 20186 19350
rect 22185 19347 22251 19350
rect 23381 19412 23447 19413
rect 23381 19408 23428 19412
rect 23492 19410 23498 19412
rect 23381 19352 23386 19408
rect 23381 19348 23428 19352
rect 23492 19350 23538 19410
rect 23492 19348 23498 19350
rect 23381 19347 23447 19348
rect 9765 19274 9831 19277
rect 13721 19274 13787 19277
rect 9765 19272 13787 19274
rect 9765 19216 9770 19272
rect 9826 19216 13726 19272
rect 13782 19216 13787 19272
rect 9765 19214 13787 19216
rect 9765 19211 9831 19214
rect 13721 19211 13787 19214
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 5993 18866 6059 18869
rect 8753 18866 8819 18869
rect 5993 18864 8819 18866
rect 5993 18808 5998 18864
rect 6054 18808 8758 18864
rect 8814 18808 8819 18864
rect 5993 18806 8819 18808
rect 5993 18803 6059 18806
rect 8753 18803 8819 18806
rect 7097 18730 7163 18733
rect 7230 18730 7236 18732
rect 7097 18728 7236 18730
rect 7097 18672 7102 18728
rect 7158 18672 7236 18728
rect 7097 18670 7236 18672
rect 7097 18667 7163 18670
rect 7230 18668 7236 18670
rect 7300 18668 7306 18732
rect 8886 18532 8892 18596
rect 8956 18594 8962 18596
rect 9489 18594 9555 18597
rect 8956 18592 9555 18594
rect 8956 18536 9494 18592
rect 9550 18536 9555 18592
rect 8956 18534 9555 18536
rect 8956 18532 8962 18534
rect 9489 18531 9555 18534
rect 22185 18594 22251 18597
rect 22318 18594 22324 18596
rect 22185 18592 22324 18594
rect 22185 18536 22190 18592
rect 22246 18536 22324 18592
rect 22185 18534 22324 18536
rect 22185 18531 22251 18534
rect 22318 18532 22324 18534
rect 22388 18594 22394 18596
rect 23105 18594 23171 18597
rect 22388 18592 23171 18594
rect 22388 18536 23110 18592
rect 23166 18536 23171 18592
rect 22388 18534 23171 18536
rect 22388 18532 22394 18534
rect 23105 18531 23171 18534
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 0 18050 400 18080
rect 3877 18050 3943 18053
rect 0 18048 3943 18050
rect 0 17992 3882 18048
rect 3938 17992 3943 18048
rect 0 17990 3943 17992
rect 0 17960 400 17990
rect 3877 17987 3943 17990
rect 15694 17988 15700 18052
rect 15764 18050 15770 18052
rect 17953 18050 18019 18053
rect 15764 18048 18019 18050
rect 15764 17992 17958 18048
rect 18014 17992 18019 18048
rect 15764 17990 18019 17992
rect 15764 17988 15770 17990
rect 17953 17987 18019 17990
rect 20478 17988 20484 18052
rect 20548 18050 20554 18052
rect 24393 18050 24459 18053
rect 20548 18048 24459 18050
rect 20548 17992 24398 18048
rect 24454 17992 24459 18048
rect 20548 17990 24459 17992
rect 20548 17988 20554 17990
rect 24393 17987 24459 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 7465 17642 7531 17645
rect 7598 17642 7604 17644
rect 7465 17640 7604 17642
rect 7465 17584 7470 17640
rect 7526 17584 7604 17640
rect 7465 17582 7604 17584
rect 7465 17579 7531 17582
rect 7598 17580 7604 17582
rect 7668 17580 7674 17644
rect 9489 17642 9555 17645
rect 15285 17642 15351 17645
rect 9489 17640 15351 17642
rect 9489 17584 9494 17640
rect 9550 17584 15290 17640
rect 15346 17584 15351 17640
rect 9489 17582 15351 17584
rect 9489 17579 9555 17582
rect 15285 17579 15351 17582
rect 6269 17506 6335 17509
rect 6494 17506 6500 17508
rect 6269 17504 6500 17506
rect 6269 17448 6274 17504
rect 6330 17448 6500 17504
rect 6269 17446 6500 17448
rect 6269 17443 6335 17446
rect 6494 17444 6500 17446
rect 6564 17444 6570 17508
rect 12893 17506 12959 17509
rect 14365 17506 14431 17509
rect 12893 17504 14431 17506
rect 12893 17448 12898 17504
rect 12954 17448 14370 17504
rect 14426 17448 14431 17504
rect 12893 17446 14431 17448
rect 12893 17443 12959 17446
rect 14365 17443 14431 17446
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 9121 16826 9187 16829
rect 9581 16826 9647 16829
rect 9121 16824 9647 16826
rect 9121 16768 9126 16824
rect 9182 16768 9586 16824
rect 9642 16768 9647 16824
rect 9121 16766 9647 16768
rect 9121 16763 9187 16766
rect 9581 16763 9647 16766
rect 18781 16826 18847 16829
rect 19333 16826 19399 16829
rect 18781 16824 19399 16826
rect 18781 16768 18786 16824
rect 18842 16768 19338 16824
rect 19394 16768 19399 16824
rect 18781 16766 19399 16768
rect 18781 16763 18847 16766
rect 19333 16763 19399 16766
rect 9305 16692 9371 16693
rect 9254 16690 9260 16692
rect 9214 16630 9260 16690
rect 9324 16688 9371 16692
rect 9366 16632 9371 16688
rect 9254 16628 9260 16630
rect 9324 16628 9371 16632
rect 9305 16627 9371 16628
rect 11697 16690 11763 16693
rect 11830 16690 11836 16692
rect 11697 16688 11836 16690
rect 11697 16632 11702 16688
rect 11758 16632 11836 16688
rect 11697 16630 11836 16632
rect 11697 16627 11763 16630
rect 11830 16628 11836 16630
rect 11900 16628 11906 16692
rect 17718 16628 17724 16692
rect 17788 16690 17794 16692
rect 17861 16690 17927 16693
rect 17788 16688 17927 16690
rect 17788 16632 17866 16688
rect 17922 16632 17927 16688
rect 17788 16630 17927 16632
rect 17788 16628 17794 16630
rect 17861 16627 17927 16630
rect 20437 16690 20503 16693
rect 23197 16690 23263 16693
rect 20437 16688 23263 16690
rect 20437 16632 20442 16688
rect 20498 16632 23202 16688
rect 23258 16632 23263 16688
rect 20437 16630 23263 16632
rect 20437 16627 20503 16630
rect 23197 16627 23263 16630
rect 8937 16554 9003 16557
rect 9622 16554 9628 16556
rect 8937 16552 9628 16554
rect 8937 16496 8942 16552
rect 8998 16496 9628 16552
rect 8937 16494 9628 16496
rect 8937 16491 9003 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 16297 16554 16363 16557
rect 21265 16554 21331 16557
rect 16297 16552 21331 16554
rect 16297 16496 16302 16552
rect 16358 16496 21270 16552
rect 21326 16496 21331 16552
rect 16297 16494 21331 16496
rect 16297 16491 16363 16494
rect 21265 16491 21331 16494
rect 18137 16418 18203 16421
rect 19425 16418 19491 16421
rect 18137 16416 19491 16418
rect 18137 16360 18142 16416
rect 18198 16360 19430 16416
rect 19486 16360 19491 16416
rect 18137 16358 19491 16360
rect 18137 16355 18203 16358
rect 19425 16355 19491 16358
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 19425 16282 19491 16285
rect 19977 16282 20043 16285
rect 19425 16280 20043 16282
rect 19425 16224 19430 16280
rect 19486 16224 19982 16280
rect 20038 16224 20043 16280
rect 19425 16222 20043 16224
rect 19425 16219 19491 16222
rect 19977 16219 20043 16222
rect 23473 16282 23539 16285
rect 23749 16282 23815 16285
rect 23473 16280 23815 16282
rect 23473 16224 23478 16280
rect 23534 16224 23754 16280
rect 23810 16224 23815 16280
rect 23473 16222 23815 16224
rect 23473 16219 23539 16222
rect 23749 16219 23815 16222
rect 6269 16146 6335 16149
rect 8109 16146 8175 16149
rect 6269 16144 8175 16146
rect 6269 16088 6274 16144
rect 6330 16088 8114 16144
rect 8170 16088 8175 16144
rect 6269 16086 8175 16088
rect 6269 16083 6335 16086
rect 8109 16083 8175 16086
rect 9673 16146 9739 16149
rect 11145 16146 11211 16149
rect 9673 16144 11211 16146
rect 9673 16088 9678 16144
rect 9734 16088 11150 16144
rect 11206 16088 11211 16144
rect 9673 16086 11211 16088
rect 9673 16083 9739 16086
rect 11145 16083 11211 16086
rect 19701 16146 19767 16149
rect 22645 16146 22711 16149
rect 23473 16146 23539 16149
rect 19701 16144 23539 16146
rect 19701 16088 19706 16144
rect 19762 16088 22650 16144
rect 22706 16088 23478 16144
rect 23534 16088 23539 16144
rect 19701 16086 23539 16088
rect 19701 16083 19767 16086
rect 22645 16083 22711 16086
rect 23473 16083 23539 16086
rect 0 16010 400 16040
rect 657 16010 723 16013
rect 0 16008 723 16010
rect 0 15952 662 16008
rect 718 15952 723 16008
rect 0 15950 723 15952
rect 0 15920 400 15950
rect 657 15947 723 15950
rect 4102 15948 4108 16012
rect 4172 16010 4178 16012
rect 4521 16010 4587 16013
rect 4172 16008 4587 16010
rect 4172 15952 4526 16008
rect 4582 15952 4587 16008
rect 4172 15950 4587 15952
rect 4172 15948 4178 15950
rect 4521 15947 4587 15950
rect 6126 15948 6132 16012
rect 6196 16010 6202 16012
rect 6913 16010 6979 16013
rect 6196 16008 6979 16010
rect 6196 15952 6918 16008
rect 6974 15952 6979 16008
rect 6196 15950 6979 15952
rect 6196 15948 6202 15950
rect 6913 15947 6979 15950
rect 18781 16010 18847 16013
rect 21265 16010 21331 16013
rect 18781 16008 21331 16010
rect 18781 15952 18786 16008
rect 18842 15952 21270 16008
rect 21326 15952 21331 16008
rect 18781 15950 21331 15952
rect 18781 15947 18847 15950
rect 21265 15947 21331 15950
rect 19149 15874 19215 15877
rect 20253 15874 20319 15877
rect 19149 15872 20319 15874
rect 19149 15816 19154 15872
rect 19210 15816 20258 15872
rect 20314 15816 20319 15872
rect 19149 15814 20319 15816
rect 19149 15811 19215 15814
rect 20253 15811 20319 15814
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 19241 15738 19307 15741
rect 22737 15738 22803 15741
rect 19241 15736 22803 15738
rect 19241 15680 19246 15736
rect 19302 15680 22742 15736
rect 22798 15680 22803 15736
rect 19241 15678 22803 15680
rect 19241 15675 19307 15678
rect 22737 15675 22803 15678
rect 3049 15602 3115 15605
rect 6085 15602 6151 15605
rect 9397 15604 9463 15605
rect 3049 15600 6151 15602
rect 3049 15544 3054 15600
rect 3110 15544 6090 15600
rect 6146 15544 6151 15600
rect 3049 15542 6151 15544
rect 3049 15539 3115 15542
rect 6085 15539 6151 15542
rect 7414 15540 7420 15604
rect 7484 15602 7490 15604
rect 9397 15602 9444 15604
rect 7484 15600 9444 15602
rect 9508 15602 9514 15604
rect 10869 15602 10935 15605
rect 18086 15602 18092 15604
rect 7484 15544 9402 15600
rect 7484 15542 9444 15544
rect 7484 15540 7490 15542
rect 9397 15540 9444 15542
rect 9508 15542 9590 15602
rect 10869 15600 18092 15602
rect 10869 15544 10874 15600
rect 10930 15544 18092 15600
rect 10869 15542 18092 15544
rect 9508 15540 9514 15542
rect 9397 15539 9463 15540
rect 10869 15539 10935 15542
rect 18086 15540 18092 15542
rect 18156 15540 18162 15604
rect 21398 15540 21404 15604
rect 21468 15602 21474 15604
rect 21909 15602 21975 15605
rect 21468 15600 21975 15602
rect 21468 15544 21914 15600
rect 21970 15544 21975 15600
rect 21468 15542 21975 15544
rect 21468 15540 21474 15542
rect 21909 15539 21975 15542
rect 8385 15466 8451 15469
rect 9305 15466 9371 15469
rect 8385 15464 9371 15466
rect 8385 15408 8390 15464
rect 8446 15408 9310 15464
rect 9366 15408 9371 15464
rect 8385 15406 9371 15408
rect 8385 15403 8451 15406
rect 9305 15403 9371 15406
rect 14590 15404 14596 15468
rect 14660 15466 14666 15468
rect 20713 15466 20779 15469
rect 14660 15464 20779 15466
rect 14660 15408 20718 15464
rect 20774 15408 20779 15464
rect 14660 15406 20779 15408
rect 14660 15404 14666 15406
rect 20713 15403 20779 15406
rect 21725 15466 21791 15469
rect 24117 15466 24183 15469
rect 21725 15464 24183 15466
rect 21725 15408 21730 15464
rect 21786 15408 24122 15464
rect 24178 15408 24183 15464
rect 21725 15406 24183 15408
rect 21725 15403 21791 15406
rect 24117 15403 24183 15406
rect 11605 15330 11671 15333
rect 13854 15330 13860 15332
rect 11605 15328 13860 15330
rect 11605 15272 11610 15328
rect 11666 15272 13860 15328
rect 11605 15270 13860 15272
rect 11605 15267 11671 15270
rect 13854 15268 13860 15270
rect 13924 15268 13930 15332
rect 17902 15268 17908 15332
rect 17972 15330 17978 15332
rect 18321 15330 18387 15333
rect 17972 15328 18387 15330
rect 17972 15272 18326 15328
rect 18382 15272 18387 15328
rect 17972 15270 18387 15272
rect 17972 15268 17978 15270
rect 18321 15267 18387 15270
rect 22502 15268 22508 15332
rect 22572 15330 22578 15332
rect 22829 15330 22895 15333
rect 22572 15328 22895 15330
rect 22572 15272 22834 15328
rect 22890 15272 22895 15328
rect 22572 15270 22895 15272
rect 22572 15268 22578 15270
rect 22829 15267 22895 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 8937 15194 9003 15197
rect 8710 15192 9003 15194
rect 8710 15136 8942 15192
rect 8998 15136 9003 15192
rect 8710 15134 9003 15136
rect 3366 14996 3372 15060
rect 3436 15058 3442 15060
rect 8710 15058 8770 15134
rect 8937 15131 9003 15134
rect 3436 14998 8770 15058
rect 3436 14996 3442 14998
rect 19926 14996 19932 15060
rect 19996 15058 20002 15060
rect 20069 15058 20135 15061
rect 19996 15056 20135 15058
rect 19996 15000 20074 15056
rect 20130 15000 20135 15056
rect 19996 14998 20135 15000
rect 19996 14996 20002 14998
rect 20069 14995 20135 14998
rect 7230 14860 7236 14924
rect 7300 14922 7306 14924
rect 9581 14922 9647 14925
rect 7300 14920 9647 14922
rect 7300 14864 9586 14920
rect 9642 14864 9647 14920
rect 7300 14862 9647 14864
rect 7300 14860 7306 14862
rect 9581 14859 9647 14862
rect 8017 14786 8083 14789
rect 9305 14786 9371 14789
rect 9581 14786 9647 14789
rect 8017 14784 9647 14786
rect 8017 14728 8022 14784
rect 8078 14728 9310 14784
rect 9366 14728 9586 14784
rect 9642 14728 9647 14784
rect 8017 14726 9647 14728
rect 8017 14723 8083 14726
rect 9305 14723 9371 14726
rect 9581 14723 9647 14726
rect 21030 14724 21036 14788
rect 21100 14786 21106 14788
rect 21173 14786 21239 14789
rect 21100 14784 21239 14786
rect 21100 14728 21178 14784
rect 21234 14728 21239 14784
rect 21100 14726 21239 14728
rect 21100 14724 21106 14726
rect 21173 14723 21239 14726
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 10225 14514 10291 14517
rect 11789 14514 11855 14517
rect 10225 14512 11855 14514
rect 10225 14456 10230 14512
rect 10286 14456 11794 14512
rect 11850 14456 11855 14512
rect 10225 14454 11855 14456
rect 10225 14451 10291 14454
rect 11789 14451 11855 14454
rect 9121 14378 9187 14381
rect 9489 14378 9555 14381
rect 9121 14376 9555 14378
rect 9121 14320 9126 14376
rect 9182 14320 9494 14376
rect 9550 14320 9555 14376
rect 9121 14318 9555 14320
rect 9121 14315 9187 14318
rect 9489 14315 9555 14318
rect 8886 14180 8892 14244
rect 8956 14242 8962 14244
rect 12709 14242 12775 14245
rect 8956 14240 12775 14242
rect 8956 14184 12714 14240
rect 12770 14184 12775 14240
rect 8956 14182 12775 14184
rect 8956 14180 8962 14182
rect 12709 14179 12775 14182
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 0 13970 400 14000
rect 565 13970 631 13973
rect 0 13968 631 13970
rect 0 13912 570 13968
rect 626 13912 631 13968
rect 0 13910 631 13912
rect 0 13880 400 13910
rect 565 13907 631 13910
rect 16665 13970 16731 13973
rect 18689 13970 18755 13973
rect 16665 13968 18755 13970
rect 16665 13912 16670 13968
rect 16726 13912 18694 13968
rect 18750 13912 18755 13968
rect 16665 13910 18755 13912
rect 16665 13907 16731 13910
rect 18689 13907 18755 13910
rect 20253 13970 20319 13973
rect 21030 13970 21036 13972
rect 20253 13968 21036 13970
rect 20253 13912 20258 13968
rect 20314 13912 21036 13968
rect 20253 13910 21036 13912
rect 20253 13907 20319 13910
rect 21030 13908 21036 13910
rect 21100 13908 21106 13972
rect 8293 13834 8359 13837
rect 9622 13834 9628 13836
rect 8293 13832 9628 13834
rect 8293 13776 8298 13832
rect 8354 13776 9628 13832
rect 8293 13774 9628 13776
rect 8293 13771 8359 13774
rect 9622 13772 9628 13774
rect 9692 13772 9698 13836
rect 15469 13834 15535 13837
rect 17309 13834 17375 13837
rect 18321 13834 18387 13837
rect 15469 13832 18387 13834
rect 15469 13776 15474 13832
rect 15530 13776 17314 13832
rect 17370 13776 18326 13832
rect 18382 13776 18387 13832
rect 15469 13774 18387 13776
rect 15469 13771 15535 13774
rect 17309 13771 17375 13774
rect 18321 13771 18387 13774
rect 11830 13636 11836 13700
rect 11900 13698 11906 13700
rect 17350 13698 17356 13700
rect 11900 13638 17356 13698
rect 11900 13636 11906 13638
rect 17350 13636 17356 13638
rect 17420 13636 17426 13700
rect 22185 13698 22251 13701
rect 22318 13698 22324 13700
rect 22185 13696 22324 13698
rect 22185 13640 22190 13696
rect 22246 13640 22324 13696
rect 22185 13638 22324 13640
rect 22185 13635 22251 13638
rect 22318 13636 22324 13638
rect 22388 13636 22394 13700
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 14457 13562 14523 13565
rect 15377 13562 15443 13565
rect 14457 13560 15443 13562
rect 14457 13504 14462 13560
rect 14518 13504 15382 13560
rect 15438 13504 15443 13560
rect 14457 13502 15443 13504
rect 14457 13499 14523 13502
rect 15377 13499 15443 13502
rect 15653 13562 15719 13565
rect 16389 13562 16455 13565
rect 15653 13560 16455 13562
rect 15653 13504 15658 13560
rect 15714 13504 16394 13560
rect 16450 13504 16455 13560
rect 15653 13502 16455 13504
rect 15653 13499 15719 13502
rect 16389 13499 16455 13502
rect 12433 13426 12499 13429
rect 16113 13426 16179 13429
rect 12433 13424 16179 13426
rect 12433 13368 12438 13424
rect 12494 13368 16118 13424
rect 16174 13368 16179 13424
rect 12433 13366 16179 13368
rect 12433 13363 12499 13366
rect 16113 13363 16179 13366
rect 9673 13290 9739 13293
rect 9630 13288 9739 13290
rect 9630 13232 9678 13288
rect 9734 13232 9739 13288
rect 9630 13227 9739 13232
rect 15929 13290 15995 13293
rect 19701 13290 19767 13293
rect 20253 13292 20319 13293
rect 20253 13290 20300 13292
rect 15929 13288 19767 13290
rect 15929 13232 15934 13288
rect 15990 13232 19706 13288
rect 19762 13232 19767 13288
rect 15929 13230 19767 13232
rect 20208 13288 20300 13290
rect 20208 13232 20258 13288
rect 20208 13230 20300 13232
rect 15929 13227 15995 13230
rect 19701 13227 19767 13230
rect 20253 13228 20300 13230
rect 20364 13228 20370 13292
rect 20253 13227 20319 13228
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 9630 13021 9690 13227
rect 16941 13154 17007 13157
rect 18781 13154 18847 13157
rect 16941 13152 18847 13154
rect 16941 13096 16946 13152
rect 17002 13096 18786 13152
rect 18842 13096 18847 13152
rect 16941 13094 18847 13096
rect 16941 13091 17007 13094
rect 18781 13091 18847 13094
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 9630 13016 9739 13021
rect 9630 12960 9678 13016
rect 9734 12960 9739 13016
rect 9630 12958 9739 12960
rect 9673 12955 9739 12958
rect 16982 12956 16988 13020
rect 17052 13018 17058 13020
rect 17493 13018 17559 13021
rect 17052 13016 17559 13018
rect 17052 12960 17498 13016
rect 17554 12960 17559 13016
rect 17052 12958 17559 12960
rect 17052 12956 17058 12958
rect 17493 12955 17559 12958
rect 9438 12820 9444 12884
rect 9508 12882 9514 12884
rect 9581 12882 9647 12885
rect 9508 12880 9647 12882
rect 9508 12824 9586 12880
rect 9642 12824 9647 12880
rect 9508 12822 9647 12824
rect 9508 12820 9514 12822
rect 9581 12819 9647 12822
rect 15653 12882 15719 12885
rect 22502 12882 22508 12884
rect 15653 12880 22508 12882
rect 15653 12824 15658 12880
rect 15714 12824 22508 12880
rect 15653 12822 22508 12824
rect 15653 12819 15719 12822
rect 22502 12820 22508 12822
rect 22572 12820 22578 12884
rect 17769 12746 17835 12749
rect 18045 12746 18111 12749
rect 17769 12744 18111 12746
rect 17769 12688 17774 12744
rect 17830 12688 18050 12744
rect 18106 12688 18111 12744
rect 17769 12686 18111 12688
rect 17769 12683 17835 12686
rect 18045 12683 18111 12686
rect 19885 12746 19951 12749
rect 22829 12746 22895 12749
rect 19885 12744 22895 12746
rect 19885 12688 19890 12744
rect 19946 12688 22834 12744
rect 22890 12688 22895 12744
rect 19885 12686 22895 12688
rect 19885 12683 19951 12686
rect 22829 12683 22895 12686
rect 13813 12610 13879 12613
rect 17953 12610 18019 12613
rect 13813 12608 18019 12610
rect 13813 12552 13818 12608
rect 13874 12552 17958 12608
rect 18014 12552 18019 12608
rect 13813 12550 18019 12552
rect 13813 12547 13879 12550
rect 17953 12547 18019 12550
rect 25814 12548 25820 12612
rect 25884 12610 25890 12612
rect 26141 12610 26207 12613
rect 25884 12608 26207 12610
rect 25884 12552 26146 12608
rect 26202 12552 26207 12608
rect 25884 12550 26207 12552
rect 25884 12548 25890 12550
rect 26141 12547 26207 12550
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 18137 12340 18203 12341
rect 18086 12276 18092 12340
rect 18156 12338 18203 12340
rect 19517 12338 19583 12341
rect 19977 12338 20043 12341
rect 18156 12336 18248 12338
rect 18198 12280 18248 12336
rect 18156 12278 18248 12280
rect 19517 12336 20043 12338
rect 19517 12280 19522 12336
rect 19578 12280 19982 12336
rect 20038 12280 20043 12336
rect 19517 12278 20043 12280
rect 18156 12276 18203 12278
rect 18137 12275 18203 12276
rect 19517 12275 19583 12278
rect 19977 12275 20043 12278
rect 20253 12338 20319 12341
rect 20253 12336 22570 12338
rect 20253 12280 20258 12336
rect 20314 12280 22570 12336
rect 20253 12278 22570 12280
rect 20253 12275 20319 12278
rect 5073 12202 5139 12205
rect 5257 12202 5323 12205
rect 9213 12202 9279 12205
rect 5073 12200 9279 12202
rect 5073 12144 5078 12200
rect 5134 12144 5262 12200
rect 5318 12144 9218 12200
rect 9274 12144 9279 12200
rect 5073 12142 9279 12144
rect 5073 12139 5139 12142
rect 5257 12139 5323 12142
rect 9213 12139 9279 12142
rect 12801 12202 12867 12205
rect 13261 12202 13327 12205
rect 21173 12202 21239 12205
rect 12801 12200 21239 12202
rect 12801 12144 12806 12200
rect 12862 12144 13266 12200
rect 13322 12144 21178 12200
rect 21234 12144 21239 12200
rect 12801 12142 21239 12144
rect 22510 12202 22570 12278
rect 26509 12202 26575 12205
rect 22510 12200 26575 12202
rect 22510 12144 26514 12200
rect 26570 12144 26575 12200
rect 22510 12142 26575 12144
rect 12801 12139 12867 12142
rect 13261 12139 13327 12142
rect 21173 12139 21239 12142
rect 26509 12139 26575 12142
rect 22737 12066 22803 12069
rect 25037 12066 25103 12069
rect 22737 12064 25103 12066
rect 22737 12008 22742 12064
rect 22798 12008 25042 12064
rect 25098 12008 25103 12064
rect 22737 12006 25103 12008
rect 22737 12003 22803 12006
rect 25037 12003 25103 12006
rect 7892 12000 8208 12001
rect 0 11930 400 11960
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 749 11930 815 11933
rect 0 11928 815 11930
rect 0 11872 754 11928
rect 810 11872 815 11928
rect 0 11870 815 11872
rect 0 11840 400 11870
rect 749 11867 815 11870
rect 23422 11868 23428 11932
rect 23492 11930 23498 11932
rect 25037 11930 25103 11933
rect 23492 11928 25103 11930
rect 23492 11872 25042 11928
rect 25098 11872 25103 11928
rect 23492 11870 25103 11872
rect 23492 11868 23498 11870
rect 25037 11867 25103 11870
rect 13854 11732 13860 11796
rect 13924 11794 13930 11796
rect 15009 11794 15075 11797
rect 13924 11792 15075 11794
rect 13924 11736 15014 11792
rect 15070 11736 15075 11792
rect 13924 11734 15075 11736
rect 13924 11732 13930 11734
rect 15009 11731 15075 11734
rect 15929 11794 15995 11797
rect 17718 11794 17724 11796
rect 15929 11792 17724 11794
rect 15929 11736 15934 11792
rect 15990 11736 17724 11792
rect 15929 11734 17724 11736
rect 15929 11731 15995 11734
rect 17718 11732 17724 11734
rect 17788 11794 17794 11796
rect 17861 11794 17927 11797
rect 17788 11792 17927 11794
rect 17788 11736 17866 11792
rect 17922 11736 17927 11792
rect 17788 11734 17927 11736
rect 17788 11732 17794 11734
rect 17861 11731 17927 11734
rect 24301 11794 24367 11797
rect 26417 11794 26483 11797
rect 27521 11794 27587 11797
rect 24301 11792 27587 11794
rect 24301 11736 24306 11792
rect 24362 11736 26422 11792
rect 26478 11736 27526 11792
rect 27582 11736 27587 11792
rect 24301 11734 27587 11736
rect 24301 11731 24367 11734
rect 26417 11731 26483 11734
rect 27521 11731 27587 11734
rect 14089 11658 14155 11661
rect 15285 11658 15351 11661
rect 14089 11656 15351 11658
rect 14089 11600 14094 11656
rect 14150 11600 15290 11656
rect 15346 11600 15351 11656
rect 14089 11598 15351 11600
rect 14089 11595 14155 11598
rect 15285 11595 15351 11598
rect 21449 11522 21515 11525
rect 24761 11522 24827 11525
rect 21449 11520 24827 11522
rect 21449 11464 21454 11520
rect 21510 11464 24766 11520
rect 24822 11464 24827 11520
rect 21449 11462 24827 11464
rect 21449 11459 21515 11462
rect 24761 11459 24827 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 20621 11386 20687 11389
rect 21449 11386 21515 11389
rect 24301 11386 24367 11389
rect 20621 11384 24367 11386
rect 20621 11328 20626 11384
rect 20682 11328 21454 11384
rect 21510 11328 24306 11384
rect 24362 11328 24367 11384
rect 20621 11326 24367 11328
rect 20621 11323 20687 11326
rect 21449 11323 21515 11326
rect 24301 11323 24367 11326
rect 16481 11250 16547 11253
rect 19885 11250 19951 11253
rect 16481 11248 19951 11250
rect 16481 11192 16486 11248
rect 16542 11192 19890 11248
rect 19946 11192 19951 11248
rect 16481 11190 19951 11192
rect 16481 11187 16547 11190
rect 19885 11187 19951 11190
rect 23105 11250 23171 11253
rect 24393 11250 24459 11253
rect 23105 11248 24459 11250
rect 23105 11192 23110 11248
rect 23166 11192 24398 11248
rect 24454 11192 24459 11248
rect 23105 11190 24459 11192
rect 23105 11187 23171 11190
rect 24393 11187 24459 11190
rect 5257 11114 5323 11117
rect 6637 11114 6703 11117
rect 5257 11112 6703 11114
rect 5257 11056 5262 11112
rect 5318 11056 6642 11112
rect 6698 11056 6703 11112
rect 5257 11054 6703 11056
rect 5257 11051 5323 11054
rect 6637 11051 6703 11054
rect 7414 11052 7420 11116
rect 7484 11114 7490 11116
rect 8201 11114 8267 11117
rect 7484 11112 8267 11114
rect 7484 11056 8206 11112
rect 8262 11056 8267 11112
rect 7484 11054 8267 11056
rect 7484 11052 7490 11054
rect 8201 11051 8267 11054
rect 9622 11052 9628 11116
rect 9692 11114 9698 11116
rect 9692 11054 16498 11114
rect 9692 11052 9698 11054
rect 16438 10978 16498 11054
rect 16614 11052 16620 11116
rect 16684 11114 16690 11116
rect 16849 11114 16915 11117
rect 23289 11114 23355 11117
rect 16684 11112 23355 11114
rect 16684 11056 16854 11112
rect 16910 11056 23294 11112
rect 23350 11056 23355 11112
rect 16684 11054 23355 11056
rect 16684 11052 16690 11054
rect 16849 11051 16915 11054
rect 23289 11051 23355 11054
rect 18137 10978 18203 10981
rect 16438 10976 18203 10978
rect 16438 10920 18142 10976
rect 18198 10920 18203 10976
rect 16438 10918 18203 10920
rect 18137 10915 18203 10918
rect 20989 10980 21055 10981
rect 20989 10976 21036 10980
rect 21100 10978 21106 10980
rect 20989 10920 20994 10976
rect 20989 10916 21036 10920
rect 21100 10918 21146 10978
rect 21100 10916 21106 10918
rect 20989 10915 21055 10916
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 22185 10842 22251 10845
rect 23381 10842 23447 10845
rect 22185 10840 23447 10842
rect 22185 10784 22190 10840
rect 22246 10784 23386 10840
rect 23442 10784 23447 10840
rect 22185 10782 23447 10784
rect 22185 10779 22251 10782
rect 23381 10779 23447 10782
rect 19885 10706 19951 10709
rect 22369 10706 22435 10709
rect 19885 10704 22435 10706
rect 19885 10648 19890 10704
rect 19946 10648 22374 10704
rect 22430 10648 22435 10704
rect 19885 10646 22435 10648
rect 19885 10643 19951 10646
rect 22369 10643 22435 10646
rect 22829 10706 22895 10709
rect 27521 10706 27587 10709
rect 22829 10704 27587 10706
rect 22829 10648 22834 10704
rect 22890 10648 27526 10704
rect 27582 10648 27587 10704
rect 22829 10646 27587 10648
rect 22829 10643 22895 10646
rect 27521 10643 27587 10646
rect 13721 10570 13787 10573
rect 20621 10570 20687 10573
rect 13721 10568 20687 10570
rect 13721 10512 13726 10568
rect 13782 10512 20626 10568
rect 20682 10512 20687 10568
rect 13721 10510 20687 10512
rect 13721 10507 13787 10510
rect 20621 10507 20687 10510
rect 22093 10570 22159 10573
rect 22461 10570 22527 10573
rect 25221 10570 25287 10573
rect 22093 10568 25287 10570
rect 22093 10512 22098 10568
rect 22154 10512 22466 10568
rect 22522 10512 25226 10568
rect 25282 10512 25287 10568
rect 22093 10510 25287 10512
rect 22093 10507 22159 10510
rect 22461 10507 22527 10510
rect 25221 10507 25287 10510
rect 13997 10434 14063 10437
rect 16665 10434 16731 10437
rect 13997 10432 16731 10434
rect 13997 10376 14002 10432
rect 14058 10376 16670 10432
rect 16726 10376 16731 10432
rect 13997 10374 16731 10376
rect 13997 10371 14063 10374
rect 16665 10371 16731 10374
rect 18689 10434 18755 10437
rect 19885 10434 19951 10437
rect 18689 10432 19951 10434
rect 18689 10376 18694 10432
rect 18750 10376 19890 10432
rect 19946 10376 19951 10432
rect 18689 10374 19951 10376
rect 18689 10371 18755 10374
rect 19885 10371 19951 10374
rect 21081 10434 21147 10437
rect 23197 10434 23263 10437
rect 21081 10432 23263 10434
rect 21081 10376 21086 10432
rect 21142 10376 23202 10432
rect 23258 10376 23263 10432
rect 21081 10374 23263 10376
rect 21081 10371 21147 10374
rect 23197 10371 23263 10374
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 19609 10298 19675 10301
rect 21725 10298 21791 10301
rect 19609 10296 21791 10298
rect 19609 10240 19614 10296
rect 19670 10240 21730 10296
rect 21786 10240 21791 10296
rect 19609 10238 21791 10240
rect 19609 10235 19675 10238
rect 21725 10235 21791 10238
rect 19333 10162 19399 10165
rect 19609 10162 19675 10165
rect 19333 10160 19675 10162
rect 19333 10104 19338 10160
rect 19394 10104 19614 10160
rect 19670 10104 19675 10160
rect 19333 10102 19675 10104
rect 19333 10099 19399 10102
rect 19609 10099 19675 10102
rect 21357 10162 21423 10165
rect 24485 10162 24551 10165
rect 21357 10160 24551 10162
rect 21357 10104 21362 10160
rect 21418 10104 24490 10160
rect 24546 10104 24551 10160
rect 21357 10102 24551 10104
rect 21357 10099 21423 10102
rect 24485 10099 24551 10102
rect 24761 10162 24827 10165
rect 26233 10162 26299 10165
rect 24761 10160 26299 10162
rect 24761 10104 24766 10160
rect 24822 10104 26238 10160
rect 26294 10104 26299 10160
rect 24761 10102 26299 10104
rect 24761 10099 24827 10102
rect 26233 10099 26299 10102
rect 16665 10026 16731 10029
rect 22645 10026 22711 10029
rect 16665 10024 22711 10026
rect 16665 9968 16670 10024
rect 16726 9968 22650 10024
rect 22706 9968 22711 10024
rect 16665 9966 22711 9968
rect 16665 9963 16731 9966
rect 22645 9963 22711 9966
rect 0 9890 400 9920
rect 841 9890 907 9893
rect 0 9888 907 9890
rect 0 9832 846 9888
rect 902 9832 907 9888
rect 0 9830 907 9832
rect 0 9800 400 9830
rect 841 9827 907 9830
rect 19517 9890 19583 9893
rect 19517 9888 20178 9890
rect 19517 9832 19522 9888
rect 19578 9832 20178 9888
rect 19517 9830 20178 9832
rect 19517 9827 19583 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 6177 9754 6243 9757
rect 7230 9754 7236 9756
rect 6177 9752 7236 9754
rect 6177 9696 6182 9752
rect 6238 9696 7236 9752
rect 6177 9694 7236 9696
rect 6177 9691 6243 9694
rect 7230 9692 7236 9694
rect 7300 9692 7306 9756
rect 19333 9754 19399 9757
rect 19885 9754 19951 9757
rect 19333 9752 19951 9754
rect 19333 9696 19338 9752
rect 19394 9696 19890 9752
rect 19946 9696 19951 9752
rect 19333 9694 19951 9696
rect 20118 9754 20178 9830
rect 20294 9828 20300 9892
rect 20364 9890 20370 9892
rect 20989 9890 21055 9893
rect 20364 9888 21055 9890
rect 20364 9832 20994 9888
rect 21050 9832 21055 9888
rect 20364 9830 21055 9832
rect 20364 9828 20370 9830
rect 20989 9827 21055 9830
rect 22461 9890 22527 9893
rect 25497 9890 25563 9893
rect 22461 9888 25563 9890
rect 22461 9832 22466 9888
rect 22522 9832 25502 9888
rect 25558 9832 25563 9888
rect 22461 9830 25563 9832
rect 22461 9827 22527 9830
rect 25497 9827 25563 9830
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 21357 9754 21423 9757
rect 20118 9752 21423 9754
rect 20118 9696 21362 9752
rect 21418 9696 21423 9752
rect 20118 9694 21423 9696
rect 19333 9691 19399 9694
rect 19885 9691 19951 9694
rect 21357 9691 21423 9694
rect 22553 9754 22619 9757
rect 24117 9754 24183 9757
rect 22553 9752 24183 9754
rect 22553 9696 22558 9752
rect 22614 9696 24122 9752
rect 24178 9696 24183 9752
rect 22553 9694 24183 9696
rect 22553 9691 22619 9694
rect 24117 9691 24183 9694
rect 19517 9618 19583 9621
rect 19885 9620 19951 9621
rect 19742 9618 19748 9620
rect 19517 9616 19748 9618
rect 19517 9560 19522 9616
rect 19578 9560 19748 9616
rect 19517 9558 19748 9560
rect 19517 9555 19583 9558
rect 19742 9556 19748 9558
rect 19812 9556 19818 9620
rect 19885 9616 19932 9620
rect 19996 9618 20002 9620
rect 19885 9560 19890 9616
rect 19885 9556 19932 9560
rect 19996 9558 20042 9618
rect 19996 9556 20002 9558
rect 20294 9556 20300 9620
rect 20364 9618 20370 9620
rect 20621 9618 20687 9621
rect 20364 9616 20687 9618
rect 20364 9560 20626 9616
rect 20682 9560 20687 9616
rect 20364 9558 20687 9560
rect 20364 9556 20370 9558
rect 19885 9555 19951 9556
rect 20621 9555 20687 9558
rect 22737 9618 22803 9621
rect 27705 9618 27771 9621
rect 22737 9616 27771 9618
rect 22737 9560 22742 9616
rect 22798 9560 27710 9616
rect 27766 9560 27771 9616
rect 22737 9558 27771 9560
rect 22737 9555 22803 9558
rect 27705 9555 27771 9558
rect 18137 9482 18203 9485
rect 20478 9482 20484 9484
rect 18137 9480 20484 9482
rect 18137 9424 18142 9480
rect 18198 9424 20484 9480
rect 18137 9422 20484 9424
rect 18137 9419 18203 9422
rect 20478 9420 20484 9422
rect 20548 9420 20554 9484
rect 25405 9482 25471 9485
rect 26693 9482 26759 9485
rect 25405 9480 26759 9482
rect 25405 9424 25410 9480
rect 25466 9424 26698 9480
rect 26754 9424 26759 9480
rect 25405 9422 26759 9424
rect 25405 9419 25471 9422
rect 26693 9419 26759 9422
rect 19609 9346 19675 9349
rect 23422 9346 23428 9348
rect 19609 9344 23428 9346
rect 19609 9288 19614 9344
rect 19670 9288 23428 9344
rect 19609 9286 23428 9288
rect 19609 9283 19675 9286
rect 23422 9284 23428 9286
rect 23492 9284 23498 9348
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 13629 9210 13695 9213
rect 17953 9210 18019 9213
rect 13629 9208 18019 9210
rect 13629 9152 13634 9208
rect 13690 9152 17958 9208
rect 18014 9152 18019 9208
rect 13629 9150 18019 9152
rect 13629 9147 13695 9150
rect 17953 9147 18019 9150
rect 19742 9148 19748 9212
rect 19812 9210 19818 9212
rect 19812 9150 20178 9210
rect 19812 9148 19818 9150
rect 15653 9076 15719 9077
rect 15653 9072 15700 9076
rect 15764 9074 15770 9076
rect 15653 9016 15658 9072
rect 15653 9012 15700 9016
rect 15764 9014 15810 9074
rect 15764 9012 15770 9014
rect 16430 9012 16436 9076
rect 16500 9074 16506 9076
rect 16941 9074 17007 9077
rect 16500 9072 17007 9074
rect 16500 9016 16946 9072
rect 17002 9016 17007 9072
rect 16500 9014 17007 9016
rect 16500 9012 16506 9014
rect 15653 9011 15719 9012
rect 16941 9011 17007 9014
rect 17350 9012 17356 9076
rect 17420 9074 17426 9076
rect 18321 9074 18387 9077
rect 17420 9072 18387 9074
rect 17420 9016 18326 9072
rect 18382 9016 18387 9072
rect 17420 9014 18387 9016
rect 20118 9074 20178 9150
rect 24025 9074 24091 9077
rect 20118 9072 24091 9074
rect 20118 9016 24030 9072
rect 24086 9016 24091 9072
rect 20118 9014 24091 9016
rect 17420 9012 17426 9014
rect 18321 9011 18387 9014
rect 24025 9011 24091 9014
rect 12525 8938 12591 8941
rect 15285 8938 15351 8941
rect 12525 8936 15351 8938
rect 12525 8880 12530 8936
rect 12586 8880 15290 8936
rect 15346 8880 15351 8936
rect 12525 8878 15351 8880
rect 12525 8875 12591 8878
rect 15285 8875 15351 8878
rect 20621 8938 20687 8941
rect 23933 8938 23999 8941
rect 20621 8936 23999 8938
rect 20621 8880 20626 8936
rect 20682 8880 23938 8936
rect 23994 8880 23999 8936
rect 20621 8878 23999 8880
rect 20621 8875 20687 8878
rect 23933 8875 23999 8878
rect 18045 8802 18111 8805
rect 19701 8802 19767 8805
rect 18045 8800 19767 8802
rect 18045 8744 18050 8800
rect 18106 8744 19706 8800
rect 19762 8744 19767 8800
rect 18045 8742 19767 8744
rect 18045 8739 18111 8742
rect 19701 8739 19767 8742
rect 24393 8802 24459 8805
rect 25313 8802 25379 8805
rect 25814 8802 25820 8804
rect 24393 8800 25820 8802
rect 24393 8744 24398 8800
rect 24454 8744 25318 8800
rect 25374 8744 25820 8800
rect 24393 8742 25820 8744
rect 24393 8739 24459 8742
rect 25313 8739 25379 8742
rect 25814 8740 25820 8742
rect 25884 8740 25890 8804
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 19333 8666 19399 8669
rect 20621 8666 20687 8669
rect 19333 8664 20687 8666
rect 19333 8608 19338 8664
rect 19394 8608 20626 8664
rect 20682 8608 20687 8664
rect 19333 8606 20687 8608
rect 19333 8603 19399 8606
rect 17953 8530 18019 8533
rect 18321 8530 18387 8533
rect 17953 8528 18387 8530
rect 17953 8472 17958 8528
rect 18014 8472 18326 8528
rect 18382 8472 18387 8528
rect 17953 8470 18387 8472
rect 17953 8467 18019 8470
rect 18321 8467 18387 8470
rect 19566 8397 19626 8606
rect 20621 8603 20687 8606
rect 13670 8332 13676 8396
rect 13740 8394 13746 8396
rect 16982 8394 16988 8396
rect 13740 8334 16988 8394
rect 13740 8332 13746 8334
rect 16982 8332 16988 8334
rect 17052 8332 17058 8396
rect 18045 8394 18111 8397
rect 18873 8394 18939 8397
rect 18045 8392 18939 8394
rect 18045 8336 18050 8392
rect 18106 8336 18878 8392
rect 18934 8336 18939 8392
rect 18045 8334 18939 8336
rect 19566 8392 19675 8397
rect 19566 8336 19614 8392
rect 19670 8336 19675 8392
rect 19566 8334 19675 8336
rect 18045 8331 18111 8334
rect 18873 8331 18939 8334
rect 19609 8331 19675 8334
rect 14273 8258 14339 8261
rect 17902 8258 17908 8260
rect 14273 8256 17908 8258
rect 14273 8200 14278 8256
rect 14334 8200 17908 8256
rect 14273 8198 17908 8200
rect 14273 8195 14339 8198
rect 17902 8196 17908 8198
rect 17972 8196 17978 8260
rect 19425 8258 19491 8261
rect 22277 8258 22343 8261
rect 19425 8256 22343 8258
rect 19425 8200 19430 8256
rect 19486 8200 22282 8256
rect 22338 8200 22343 8256
rect 19425 8198 22343 8200
rect 19425 8195 19491 8198
rect 22277 8195 22343 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 19425 8122 19491 8125
rect 20294 8122 20300 8124
rect 19425 8120 20300 8122
rect 19425 8064 19430 8120
rect 19486 8064 20300 8120
rect 19425 8062 20300 8064
rect 19425 8059 19491 8062
rect 20294 8060 20300 8062
rect 20364 8060 20370 8124
rect 22277 7986 22343 7989
rect 22737 7986 22803 7989
rect 22277 7984 22803 7986
rect 22277 7928 22282 7984
rect 22338 7928 22742 7984
rect 22798 7928 22803 7984
rect 22277 7926 22803 7928
rect 22277 7923 22343 7926
rect 22737 7923 22803 7926
rect 0 7850 400 7880
rect 933 7850 999 7853
rect 0 7848 999 7850
rect 0 7792 938 7848
rect 994 7792 999 7848
rect 0 7790 999 7792
rect 0 7760 400 7790
rect 933 7787 999 7790
rect 3550 7788 3556 7852
rect 3620 7850 3626 7852
rect 13118 7850 13124 7852
rect 3620 7790 13124 7850
rect 3620 7788 3626 7790
rect 13118 7788 13124 7790
rect 13188 7788 13194 7852
rect 21817 7850 21883 7853
rect 23381 7850 23447 7853
rect 21817 7848 23447 7850
rect 21817 7792 21822 7848
rect 21878 7792 23386 7848
rect 23442 7792 23447 7848
rect 21817 7790 23447 7792
rect 21817 7787 21883 7790
rect 23381 7787 23447 7790
rect 11881 7714 11947 7717
rect 12433 7714 12499 7717
rect 11881 7712 12499 7714
rect 11881 7656 11886 7712
rect 11942 7656 12438 7712
rect 12494 7656 12499 7712
rect 11881 7654 12499 7656
rect 11881 7651 11947 7654
rect 12433 7651 12499 7654
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 13077 7442 13143 7445
rect 15837 7442 15903 7445
rect 17125 7442 17191 7445
rect 13077 7440 17191 7442
rect 13077 7384 13082 7440
rect 13138 7384 15842 7440
rect 15898 7384 17130 7440
rect 17186 7384 17191 7440
rect 13077 7382 17191 7384
rect 13077 7379 13143 7382
rect 15837 7379 15903 7382
rect 17125 7379 17191 7382
rect 15009 7306 15075 7309
rect 21081 7306 21147 7309
rect 15009 7304 21147 7306
rect 15009 7248 15014 7304
rect 15070 7248 21086 7304
rect 21142 7248 21147 7304
rect 15009 7246 21147 7248
rect 15009 7243 15075 7246
rect 21081 7243 21147 7246
rect 14549 7170 14615 7173
rect 17309 7170 17375 7173
rect 14549 7168 17375 7170
rect 14549 7112 14554 7168
rect 14610 7112 17314 7168
rect 17370 7112 17375 7168
rect 14549 7110 17375 7112
rect 14549 7107 14615 7110
rect 17309 7107 17375 7110
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 4797 7034 4863 7037
rect 6126 7034 6132 7036
rect 4797 7032 6132 7034
rect 4797 6976 4802 7032
rect 4858 6976 6132 7032
rect 4797 6974 6132 6976
rect 4797 6971 4863 6974
rect 6126 6972 6132 6974
rect 6196 6972 6202 7036
rect 2681 6898 2747 6901
rect 4102 6898 4108 6900
rect 2681 6896 4108 6898
rect 2681 6840 2686 6896
rect 2742 6840 4108 6896
rect 2681 6838 4108 6840
rect 2681 6835 2747 6838
rect 4102 6836 4108 6838
rect 4172 6836 4178 6900
rect 10041 6898 10107 6901
rect 13721 6900 13787 6901
rect 10174 6898 10180 6900
rect 10041 6896 10180 6898
rect 10041 6840 10046 6896
rect 10102 6840 10180 6896
rect 10041 6838 10180 6840
rect 10041 6835 10107 6838
rect 10174 6836 10180 6838
rect 10244 6836 10250 6900
rect 13670 6836 13676 6900
rect 13740 6898 13787 6900
rect 20069 6898 20135 6901
rect 21817 6898 21883 6901
rect 13740 6896 13832 6898
rect 13782 6840 13832 6896
rect 13740 6838 13832 6840
rect 20069 6896 21883 6898
rect 20069 6840 20074 6896
rect 20130 6840 21822 6896
rect 21878 6840 21883 6896
rect 20069 6838 21883 6840
rect 13740 6836 13787 6838
rect 13721 6835 13787 6836
rect 20069 6835 20135 6838
rect 21817 6835 21883 6838
rect 15837 6762 15903 6765
rect 18689 6762 18755 6765
rect 15837 6760 18755 6762
rect 15837 6704 15842 6760
rect 15898 6704 18694 6760
rect 18750 6704 18755 6760
rect 15837 6702 18755 6704
rect 15837 6699 15903 6702
rect 18689 6699 18755 6702
rect 20529 6762 20595 6765
rect 24301 6762 24367 6765
rect 26417 6762 26483 6765
rect 20529 6760 26483 6762
rect 20529 6704 20534 6760
rect 20590 6704 24306 6760
rect 24362 6704 26422 6760
rect 26478 6704 26483 6760
rect 20529 6702 26483 6704
rect 20529 6699 20595 6702
rect 24301 6699 24367 6702
rect 26417 6699 26483 6702
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 14590 6292 14596 6356
rect 14660 6354 14666 6356
rect 14825 6354 14891 6357
rect 14660 6352 14891 6354
rect 14660 6296 14830 6352
rect 14886 6296 14891 6352
rect 14660 6294 14891 6296
rect 14660 6292 14666 6294
rect 14825 6291 14891 6294
rect 10501 6218 10567 6221
rect 14917 6218 14983 6221
rect 17309 6218 17375 6221
rect 10501 6216 14842 6218
rect 10501 6160 10506 6216
rect 10562 6160 14842 6216
rect 10501 6158 14842 6160
rect 10501 6155 10567 6158
rect 14782 6082 14842 6158
rect 14917 6216 17375 6218
rect 14917 6160 14922 6216
rect 14978 6160 17314 6216
rect 17370 6160 17375 6216
rect 14917 6158 17375 6160
rect 14917 6155 14983 6158
rect 17309 6155 17375 6158
rect 17769 6218 17835 6221
rect 19793 6218 19859 6221
rect 22277 6218 22343 6221
rect 22553 6218 22619 6221
rect 17769 6216 22619 6218
rect 17769 6160 17774 6216
rect 17830 6160 19798 6216
rect 19854 6160 22282 6216
rect 22338 6160 22558 6216
rect 22614 6160 22619 6216
rect 17769 6158 22619 6160
rect 17769 6155 17835 6158
rect 19793 6155 19859 6158
rect 22277 6155 22343 6158
rect 22553 6155 22619 6158
rect 15009 6082 15075 6085
rect 14782 6080 15075 6082
rect 14782 6024 15014 6080
rect 15070 6024 15075 6080
rect 14782 6022 15075 6024
rect 15009 6019 15075 6022
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 0 5810 400 5840
rect 1761 5810 1827 5813
rect 0 5808 1827 5810
rect 0 5752 1766 5808
rect 1822 5752 1827 5808
rect 0 5750 1827 5752
rect 0 5720 400 5750
rect 1761 5747 1827 5750
rect 8293 5810 8359 5813
rect 9254 5810 9260 5812
rect 8293 5808 9260 5810
rect 8293 5752 8298 5808
rect 8354 5752 9260 5808
rect 8293 5750 9260 5752
rect 8293 5747 8359 5750
rect 9254 5748 9260 5750
rect 9324 5810 9330 5812
rect 15009 5810 15075 5813
rect 18413 5810 18479 5813
rect 9324 5750 13876 5810
rect 9324 5748 9330 5750
rect 12985 5674 13051 5677
rect 9630 5672 13051 5674
rect 9630 5616 12990 5672
rect 13046 5616 13051 5672
rect 9630 5614 13051 5616
rect 13816 5674 13876 5750
rect 15009 5808 18479 5810
rect 15009 5752 15014 5808
rect 15070 5752 18418 5808
rect 18474 5752 18479 5808
rect 15009 5750 18479 5752
rect 15009 5747 15075 5750
rect 18413 5747 18479 5750
rect 16573 5676 16639 5677
rect 16573 5674 16620 5676
rect 13816 5672 16620 5674
rect 13816 5616 16578 5672
rect 13816 5614 16620 5616
rect 9397 5538 9463 5541
rect 9630 5538 9690 5614
rect 12985 5611 13051 5614
rect 16573 5612 16620 5614
rect 16684 5612 16690 5676
rect 16573 5611 16639 5612
rect 9397 5536 9690 5538
rect 9397 5480 9402 5536
rect 9458 5480 9690 5536
rect 9397 5478 9690 5480
rect 9397 5475 9463 5478
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 12433 5266 12499 5269
rect 12893 5266 12959 5269
rect 13077 5266 13143 5269
rect 17585 5266 17651 5269
rect 12433 5264 17651 5266
rect 12433 5208 12438 5264
rect 12494 5208 12898 5264
rect 12954 5208 13082 5264
rect 13138 5208 17590 5264
rect 17646 5208 17651 5264
rect 12433 5206 17651 5208
rect 12433 5203 12499 5206
rect 12893 5203 12959 5206
rect 13077 5203 13143 5206
rect 17585 5203 17651 5206
rect 3141 5130 3207 5133
rect 7598 5130 7604 5132
rect 3141 5128 7604 5130
rect 3141 5072 3146 5128
rect 3202 5072 7604 5128
rect 3141 5070 7604 5072
rect 3141 5067 3207 5070
rect 7598 5068 7604 5070
rect 7668 5068 7674 5132
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 12157 4586 12223 4589
rect 18137 4586 18203 4589
rect 12157 4584 18203 4586
rect 12157 4528 12162 4584
rect 12218 4528 18142 4584
rect 18198 4528 18203 4584
rect 12157 4526 18203 4528
rect 12157 4523 12223 4526
rect 18137 4523 18203 4526
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 3049 4042 3115 4045
rect 7414 4042 7420 4044
rect 3049 4040 7420 4042
rect 3049 3984 3054 4040
rect 3110 3984 7420 4040
rect 3049 3982 7420 3984
rect 3049 3979 3115 3982
rect 7414 3980 7420 3982
rect 7484 3980 7490 4044
rect 4419 3840 4735 3841
rect 0 3770 400 3800
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 1301 3770 1367 3773
rect 0 3768 1367 3770
rect 0 3712 1306 3768
rect 1362 3712 1367 3768
rect 0 3710 1367 3712
rect 0 3680 400 3710
rect 1301 3707 1367 3710
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 12985 3090 13051 3093
rect 15009 3090 15075 3093
rect 17033 3090 17099 3093
rect 12985 3088 17099 3090
rect 12985 3032 12990 3088
rect 13046 3032 15014 3088
rect 15070 3032 17038 3088
rect 17094 3032 17099 3088
rect 12985 3030 17099 3032
rect 12985 3027 13051 3030
rect 15009 3027 15075 3030
rect 17033 3027 17099 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 3325 2684 3391 2685
rect 3325 2682 3372 2684
rect 3280 2680 3372 2682
rect 3280 2624 3330 2680
rect 3280 2622 3372 2624
rect 3325 2620 3372 2622
rect 3436 2620 3442 2684
rect 17309 2682 17375 2685
rect 17769 2682 17835 2685
rect 17309 2680 17835 2682
rect 17309 2624 17314 2680
rect 17370 2624 17774 2680
rect 17830 2624 17835 2680
rect 17309 2622 17835 2624
rect 3325 2619 3391 2620
rect 17309 2619 17375 2622
rect 17769 2619 17835 2622
rect 17309 2546 17375 2549
rect 18321 2546 18387 2549
rect 17309 2544 18387 2546
rect 17309 2488 17314 2544
rect 17370 2488 18326 2544
rect 18382 2488 18387 2544
rect 17309 2486 18387 2488
rect 17309 2483 17375 2486
rect 18321 2483 18387 2486
rect 17309 2274 17375 2277
rect 18965 2274 19031 2277
rect 17309 2272 19031 2274
rect 17309 2216 17314 2272
rect 17370 2216 18970 2272
rect 19026 2216 19031 2272
rect 17309 2214 19031 2216
rect 17309 2211 17375 2214
rect 18965 2211 19031 2214
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 3417 2002 3483 2005
rect 3550 2002 3556 2004
rect 3417 2000 3556 2002
rect 3417 1944 3422 2000
rect 3478 1944 3556 2000
rect 3417 1942 3556 1944
rect 3417 1939 3483 1942
rect 3550 1940 3556 1942
rect 3620 1940 3626 2004
rect 0 1730 400 1760
rect 2865 1730 2931 1733
rect 0 1728 2931 1730
rect 0 1672 2870 1728
rect 2926 1672 2931 1728
rect 0 1670 2931 1672
rect 0 1640 400 1670
rect 2865 1667 2931 1670
rect 4419 1664 4735 1665
rect 4419 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4735 1664
rect 4419 1599 4735 1600
rect 11365 1664 11681 1665
rect 11365 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11681 1664
rect 11365 1599 11681 1600
rect 18311 1664 18627 1665
rect 18311 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18627 1664
rect 18311 1599 18627 1600
rect 25257 1664 25573 1665
rect 25257 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25573 1664
rect 25257 1599 25573 1600
rect 12433 1458 12499 1461
rect 16113 1458 16179 1461
rect 21081 1458 21147 1461
rect 12433 1456 21147 1458
rect 12433 1400 12438 1456
rect 12494 1400 16118 1456
rect 16174 1400 21086 1456
rect 21142 1400 21147 1456
rect 12433 1398 21147 1400
rect 12433 1395 12499 1398
rect 16113 1395 16179 1398
rect 21081 1395 21147 1398
rect 3325 1322 3391 1325
rect 8886 1322 8892 1324
rect 3325 1320 8892 1322
rect 3325 1264 3330 1320
rect 3386 1264 8892 1320
rect 3325 1262 8892 1264
rect 3325 1259 3391 1262
rect 8886 1260 8892 1262
rect 8956 1260 8962 1324
rect 11973 1322 12039 1325
rect 12934 1322 12940 1324
rect 11973 1320 12940 1322
rect 11973 1264 11978 1320
rect 12034 1264 12940 1320
rect 11973 1262 12940 1264
rect 11973 1259 12039 1262
rect 12934 1260 12940 1262
rect 13004 1260 13010 1324
rect 7892 1120 8208 1121
rect 7892 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8208 1120
rect 7892 1055 8208 1056
rect 14838 1120 15154 1121
rect 14838 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15154 1120
rect 14838 1055 15154 1056
rect 21784 1120 22100 1121
rect 21784 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22100 1120
rect 21784 1055 22100 1056
rect 28730 1120 29046 1121
rect 28730 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29046 1120
rect 28730 1055 29046 1056
rect 2221 914 2287 917
rect 15878 914 15884 916
rect 2221 912 15884 914
rect 2221 856 2226 912
rect 2282 856 15884 912
rect 2221 854 15884 856
rect 2221 851 2287 854
rect 15878 852 15884 854
rect 15948 852 15954 916
rect 5349 778 5415 781
rect 11094 778 11100 780
rect 5349 776 11100 778
rect 5349 720 5354 776
rect 5410 720 11100 776
rect 5349 718 11100 720
rect 5349 715 5415 718
rect 11094 716 11100 718
rect 11164 716 11170 780
<< via3 >>
rect 7898 32668 7962 32672
rect 7898 32612 7902 32668
rect 7902 32612 7958 32668
rect 7958 32612 7962 32668
rect 7898 32608 7962 32612
rect 7978 32668 8042 32672
rect 7978 32612 7982 32668
rect 7982 32612 8038 32668
rect 8038 32612 8042 32668
rect 7978 32608 8042 32612
rect 8058 32668 8122 32672
rect 8058 32612 8062 32668
rect 8062 32612 8118 32668
rect 8118 32612 8122 32668
rect 8058 32608 8122 32612
rect 8138 32668 8202 32672
rect 8138 32612 8142 32668
rect 8142 32612 8198 32668
rect 8198 32612 8202 32668
rect 8138 32608 8202 32612
rect 14844 32668 14908 32672
rect 14844 32612 14848 32668
rect 14848 32612 14904 32668
rect 14904 32612 14908 32668
rect 14844 32608 14908 32612
rect 14924 32668 14988 32672
rect 14924 32612 14928 32668
rect 14928 32612 14984 32668
rect 14984 32612 14988 32668
rect 14924 32608 14988 32612
rect 15004 32668 15068 32672
rect 15004 32612 15008 32668
rect 15008 32612 15064 32668
rect 15064 32612 15068 32668
rect 15004 32608 15068 32612
rect 15084 32668 15148 32672
rect 15084 32612 15088 32668
rect 15088 32612 15144 32668
rect 15144 32612 15148 32668
rect 15084 32608 15148 32612
rect 21790 32668 21854 32672
rect 21790 32612 21794 32668
rect 21794 32612 21850 32668
rect 21850 32612 21854 32668
rect 21790 32608 21854 32612
rect 21870 32668 21934 32672
rect 21870 32612 21874 32668
rect 21874 32612 21930 32668
rect 21930 32612 21934 32668
rect 21870 32608 21934 32612
rect 21950 32668 22014 32672
rect 21950 32612 21954 32668
rect 21954 32612 22010 32668
rect 22010 32612 22014 32668
rect 21950 32608 22014 32612
rect 22030 32668 22094 32672
rect 22030 32612 22034 32668
rect 22034 32612 22090 32668
rect 22090 32612 22094 32668
rect 22030 32608 22094 32612
rect 28736 32668 28800 32672
rect 28736 32612 28740 32668
rect 28740 32612 28796 32668
rect 28796 32612 28800 32668
rect 28736 32608 28800 32612
rect 28816 32668 28880 32672
rect 28816 32612 28820 32668
rect 28820 32612 28876 32668
rect 28876 32612 28880 32668
rect 28816 32608 28880 32612
rect 28896 32668 28960 32672
rect 28896 32612 28900 32668
rect 28900 32612 28956 32668
rect 28956 32612 28960 32668
rect 28896 32608 28960 32612
rect 28976 32668 29040 32672
rect 28976 32612 28980 32668
rect 28980 32612 29036 32668
rect 29036 32612 29040 32668
rect 28976 32608 29040 32612
rect 4425 32124 4489 32128
rect 4425 32068 4429 32124
rect 4429 32068 4485 32124
rect 4485 32068 4489 32124
rect 4425 32064 4489 32068
rect 4505 32124 4569 32128
rect 4505 32068 4509 32124
rect 4509 32068 4565 32124
rect 4565 32068 4569 32124
rect 4505 32064 4569 32068
rect 4585 32124 4649 32128
rect 4585 32068 4589 32124
rect 4589 32068 4645 32124
rect 4645 32068 4649 32124
rect 4585 32064 4649 32068
rect 4665 32124 4729 32128
rect 4665 32068 4669 32124
rect 4669 32068 4725 32124
rect 4725 32068 4729 32124
rect 4665 32064 4729 32068
rect 11371 32124 11435 32128
rect 11371 32068 11375 32124
rect 11375 32068 11431 32124
rect 11431 32068 11435 32124
rect 11371 32064 11435 32068
rect 11451 32124 11515 32128
rect 11451 32068 11455 32124
rect 11455 32068 11511 32124
rect 11511 32068 11515 32124
rect 11451 32064 11515 32068
rect 11531 32124 11595 32128
rect 11531 32068 11535 32124
rect 11535 32068 11591 32124
rect 11591 32068 11595 32124
rect 11531 32064 11595 32068
rect 11611 32124 11675 32128
rect 11611 32068 11615 32124
rect 11615 32068 11671 32124
rect 11671 32068 11675 32124
rect 11611 32064 11675 32068
rect 18317 32124 18381 32128
rect 18317 32068 18321 32124
rect 18321 32068 18377 32124
rect 18377 32068 18381 32124
rect 18317 32064 18381 32068
rect 18397 32124 18461 32128
rect 18397 32068 18401 32124
rect 18401 32068 18457 32124
rect 18457 32068 18461 32124
rect 18397 32064 18461 32068
rect 18477 32124 18541 32128
rect 18477 32068 18481 32124
rect 18481 32068 18537 32124
rect 18537 32068 18541 32124
rect 18477 32064 18541 32068
rect 18557 32124 18621 32128
rect 18557 32068 18561 32124
rect 18561 32068 18617 32124
rect 18617 32068 18621 32124
rect 18557 32064 18621 32068
rect 25263 32124 25327 32128
rect 25263 32068 25267 32124
rect 25267 32068 25323 32124
rect 25323 32068 25327 32124
rect 25263 32064 25327 32068
rect 25343 32124 25407 32128
rect 25343 32068 25347 32124
rect 25347 32068 25403 32124
rect 25403 32068 25407 32124
rect 25343 32064 25407 32068
rect 25423 32124 25487 32128
rect 25423 32068 25427 32124
rect 25427 32068 25483 32124
rect 25483 32068 25487 32124
rect 25423 32064 25487 32068
rect 25503 32124 25567 32128
rect 25503 32068 25507 32124
rect 25507 32068 25563 32124
rect 25563 32068 25567 32124
rect 25503 32064 25567 32068
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7420 26284 7484 26348
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 10180 25332 10244 25396
rect 13124 25196 13188 25260
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 12940 24788 13004 24852
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 21404 22612 21468 22676
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 15884 20768 15948 20772
rect 15884 20712 15898 20768
rect 15898 20712 15948 20768
rect 15884 20708 15948 20712
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 7236 20436 7300 20500
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 16436 19892 16500 19956
rect 11100 19756 11164 19820
rect 6500 19680 6564 19684
rect 6500 19624 6550 19680
rect 6550 19624 6564 19680
rect 6500 19620 6564 19624
rect 9812 19680 9876 19684
rect 9812 19624 9826 19680
rect 9826 19624 9876 19680
rect 9812 19620 9876 19624
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 6132 19348 6196 19412
rect 20116 19348 20180 19412
rect 23428 19408 23492 19412
rect 23428 19352 23442 19408
rect 23442 19352 23492 19408
rect 23428 19348 23492 19352
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7236 18668 7300 18732
rect 8892 18532 8956 18596
rect 22324 18532 22388 18596
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 15700 17988 15764 18052
rect 20484 17988 20548 18052
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7604 17580 7668 17644
rect 6500 17444 6564 17508
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 9260 16688 9324 16692
rect 9260 16632 9310 16688
rect 9310 16632 9324 16688
rect 9260 16628 9324 16632
rect 11836 16628 11900 16692
rect 17724 16628 17788 16692
rect 9628 16492 9692 16556
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4108 15948 4172 16012
rect 6132 15948 6196 16012
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7420 15540 7484 15604
rect 9444 15600 9508 15604
rect 9444 15544 9458 15600
rect 9458 15544 9508 15600
rect 9444 15540 9508 15544
rect 18092 15540 18156 15604
rect 21404 15540 21468 15604
rect 14596 15404 14660 15468
rect 13860 15268 13924 15332
rect 17908 15268 17972 15332
rect 22508 15268 22572 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 3372 14996 3436 15060
rect 19932 14996 19996 15060
rect 7236 14860 7300 14924
rect 21036 14724 21100 14788
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 8892 14180 8956 14244
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 21036 13908 21100 13972
rect 9628 13772 9692 13836
rect 11836 13636 11900 13700
rect 17356 13636 17420 13700
rect 22324 13636 22388 13700
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 20300 13288 20364 13292
rect 20300 13232 20314 13288
rect 20314 13232 20364 13288
rect 20300 13228 20364 13232
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 16988 12956 17052 13020
rect 9444 12820 9508 12884
rect 22508 12820 22572 12884
rect 25820 12548 25884 12612
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 18092 12336 18156 12340
rect 18092 12280 18142 12336
rect 18142 12280 18156 12336
rect 18092 12276 18156 12280
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 23428 11868 23492 11932
rect 13860 11732 13924 11796
rect 17724 11732 17788 11796
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7420 11052 7484 11116
rect 9628 11052 9692 11116
rect 16620 11052 16684 11116
rect 21036 10976 21100 10980
rect 21036 10920 21050 10976
rect 21050 10920 21100 10976
rect 21036 10916 21100 10920
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 7236 9692 7300 9756
rect 20300 9828 20364 9892
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 19748 9556 19812 9620
rect 19932 9616 19996 9620
rect 19932 9560 19946 9616
rect 19946 9560 19996 9616
rect 19932 9556 19996 9560
rect 20300 9556 20364 9620
rect 20484 9420 20548 9484
rect 23428 9284 23492 9348
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 19748 9148 19812 9212
rect 15700 9072 15764 9076
rect 15700 9016 15714 9072
rect 15714 9016 15764 9072
rect 15700 9012 15764 9016
rect 16436 9012 16500 9076
rect 17356 9012 17420 9076
rect 25820 8740 25884 8804
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 13676 8332 13740 8396
rect 16988 8332 17052 8396
rect 17908 8196 17972 8260
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 20300 8060 20364 8124
rect 3556 7788 3620 7852
rect 13124 7788 13188 7852
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 6132 6972 6196 7036
rect 4108 6836 4172 6900
rect 10180 6836 10244 6900
rect 13676 6896 13740 6900
rect 13676 6840 13726 6896
rect 13726 6840 13740 6896
rect 13676 6836 13740 6840
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 14596 6292 14660 6356
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 9260 5748 9324 5812
rect 16620 5672 16684 5676
rect 16620 5616 16634 5672
rect 16634 5616 16684 5672
rect 16620 5612 16684 5616
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 7604 5068 7668 5132
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 7420 3980 7484 4044
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 3372 2680 3436 2684
rect 3372 2624 3386 2680
rect 3386 2624 3436 2680
rect 3372 2620 3436 2624
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
rect 3556 1940 3620 2004
rect 4425 1660 4489 1664
rect 4425 1604 4429 1660
rect 4429 1604 4485 1660
rect 4485 1604 4489 1660
rect 4425 1600 4489 1604
rect 4505 1660 4569 1664
rect 4505 1604 4509 1660
rect 4509 1604 4565 1660
rect 4565 1604 4569 1660
rect 4505 1600 4569 1604
rect 4585 1660 4649 1664
rect 4585 1604 4589 1660
rect 4589 1604 4645 1660
rect 4645 1604 4649 1660
rect 4585 1600 4649 1604
rect 4665 1660 4729 1664
rect 4665 1604 4669 1660
rect 4669 1604 4725 1660
rect 4725 1604 4729 1660
rect 4665 1600 4729 1604
rect 11371 1660 11435 1664
rect 11371 1604 11375 1660
rect 11375 1604 11431 1660
rect 11431 1604 11435 1660
rect 11371 1600 11435 1604
rect 11451 1660 11515 1664
rect 11451 1604 11455 1660
rect 11455 1604 11511 1660
rect 11511 1604 11515 1660
rect 11451 1600 11515 1604
rect 11531 1660 11595 1664
rect 11531 1604 11535 1660
rect 11535 1604 11591 1660
rect 11591 1604 11595 1660
rect 11531 1600 11595 1604
rect 11611 1660 11675 1664
rect 11611 1604 11615 1660
rect 11615 1604 11671 1660
rect 11671 1604 11675 1660
rect 11611 1600 11675 1604
rect 18317 1660 18381 1664
rect 18317 1604 18321 1660
rect 18321 1604 18377 1660
rect 18377 1604 18381 1660
rect 18317 1600 18381 1604
rect 18397 1660 18461 1664
rect 18397 1604 18401 1660
rect 18401 1604 18457 1660
rect 18457 1604 18461 1660
rect 18397 1600 18461 1604
rect 18477 1660 18541 1664
rect 18477 1604 18481 1660
rect 18481 1604 18537 1660
rect 18537 1604 18541 1660
rect 18477 1600 18541 1604
rect 18557 1660 18621 1664
rect 18557 1604 18561 1660
rect 18561 1604 18617 1660
rect 18617 1604 18621 1660
rect 18557 1600 18621 1604
rect 25263 1660 25327 1664
rect 25263 1604 25267 1660
rect 25267 1604 25323 1660
rect 25323 1604 25327 1660
rect 25263 1600 25327 1604
rect 25343 1660 25407 1664
rect 25343 1604 25347 1660
rect 25347 1604 25403 1660
rect 25403 1604 25407 1660
rect 25343 1600 25407 1604
rect 25423 1660 25487 1664
rect 25423 1604 25427 1660
rect 25427 1604 25483 1660
rect 25483 1604 25487 1660
rect 25423 1600 25487 1604
rect 25503 1660 25567 1664
rect 25503 1604 25507 1660
rect 25507 1604 25563 1660
rect 25563 1604 25567 1660
rect 25503 1600 25567 1604
rect 8892 1260 8956 1324
rect 12940 1260 13004 1324
rect 7898 1116 7962 1120
rect 7898 1060 7902 1116
rect 7902 1060 7958 1116
rect 7958 1060 7962 1116
rect 7898 1056 7962 1060
rect 7978 1116 8042 1120
rect 7978 1060 7982 1116
rect 7982 1060 8038 1116
rect 8038 1060 8042 1116
rect 7978 1056 8042 1060
rect 8058 1116 8122 1120
rect 8058 1060 8062 1116
rect 8062 1060 8118 1116
rect 8118 1060 8122 1116
rect 8058 1056 8122 1060
rect 8138 1116 8202 1120
rect 8138 1060 8142 1116
rect 8142 1060 8198 1116
rect 8198 1060 8202 1116
rect 8138 1056 8202 1060
rect 14844 1116 14908 1120
rect 14844 1060 14848 1116
rect 14848 1060 14904 1116
rect 14904 1060 14908 1116
rect 14844 1056 14908 1060
rect 14924 1116 14988 1120
rect 14924 1060 14928 1116
rect 14928 1060 14984 1116
rect 14984 1060 14988 1116
rect 14924 1056 14988 1060
rect 15004 1116 15068 1120
rect 15004 1060 15008 1116
rect 15008 1060 15064 1116
rect 15064 1060 15068 1116
rect 15004 1056 15068 1060
rect 15084 1116 15148 1120
rect 15084 1060 15088 1116
rect 15088 1060 15144 1116
rect 15144 1060 15148 1116
rect 15084 1056 15148 1060
rect 21790 1116 21854 1120
rect 21790 1060 21794 1116
rect 21794 1060 21850 1116
rect 21850 1060 21854 1116
rect 21790 1056 21854 1060
rect 21870 1116 21934 1120
rect 21870 1060 21874 1116
rect 21874 1060 21930 1116
rect 21930 1060 21934 1116
rect 21870 1056 21934 1060
rect 21950 1116 22014 1120
rect 21950 1060 21954 1116
rect 21954 1060 22010 1116
rect 22010 1060 22014 1116
rect 21950 1056 22014 1060
rect 22030 1116 22094 1120
rect 22030 1060 22034 1116
rect 22034 1060 22090 1116
rect 22090 1060 22094 1116
rect 22030 1056 22094 1060
rect 28736 1116 28800 1120
rect 28736 1060 28740 1116
rect 28740 1060 28796 1116
rect 28796 1060 28800 1116
rect 28736 1056 28800 1060
rect 28816 1116 28880 1120
rect 28816 1060 28820 1116
rect 28820 1060 28876 1116
rect 28876 1060 28880 1116
rect 28816 1056 28880 1060
rect 28896 1116 28960 1120
rect 28896 1060 28900 1116
rect 28900 1060 28956 1116
rect 28956 1060 28960 1116
rect 28896 1056 28960 1060
rect 28976 1116 29040 1120
rect 28976 1060 28980 1116
rect 28980 1060 29036 1116
rect 29036 1060 29040 1116
rect 28976 1056 29040 1060
rect 15884 852 15948 916
rect 11100 716 11164 780
<< metal4 >>
rect 4417 32128 4737 32688
rect 4417 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4737 32128
rect 4417 31040 4737 32064
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 7890 32672 8210 32688
rect 7890 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8210 32672
rect 7890 31584 8210 32608
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7419 26348 7485 26349
rect 7419 26284 7420 26348
rect 7484 26284 7485 26348
rect 7419 26283 7485 26284
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 7235 20500 7301 20501
rect 7235 20436 7236 20500
rect 7300 20436 7301 20500
rect 7235 20435 7301 20436
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 6499 19684 6565 19685
rect 6499 19620 6500 19684
rect 6564 19620 6565 19684
rect 6499 19619 6565 19620
rect 6131 19412 6197 19413
rect 6131 19348 6132 19412
rect 6196 19348 6197 19412
rect 6131 19347 6197 19348
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4107 16012 4173 16013
rect 4107 15948 4108 16012
rect 4172 15948 4173 16012
rect 4107 15947 4173 15948
rect 3371 15060 3437 15061
rect 3371 14996 3372 15060
rect 3436 14996 3437 15060
rect 3371 14995 3437 14996
rect 3374 2685 3434 14995
rect 3555 7852 3621 7853
rect 3555 7788 3556 7852
rect 3620 7788 3621 7852
rect 3555 7787 3621 7788
rect 3371 2684 3437 2685
rect 3371 2620 3372 2684
rect 3436 2620 3437 2684
rect 3371 2619 3437 2620
rect 3558 2005 3618 7787
rect 4110 6901 4170 15947
rect 4417 15808 4737 16832
rect 6134 16013 6194 19347
rect 6502 17509 6562 19619
rect 7238 18733 7298 20435
rect 7235 18732 7301 18733
rect 7235 18668 7236 18732
rect 7300 18668 7301 18732
rect 7235 18667 7301 18668
rect 6499 17508 6565 17509
rect 6499 17444 6500 17508
rect 6564 17444 6565 17508
rect 6499 17443 6565 17444
rect 6131 16012 6197 16013
rect 6131 15948 6132 16012
rect 6196 15948 6197 16012
rect 6131 15947 6197 15948
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4107 6900 4173 6901
rect 4107 6836 4108 6900
rect 4172 6836 4173 6900
rect 4107 6835 4173 6836
rect 4417 6016 4737 7040
rect 6134 7037 6194 15947
rect 7238 14925 7298 18667
rect 7422 15605 7482 26283
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 11363 32128 11683 32688
rect 11363 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11683 32128
rect 11363 31040 11683 32064
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 10179 25396 10245 25397
rect 10179 25332 10180 25396
rect 10244 25332 10245 25396
rect 10179 25331 10245 25332
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 9811 19684 9877 19685
rect 9811 19620 9812 19684
rect 9876 19620 9877 19684
rect 9811 19619 9877 19620
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 9814 19350 9874 19619
rect 9630 19290 9874 19350
rect 8891 18596 8957 18597
rect 8891 18532 8892 18596
rect 8956 18532 8957 18596
rect 8891 18531 8957 18532
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7603 17644 7669 17645
rect 7603 17580 7604 17644
rect 7668 17580 7669 17644
rect 7603 17579 7669 17580
rect 7419 15604 7485 15605
rect 7419 15540 7420 15604
rect 7484 15540 7485 15604
rect 7419 15539 7485 15540
rect 7235 14924 7301 14925
rect 7235 14860 7236 14924
rect 7300 14860 7301 14924
rect 7235 14859 7301 14860
rect 7238 9757 7298 14859
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 7235 9756 7301 9757
rect 7235 9692 7236 9756
rect 7300 9692 7301 9756
rect 7235 9691 7301 9692
rect 6131 7036 6197 7037
rect 6131 6972 6132 7036
rect 6196 6972 6197 7036
rect 6131 6971 6197 6972
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 7422 4045 7482 11051
rect 7606 5133 7666 17579
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 8894 14245 8954 18531
rect 9259 16692 9325 16693
rect 9259 16628 9260 16692
rect 9324 16628 9325 16692
rect 9259 16627 9325 16628
rect 8891 14244 8957 14245
rect 8891 14180 8892 14244
rect 8956 14180 8957 14244
rect 8891 14179 8957 14180
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7603 5132 7669 5133
rect 7603 5068 7604 5132
rect 7668 5068 7669 5132
rect 7603 5067 7669 5068
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 3555 2004 3621 2005
rect 3555 1940 3556 2004
rect 3620 1940 3621 2004
rect 3555 1939 3621 1940
rect 4417 1664 4737 2688
rect 4417 1600 4425 1664
rect 4489 1600 4505 1664
rect 4569 1600 4585 1664
rect 4649 1600 4665 1664
rect 4729 1600 4737 1664
rect 4417 1040 4737 1600
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 1120 8210 2144
rect 8894 1325 8954 14179
rect 9262 5813 9322 16627
rect 9630 16557 9690 19290
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9443 15604 9509 15605
rect 9443 15540 9444 15604
rect 9508 15540 9509 15604
rect 9443 15539 9509 15540
rect 9446 12885 9506 15539
rect 9627 13836 9693 13837
rect 9627 13772 9628 13836
rect 9692 13772 9693 13836
rect 9627 13771 9693 13772
rect 9443 12884 9509 12885
rect 9443 12820 9444 12884
rect 9508 12820 9509 12884
rect 9443 12819 9509 12820
rect 9630 11117 9690 13771
rect 9627 11116 9693 11117
rect 9627 11052 9628 11116
rect 9692 11052 9693 11116
rect 9627 11051 9693 11052
rect 10182 6901 10242 25331
rect 11363 24512 11683 25536
rect 14836 32672 15156 32688
rect 14836 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15156 32672
rect 14836 31584 15156 32608
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 13123 25260 13189 25261
rect 13123 25196 13124 25260
rect 13188 25196 13189 25260
rect 13123 25195 13189 25196
rect 12939 24852 13005 24853
rect 12939 24788 12940 24852
rect 13004 24788 13005 24852
rect 12939 24787 13005 24788
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11099 19820 11165 19821
rect 11099 19756 11100 19820
rect 11164 19756 11165 19820
rect 11099 19755 11165 19756
rect 10179 6900 10245 6901
rect 10179 6836 10180 6900
rect 10244 6836 10245 6900
rect 10179 6835 10245 6836
rect 9259 5812 9325 5813
rect 9259 5748 9260 5812
rect 9324 5748 9325 5812
rect 9259 5747 9325 5748
rect 8891 1324 8957 1325
rect 8891 1260 8892 1324
rect 8956 1260 8957 1324
rect 8891 1259 8957 1260
rect 7890 1056 7898 1120
rect 7962 1056 7978 1120
rect 8042 1056 8058 1120
rect 8122 1056 8138 1120
rect 8202 1056 8210 1120
rect 7890 1040 8210 1056
rect 11102 781 11162 19755
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11835 16692 11901 16693
rect 11835 16628 11836 16692
rect 11900 16628 11901 16692
rect 11835 16627 11901 16628
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11838 13701 11898 16627
rect 11835 13700 11901 13701
rect 11835 13636 11836 13700
rect 11900 13636 11901 13700
rect 11835 13635 11901 13636
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 1664 11683 2688
rect 11363 1600 11371 1664
rect 11435 1600 11451 1664
rect 11515 1600 11531 1664
rect 11595 1600 11611 1664
rect 11675 1600 11683 1664
rect 11363 1040 11683 1600
rect 12942 1325 13002 24787
rect 13126 7853 13186 25195
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 18309 32128 18629 32688
rect 18309 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18629 32128
rect 18309 31040 18629 32064
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 21782 32672 22102 32688
rect 21782 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22102 32672
rect 21782 31584 22102 32608
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21403 22676 21469 22677
rect 21403 22612 21404 22676
rect 21468 22612 21469 22676
rect 21403 22611 21469 22612
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 15699 18052 15765 18053
rect 15699 17988 15700 18052
rect 15764 17988 15765 18052
rect 15699 17987 15765 17988
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14595 15468 14661 15469
rect 14595 15404 14596 15468
rect 14660 15404 14661 15468
rect 14595 15403 14661 15404
rect 13859 15332 13925 15333
rect 13859 15268 13860 15332
rect 13924 15268 13925 15332
rect 13859 15267 13925 15268
rect 13862 11797 13922 15267
rect 13859 11796 13925 11797
rect 13859 11732 13860 11796
rect 13924 11732 13925 11796
rect 13859 11731 13925 11732
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 13123 7852 13189 7853
rect 13123 7788 13124 7852
rect 13188 7788 13189 7852
rect 13123 7787 13189 7788
rect 13678 6901 13738 8331
rect 13675 6900 13741 6901
rect 13675 6836 13676 6900
rect 13740 6836 13741 6900
rect 13675 6835 13741 6836
rect 14598 6357 14658 15403
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 15702 9077 15762 17987
rect 15699 9076 15765 9077
rect 15699 9012 15700 9076
rect 15764 9012 15765 9076
rect 15699 9011 15765 9012
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14595 6356 14661 6357
rect 14595 6292 14596 6356
rect 14660 6292 14661 6356
rect 14595 6291 14661 6292
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 12939 1324 13005 1325
rect 12939 1260 12940 1324
rect 13004 1260 13005 1324
rect 12939 1259 13005 1260
rect 14836 1120 15156 2144
rect 14836 1056 14844 1120
rect 14908 1056 14924 1120
rect 14988 1056 15004 1120
rect 15068 1056 15084 1120
rect 15148 1056 15156 1120
rect 14836 1040 15156 1056
rect 15886 917 15946 20707
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 16435 19956 16501 19957
rect 16435 19892 16436 19956
rect 16500 19892 16501 19956
rect 16435 19891 16501 19892
rect 16438 9077 16498 19891
rect 18309 19072 18629 20096
rect 20115 19412 20181 19413
rect 20115 19348 20116 19412
rect 20180 19348 20181 19412
rect 20115 19347 20181 19348
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 20118 17970 20178 19347
rect 20483 18052 20549 18053
rect 20483 17988 20484 18052
rect 20548 17988 20549 18052
rect 20483 17987 20549 17988
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17355 13700 17421 13701
rect 17355 13636 17356 13700
rect 17420 13636 17421 13700
rect 17355 13635 17421 13636
rect 16987 13020 17053 13021
rect 16987 12956 16988 13020
rect 17052 12956 17053 13020
rect 16987 12955 17053 12956
rect 16619 11116 16685 11117
rect 16619 11052 16620 11116
rect 16684 11052 16685 11116
rect 16619 11051 16685 11052
rect 16435 9076 16501 9077
rect 16435 9012 16436 9076
rect 16500 9012 16501 9076
rect 16435 9011 16501 9012
rect 16622 5677 16682 11051
rect 16990 8397 17050 12955
rect 17358 9077 17418 13635
rect 17726 11797 17786 16627
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18091 15604 18157 15605
rect 18091 15540 18092 15604
rect 18156 15540 18157 15604
rect 18091 15539 18157 15540
rect 17907 15332 17973 15333
rect 17907 15268 17908 15332
rect 17972 15268 17973 15332
rect 17907 15267 17973 15268
rect 17723 11796 17789 11797
rect 17723 11732 17724 11796
rect 17788 11732 17789 11796
rect 17723 11731 17789 11732
rect 17355 9076 17421 9077
rect 17355 9012 17356 9076
rect 17420 9012 17421 9076
rect 17355 9011 17421 9012
rect 16987 8396 17053 8397
rect 16987 8332 16988 8396
rect 17052 8332 17053 8396
rect 16987 8331 17053 8332
rect 17910 8261 17970 15267
rect 18094 12341 18154 15539
rect 18309 14720 18629 15744
rect 19934 17910 20178 17970
rect 19934 15061 19994 17910
rect 19931 15060 19997 15061
rect 19931 14996 19932 15060
rect 19996 14996 19997 15060
rect 19931 14995 19997 14996
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18091 12340 18157 12341
rect 18091 12276 18092 12340
rect 18156 12276 18157 12340
rect 18091 12275 18157 12276
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 19934 9621 19994 14995
rect 20299 13292 20365 13293
rect 20299 13228 20300 13292
rect 20364 13228 20365 13292
rect 20299 13227 20365 13228
rect 20302 9893 20362 13227
rect 20299 9892 20365 9893
rect 20299 9828 20300 9892
rect 20364 9828 20365 9892
rect 20299 9827 20365 9828
rect 19747 9620 19813 9621
rect 19747 9556 19748 9620
rect 19812 9556 19813 9620
rect 19747 9555 19813 9556
rect 19931 9620 19997 9621
rect 19931 9556 19932 9620
rect 19996 9556 19997 9620
rect 19931 9555 19997 9556
rect 20299 9620 20365 9621
rect 20299 9556 20300 9620
rect 20364 9556 20365 9620
rect 20299 9555 20365 9556
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 17907 8260 17973 8261
rect 17907 8196 17908 8260
rect 17972 8196 17973 8260
rect 17907 8195 17973 8196
rect 18309 8192 18629 9216
rect 19750 9213 19810 9555
rect 19747 9212 19813 9213
rect 19747 9148 19748 9212
rect 19812 9148 19813 9212
rect 19747 9147 19813 9148
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 20302 8125 20362 9555
rect 20486 9485 20546 17987
rect 21406 15605 21466 22611
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 25255 32128 25575 32688
rect 25255 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25575 32128
rect 25255 31040 25575 32064
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 23427 19412 23493 19413
rect 23427 19348 23428 19412
rect 23492 19348 23493 19412
rect 23427 19347 23493 19348
rect 22323 18596 22389 18597
rect 22323 18532 22324 18596
rect 22388 18532 22389 18596
rect 22323 18531 22389 18532
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21403 15604 21469 15605
rect 21403 15540 21404 15604
rect 21468 15540 21469 15604
rect 21403 15539 21469 15540
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21035 14788 21101 14789
rect 21035 14724 21036 14788
rect 21100 14724 21101 14788
rect 21035 14723 21101 14724
rect 21038 13973 21098 14723
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21035 13972 21101 13973
rect 21035 13908 21036 13972
rect 21100 13908 21101 13972
rect 21035 13907 21101 13908
rect 21038 10981 21098 13907
rect 21782 13088 22102 14112
rect 22326 13701 22386 18531
rect 22507 15332 22573 15333
rect 22507 15268 22508 15332
rect 22572 15268 22573 15332
rect 22507 15267 22573 15268
rect 22323 13700 22389 13701
rect 22323 13636 22324 13700
rect 22388 13636 22389 13700
rect 22323 13635 22389 13636
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 22510 12885 22570 15267
rect 22507 12884 22573 12885
rect 22507 12820 22508 12884
rect 22572 12820 22573 12884
rect 22507 12819 22573 12820
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21035 10980 21101 10981
rect 21035 10916 21036 10980
rect 21100 10916 21101 10980
rect 21035 10915 21101 10916
rect 21782 10912 22102 11936
rect 23430 11933 23490 19347
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 28728 32672 29048 32688
rect 28728 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29048 32672
rect 28728 31584 29048 32608
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 25819 12612 25885 12613
rect 25819 12548 25820 12612
rect 25884 12548 25885 12612
rect 25819 12547 25885 12548
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 23427 11932 23493 11933
rect 23427 11868 23428 11932
rect 23492 11868 23493 11932
rect 23427 11867 23493 11868
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 20483 9484 20549 9485
rect 20483 9420 20484 9484
rect 20548 9420 20549 9484
rect 20483 9419 20549 9420
rect 21782 8736 22102 9760
rect 23430 9349 23490 11867
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 23427 9348 23493 9349
rect 23427 9284 23428 9348
rect 23492 9284 23493 9348
rect 23427 9283 23493 9284
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 20299 8124 20365 8125
rect 20299 8060 20300 8124
rect 20364 8060 20365 8124
rect 20299 8059 20365 8060
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 16619 5676 16685 5677
rect 16619 5612 16620 5676
rect 16684 5612 16685 5676
rect 16619 5611 16685 5612
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 1664 18629 2688
rect 18309 1600 18317 1664
rect 18381 1600 18397 1664
rect 18461 1600 18477 1664
rect 18541 1600 18557 1664
rect 18621 1600 18629 1664
rect 18309 1040 18629 1600
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 1120 22102 2144
rect 21782 1056 21790 1120
rect 21854 1056 21870 1120
rect 21934 1056 21950 1120
rect 22014 1056 22030 1120
rect 22094 1056 22102 1120
rect 21782 1040 22102 1056
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25822 8805 25882 12547
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 25819 8804 25885 8805
rect 25819 8740 25820 8804
rect 25884 8740 25885 8804
rect 25819 8739 25885 8740
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 1664 25575 2688
rect 25255 1600 25263 1664
rect 25327 1600 25343 1664
rect 25407 1600 25423 1664
rect 25487 1600 25503 1664
rect 25567 1600 25575 1664
rect 25255 1040 25575 1600
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 1120 29048 2144
rect 28728 1056 28736 1120
rect 28800 1056 28816 1120
rect 28880 1056 28896 1120
rect 28960 1056 28976 1120
rect 29040 1056 29048 1120
rect 28728 1040 29048 1056
rect 15883 916 15949 917
rect 15883 852 15884 916
rect 15948 852 15949 916
rect 15883 851 15949 852
rect 11099 780 11165 781
rect 11099 716 11100 780
rect 11164 716 11165 780
rect 11099 715 11165 716
use sky130_fd_sc_hd__buf_2  _0438_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0439_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _0440_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0441_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0442_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0443_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0444_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0445_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0446_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0447_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0448_
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0449_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0450_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0451_
timestamp 1676037725
transform 1 0 7912 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1676037725
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0453_
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0454_
timestamp 1676037725
transform 1 0 5520 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0455_
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0456_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _0457_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _0458_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0459_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0460_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0461_
timestamp 1676037725
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0462_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0463_
timestamp 1676037725
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0464_
timestamp 1676037725
transform 1 0 2024 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0465_
timestamp 1676037725
transform 1 0 3496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1676037725
transform 1 0 7728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0467_
timestamp 1676037725
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0468_
timestamp 1676037725
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0469_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0470_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0471_
timestamp 1676037725
transform 1 0 9476 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0472_
timestamp 1676037725
transform 1 0 8832 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0473_
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0474_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0475_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0476_
timestamp 1676037725
transform 1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0477_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0478_
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0480_
timestamp 1676037725
transform 1 0 11408 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0481_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0482_
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0483_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0484_
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0485_
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_2  _0486_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0487_
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0488_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0489_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0490_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _0491_
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0492_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_2  _0493_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0494_
timestamp 1676037725
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0495_
timestamp 1676037725
transform 1 0 19964 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0496_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0497_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0498_
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0499_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _0500_
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0501_
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0502_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0503_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0504_
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0505_
timestamp 1676037725
transform 1 0 22632 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0506_
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0507_
timestamp 1676037725
transform 1 0 7268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0508_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0509_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0510_
timestamp 1676037725
transform 1 0 18584 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0511_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0512_
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0513_
timestamp 1676037725
transform 1 0 9568 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _0514_
timestamp 1676037725
transform 1 0 13248 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0515_
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0516_
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0517_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_2  _0518_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0519_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0520_
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0521_
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0522_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0523_
timestamp 1676037725
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0524_
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0525_
timestamp 1676037725
transform 1 0 12420 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0526_
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0527_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0528_
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _0529_
timestamp 1676037725
transform 1 0 10120 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0530_
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0531_
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0532_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0533_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0534_
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0535_
timestamp 1676037725
transform 1 0 12328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0536_
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0537_
timestamp 1676037725
transform 1 0 11224 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0538_
timestamp 1676037725
transform 1 0 13524 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0539_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0540_
timestamp 1676037725
transform 1 0 15732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0541_
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0542_
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0543_
timestamp 1676037725
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0544_
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0545_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0546_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0547_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0548_
timestamp 1676037725
transform 1 0 20240 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0549_
timestamp 1676037725
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0550_
timestamp 1676037725
transform 1 0 20884 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0551_
timestamp 1676037725
transform 1 0 17296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1676037725
transform 1 0 23460 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0553_
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0554_
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1676037725
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0556_
timestamp 1676037725
transform 1 0 15088 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0557_
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0558_
timestamp 1676037725
transform 1 0 24840 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0559_
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0560_
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0561_
timestamp 1676037725
transform 1 0 19504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0562_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0563_
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0564_
timestamp 1676037725
transform 1 0 20792 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0565_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0566_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0567_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0569_
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0570_
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0571_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0572_
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0573_
timestamp 1676037725
transform 1 0 24288 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0574_
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0575_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0576_
timestamp 1676037725
transform 1 0 23552 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0577_
timestamp 1676037725
transform 1 0 17112 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0578_
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0579_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0580_
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0581_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0582_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0583_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0584_
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0585_
timestamp 1676037725
transform 1 0 19412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0586_
timestamp 1676037725
transform 1 0 12696 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0587_
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0588_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0589_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0590_
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0591_
timestamp 1676037725
transform 1 0 14628 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp 1676037725
transform 1 0 15732 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0593_
timestamp 1676037725
transform 1 0 19872 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0594_
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0595_
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0596_
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_2  _0597_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9200 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0598_
timestamp 1676037725
transform 1 0 14628 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0599_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0600_
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0601_
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0602_
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0603_
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0605_
timestamp 1676037725
transform 1 0 17204 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0606_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0607_
timestamp 1676037725
transform 1 0 19412 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0608_
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0609_
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0610_
timestamp 1676037725
transform 1 0 13524 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0611_
timestamp 1676037725
transform 1 0 13156 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0612_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0613_
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0614_
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0616_
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0617_
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0618_
timestamp 1676037725
transform 1 0 22724 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0619_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0620_
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0621_
timestamp 1676037725
transform 1 0 23276 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0622_
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0623_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22356 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0624_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0625_
timestamp 1676037725
transform 1 0 10028 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0626_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 1676037725
transform 1 0 20884 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0628_
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0629_
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0630_
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0632_
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0633_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0634_
timestamp 1676037725
transform 1 0 17940 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1676037725
transform 1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0636_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0637_
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 1676037725
transform 1 0 11684 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0641_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14352 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0642_
timestamp 1676037725
transform 1 0 15456 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0643_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0644_
timestamp 1676037725
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0645_
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0646_
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0647_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0648_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0649_
timestamp 1676037725
transform 1 0 20148 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0650_
timestamp 1676037725
transform 1 0 25484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0651_
timestamp 1676037725
transform 1 0 22172 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _0652_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0653_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0654_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0655_
timestamp 1676037725
transform 1 0 8096 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0656_
timestamp 1676037725
transform 1 0 6532 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0657_
timestamp 1676037725
transform 1 0 6348 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0658_
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0659_
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0660_
timestamp 1676037725
transform 1 0 25668 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0661_
timestamp 1676037725
transform 1 0 20608 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0662_
timestamp 1676037725
transform 1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0663_
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0664_
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0665_
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0666_
timestamp 1676037725
transform 1 0 21804 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0667_
timestamp 1676037725
transform 1 0 16008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0668_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0669_
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0670_
timestamp 1676037725
transform 1 0 15732 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0671_
timestamp 1676037725
transform 1 0 14720 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0672_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0673_
timestamp 1676037725
transform 1 0 11960 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0674_
timestamp 1676037725
transform 1 0 11500 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0675_
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0676_
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0677_
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0678_
timestamp 1676037725
transform 1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0679_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _0680_
timestamp 1676037725
transform 1 0 7176 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0681_
timestamp 1676037725
transform 1 0 7176 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0682_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1676037725
transform 1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0684_
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0686_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0687_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0688_
timestamp 1676037725
transform 1 0 5428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0689_
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0690_
timestamp 1676037725
transform 1 0 5520 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_2  _0691_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _0692_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0694_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0695_
timestamp 1676037725
transform 1 0 4140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0696_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0697_
timestamp 1676037725
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _0698_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0699_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1676037725
transform 1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1676037725
transform 1 0 4784 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0702_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0703_
timestamp 1676037725
transform 1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0705_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 1676037725
transform 1 0 5244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0707_
timestamp 1676037725
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0708_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0709_
timestamp 1676037725
transform 1 0 5704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _0710_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5336 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0711_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0712_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0713_
timestamp 1676037725
transform 1 0 5612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _0714_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0715_
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0716_
timestamp 1676037725
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0717_
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _0718_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _0719_
timestamp 1676037725
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0720_
timestamp 1676037725
transform 1 0 2760 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0721_
timestamp 1676037725
transform 1 0 3128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0722_
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0724_
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0725_
timestamp 1676037725
transform 1 0 3864 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0726_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0727_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0728_
timestamp 1676037725
transform 1 0 10028 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1676037725
transform 1 0 8832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0730_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0731_
timestamp 1676037725
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0732_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0733_
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0734_
timestamp 1676037725
transform 1 0 5520 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0735_
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0736_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0737_
timestamp 1676037725
transform 1 0 8188 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0738_
timestamp 1676037725
transform 1 0 12696 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0739_
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0740_
timestamp 1676037725
transform 1 0 6532 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0741_
timestamp 1676037725
transform 1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _0742_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_2  _0743_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0745_
timestamp 1676037725
transform 1 0 6624 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1676037725
transform 1 0 9384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0747_
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0748_
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0749_
timestamp 1676037725
transform 1 0 10304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0750_
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0752_
timestamp 1676037725
transform 1 0 6532 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_2  _0753_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_2  _0754_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0755_
timestamp 1676037725
transform 1 0 5612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0756_
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0758_
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0759_
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0760_
timestamp 1676037725
transform 1 0 7636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0762_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0763_
timestamp 1676037725
transform 1 0 8096 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0764_
timestamp 1676037725
transform 1 0 5244 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _0765_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0766_
timestamp 1676037725
transform 1 0 12696 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0767_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0768_
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0770_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0771_
timestamp 1676037725
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0772_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0773_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _0774_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0775_
timestamp 1676037725
transform 1 0 11868 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0776_
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0777_
timestamp 1676037725
transform 1 0 5060 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0778_
timestamp 1676037725
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0779_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0780_
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0781_
timestamp 1676037725
transform 1 0 4784 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0782_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0783_
timestamp 1676037725
transform 1 0 5520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 1676037725
transform 1 0 6992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0785_
timestamp 1676037725
transform 1 0 7360 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0786_
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0787_
timestamp 1676037725
transform 1 0 6532 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0788_
timestamp 1676037725
transform 1 0 5704 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0789_
timestamp 1676037725
transform 1 0 6532 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0791_
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1676037725
transform 1 0 7544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0794_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0795_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1676037725
transform 1 0 6808 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0797_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _0798_
timestamp 1676037725
transform 1 0 3956 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0799_
timestamp 1676037725
transform 1 0 11040 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0800_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0801_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0802_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1676037725
transform 1 0 6256 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 1676037725
transform 1 0 4784 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0805_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0806_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0807_
timestamp 1676037725
transform 1 0 6532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0808_
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0809_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1676037725
transform 1 0 5796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0811_
timestamp 1676037725
transform 1 0 3220 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0812_
timestamp 1676037725
transform 1 0 5336 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0813_
timestamp 1676037725
transform 1 0 4784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0814_
timestamp 1676037725
transform 1 0 3956 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1676037725
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0817_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1676037725
transform 1 0 7360 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 1676037725
transform 1 0 9568 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1676037725
transform 1 0 8004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0821_
timestamp 1676037725
transform 1 0 7360 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0823_
timestamp 1676037725
transform 1 0 11684 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1676037725
transform 1 0 12972 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1676037725
transform 1 0 6532 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0826_
timestamp 1676037725
transform 1 0 6624 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0827_
timestamp 1676037725
transform 1 0 7452 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1676037725
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0829_
timestamp 1676037725
transform 1 0 11592 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 1676037725
transform 1 0 11868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _0831_
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1676037725
transform 1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0833_
timestamp 1676037725
transform 1 0 5796 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0834_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _0835_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _0836_
timestamp 1676037725
transform 1 0 1748 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _0837_
timestamp 1676037725
transform 1 0 6900 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _0838_
timestamp 1676037725
transform 1 0 2576 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0839_
timestamp 1676037725
transform 1 0 5520 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0840_
timestamp 1676037725
transform 1 0 4324 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0841_
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0842_
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0843_
timestamp 1676037725
transform 1 0 1748 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0844_
timestamp 1676037725
transform 1 0 4784 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _0845_
timestamp 1676037725
transform 1 0 3956 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a21boi_1  _0846_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_2  _0847_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0848_
timestamp 1676037725
transform 1 0 12328 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0849_
timestamp 1676037725
transform 1 0 12052 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _0850_
timestamp 1676037725
transform 1 0 12788 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0851_
timestamp 1676037725
transform 1 0 3772 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0852_
timestamp 1676037725
transform 1 0 14352 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0853_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _0854_
timestamp 1676037725
transform 1 0 25668 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0855_
timestamp 1676037725
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1676037725
transform 1 0 13248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0857_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0858_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0859_
timestamp 1676037725
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0861_
timestamp 1676037725
transform 1 0 15824 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0862_
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_2  _0863_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0864_
timestamp 1676037725
transform 1 0 13984 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0865_
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0867_
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0868_
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0870_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1676037725
transform 1 0 4140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _0872_
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 1676037725
transform 1 0 2944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1676037725
transform 1 0 4232 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0875_
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0876_
timestamp 1676037725
transform 1 0 3128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0877_
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _0880_
timestamp 1676037725
transform 1 0 9200 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1676037725
transform 1 0 11776 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0882_
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _0883_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4508 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1676037725
transform 1 0 6624 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1676037725
transform 1 0 4600 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1676037725
transform 1 0 6440 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1676037725
transform 1 0 8280 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1676037725
transform 1 0 11408 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1676037725
transform 1 0 25208 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1676037725
transform 1 0 26956 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1676037725
transform 1 0 25116 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1676037725
transform 1 0 23276 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1676037725
transform 1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1676037725
transform 1 0 9200 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1676037725
transform 1 0 7912 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1676037725
transform 1 0 4140 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1676037725
transform 1 0 7268 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1676037725
transform 1 0 2668 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1676037725
transform 1 0 9108 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1676037725
transform 1 0 6716 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1676037725
transform 1 0 7912 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1676037725
transform 1 0 11316 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1676037725
transform 1 0 14076 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1676037725
transform 1 0 12420 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1676037725
transform 1 0 9568 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1676037725
transform 1 0 14720 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1676037725
transform 1 0 25024 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1676037725
transform 1 0 26956 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1676037725
transform 1 0 23828 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1676037725
transform 1 0 16376 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1676037725
transform 1 0 7636 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1676037725
transform 1 0 22356 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1676037725
transform 1 0 20792 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1676037725
transform 1 0 19136 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1676037725
transform 1 0 17296 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1676037725
transform 1 0 16928 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1676037725
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1676037725
transform 1 0 9752 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1676037725
transform 1 0 12512 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1676037725
transform 1 0 10856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1676037725
transform 1 0 12328 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1676037725
transform 1 0 13248 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1676037725
transform 1 0 9752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1676037725
transform 1 0 14536 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1676037725
transform 1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1676037725
transform 1 0 9384 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1676037725
transform 1 0 9844 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1676037725
transform 1 0 23000 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1676037725
transform 1 0 22356 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1676037725
transform 1 0 19136 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1676037725
transform 1 0 19504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1676037725
transform 1 0 20516 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1676037725
transform 1 0 23276 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1676037725
transform 1 0 23828 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1676037725
transform 1 0 22356 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1676037725
transform 1 0 21988 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1676037725
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1676037725
transform 1 0 20148 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1676037725
transform 1 0 12880 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1676037725
transform 1 0 11316 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 11316 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1676037725
transform 1 0 25576 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1676037725
transform 1 0 23000 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1676037725
transform 1 0 25852 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1676037725
transform 1 0 26956 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform 1 0 26956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1676037725
transform 1 0 25208 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1676037725
transform 1 0 25024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1676037725
transform 1 0 25024 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1676037725
transform 1 0 24840 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1676037725
transform 1 0 26680 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1676037725
transform 1 0 25208 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1676037725
transform 1 0 26956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1676037725
transform 1 0 26404 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 24656 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1676037725
transform 1 0 26956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1676037725
transform 1 0 26956 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1676037725
transform 1 0 23644 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 19136 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 20700 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 21804 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 20976 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 19780 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 18768 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 12788 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 22724 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1676037725
transform 1 0 24748 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 25116 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1676037725
transform 1 0 17480 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 20516 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1676037725
transform 1 0 14904 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1676037725
transform 1 0 18768 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 22540 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 24104 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1676037725
transform 1 0 16192 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 14904 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1676037725
transform 1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 18308 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform 1 0 25944 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1676037725
transform 1 0 26956 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1676037725
transform 1 0 26496 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1676037725
transform 1 0 26220 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1676037725
transform 1 0 25116 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1676037725
transform 1 0 26956 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1676037725
transform 1 0 25208 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1676037725
transform 1 0 25208 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1676037725
transform 1 0 25208 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1676037725
transform 1 0 26864 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1075_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2760 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1076_
timestamp 1676037725
transform 1 0 1932 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1676037725
transform 1 0 2024 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1676037725
transform 1 0 2392 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1676037725
transform 1 0 2024 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1676037725
transform 1 0 3956 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1676037725
transform 1 0 3956 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1083_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1086_
timestamp 1676037725
transform -1 0 3772 0 -1 2176
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1087_
timestamp 1676037725
transform 1 0 1932 0 1 1088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1089_
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1676037725
transform 1 0 1656 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform -1 0 1840 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 1564 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 25300 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0390_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4692 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_in[0]
timestamp 1676037725
transform 1 0 2852 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net57
timestamp 1676037725
transform 1 0 1656 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 4968 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 2852 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0390_
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_io_in[0]
timestamp 1676037725
transform 1 0 2576 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net57
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 2576 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 1564 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0390_
timestamp 1676037725
transform 1 0 2576 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_io_in[0]
timestamp 1676037725
transform 1 0 2576 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net57
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.dcdel_capnode_notouch_
timestamp 1676037725
transform 1 0 1656 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1676037725
transform 1 0 2576 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout9
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1676037725
transform 1 0 11592 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout12
timestamp 1676037725
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1676037725
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1676037725
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1676037725
transform 1 0 9108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1676037725
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1676037725
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1676037725
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout23
timestamp 1676037725
transform 1 0 27140 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1676037725
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1676037725
transform 1 0 23736 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1676037725
transform 1 0 18584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1676037725
transform 1 0 9200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1676037725
transform 1 0 1748 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47
timestamp 1676037725
transform 1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1676037725
transform 1 0 13064 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_152 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1676037725
transform 1 0 15640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1676037725
transform 1 0 19780 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1676037725
transform 1 0 20516 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_8
timestamp 1676037725
transform 1 0 1840 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1676037725
transform 1 0 3772 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1676037725
transform 1 0 5612 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1676037725
transform 1 0 7820 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1676037725
transform 1 0 9384 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1676037725
transform 1 0 12144 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_140
timestamp 1676037725
transform 1 0 13984 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1676037725
transform 1 0 14720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1676037725
transform 1 0 21344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_263
timestamp 1676037725
transform 1 0 25300 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1676037725
transform 1 0 26312 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1676037725
transform 1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1676037725
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_173
timestamp 1676037725
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_217
timestamp 1676037725
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_139
timestamp 1676037725
transform 1 0 13892 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1676037725
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1676037725
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1676037725
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1676037725
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1676037725
transform 1 0 4324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_63
timestamp 1676037725
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_105
timestamp 1676037725
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1676037725
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_164
timestamp 1676037725
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1676037725
transform 1 0 17296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_227
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1676037725
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1676037725
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1676037725
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1676037725
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_195
timestamp 1676037725
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_255
timestamp 1676037725
transform 1 0 24564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1676037725
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_106
timestamp 1676037725
transform 1 0 10856 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1676037725
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_152
timestamp 1676037725
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_156
timestamp 1676037725
transform 1 0 15456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_181
timestamp 1676037725
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1676037725
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1676037725
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_291
timestamp 1676037725
transform 1 0 27876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1676037725
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1676037725
transform 1 0 4140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1676037725
transform 1 0 4508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1676037725
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_148
timestamp 1676037725
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_158
timestamp 1676037725
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_176
timestamp 1676037725
transform 1 0 17296 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1676037725
transform 1 0 18032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1676037725
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_45
timestamp 1676037725
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_57
timestamp 1676037725
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1676037725
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_157
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_171
timestamp 1676037725
transform 1 0 16836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1676037725
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1676037725
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_279
timestamp 1676037725
transform 1 0 26772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1676037725
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1676037725
transform 1 0 3036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1676037725
transform 1 0 3404 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1676037725
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_38
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1676037725
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1676037725
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_83
timestamp 1676037725
transform 1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1676037725
transform 1 0 9476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1676037725
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_143
timestamp 1676037725
transform 1 0 14260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_147
timestamp 1676037725
transform 1 0 14628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1676037725
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_212
timestamp 1676037725
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_232
timestamp 1676037725
transform 1 0 22448 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_240
timestamp 1676037725
transform 1 0 23184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 1676037725
transform 1 0 5796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1676037725
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_98
timestamp 1676037725
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_110
timestamp 1676037725
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1676037725
transform 1 0 15640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_204
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_226
timestamp 1676037725
transform 1 0 21896 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp 1676037725
transform 1 0 23368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 1676037725
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_274
timestamp 1676037725
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1676037725
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1676037725
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1676037725
transform 1 0 8188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1676037725
transform 1 0 9752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1676037725
transform 1 0 12788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1676037725
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_146
timestamp 1676037725
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1676037725
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1676037725
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_179
timestamp 1676037725
transform 1 0 17572 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp 1676037725
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_196
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_204
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1676037725
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1676037725
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1676037725
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_40
timestamp 1676037725
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1676037725
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_69
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1676037725
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_104
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_116
timestamp 1676037725
transform 1 0 11776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1676037725
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_171
timestamp 1676037725
transform 1 0 16836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1676037725
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_280
timestamp 1676037725
transform 1 0 26864 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1676037725
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1676037725
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_66
timestamp 1676037725
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_70
timestamp 1676037725
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_87
timestamp 1676037725
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_99
timestamp 1676037725
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1676037725
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_189
timestamp 1676037725
transform 1 0 18492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_197
timestamp 1676037725
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1676037725
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_231
timestamp 1676037725
transform 1 0 22356 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_251
timestamp 1676037725
transform 1 0 24196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_39
timestamp 1676037725
transform 1 0 4692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_48
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1676037725
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_73
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1676037725
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_94
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1676037725
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1676037725
transform 1 0 16652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1676037725
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1676037725
transform 1 0 28336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_24
timestamp 1676037725
transform 1 0 3312 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1676037725
transform 1 0 4048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1676037725
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1676037725
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1676037725
transform 1 0 7636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_75
timestamp 1676037725
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_88
timestamp 1676037725
transform 1 0 9200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1676037725
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_151
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1676037725
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_236
timestamp 1676037725
transform 1 0 22816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_240
timestamp 1676037725
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_257
timestamp 1676037725
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1676037725
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_19
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_37
timestamp 1676037725
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1676037725
transform 1 0 5520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_56
timestamp 1676037725
transform 1 0 6256 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1676037725
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1676037725
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_91
timestamp 1676037725
transform 1 0 9476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_104
timestamp 1676037725
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_128
timestamp 1676037725
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_224
timestamp 1676037725
transform 1 0 21712 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_231
timestamp 1676037725
transform 1 0 22356 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1676037725
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_46
timestamp 1676037725
transform 1 0 5336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 1676037725
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1676037725
transform 1 0 7912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1676037725
transform 1 0 8648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_92
timestamp 1676037725
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_96
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1676037725
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_235
timestamp 1676037725
transform 1 0 22724 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_257
timestamp 1676037725
transform 1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_290
timestamp 1676037725
transform 1 0 27784 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1676037725
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_44
timestamp 1676037725
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_117
timestamp 1676037725
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1676037725
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_211
timestamp 1676037725
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_223
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_231
timestamp 1676037725
transform 1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_242
timestamp 1676037725
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_262
timestamp 1676037725
transform 1 0 25208 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_286
timestamp 1676037725
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1676037725
transform 1 0 28520 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_64
timestamp 1676037725
transform 1 0 6992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_72
timestamp 1676037725
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_90
timestamp 1676037725
transform 1 0 9384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_139
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1676037725
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_290
timestamp 1676037725
transform 1 0 27784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1676037725
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1676037725
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1676037725
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1676037725
transform 1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_102
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1676037725
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 1676037725
transform 1 0 19872 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_228
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_65
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1676037725
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_145
timestamp 1676037725
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_186
timestamp 1676037725
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_190
timestamp 1676037725
transform 1 0 18584 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_195
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1676037725
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_40
timestamp 1676037725
transform 1 0 4784 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_48
timestamp 1676037725
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_56
timestamp 1676037725
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_67
timestamp 1676037725
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1676037725
transform 1 0 7636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1676037725
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1676037725
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1676037725
transform 1 0 10488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1676037725
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1676037725
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1676037725
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_168
timestamp 1676037725
transform 1 0 16560 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_184
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_232
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_240
timestamp 1676037725
transform 1 0 23184 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_272
timestamp 1676037725
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_292
timestamp 1676037725
transform 1 0 27968 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1676037725
transform 1 0 28520 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_30
timestamp 1676037725
transform 1 0 3864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_38
timestamp 1676037725
transform 1 0 4600 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1676037725
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_144
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1676037725
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_232
timestamp 1676037725
transform 1 0 22448 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_240
timestamp 1676037725
transform 1 0 23184 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1676037725
transform 1 0 23736 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_266
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1676037725
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_9
timestamp 1676037725
transform 1 0 1932 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1676037725
transform 1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_38
timestamp 1676037725
transform 1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1676037725
transform 1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_55
timestamp 1676037725
transform 1 0 6164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1676037725
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1676037725
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_173
timestamp 1676037725
transform 1 0 17020 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1676037725
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_203
timestamp 1676037725
transform 1 0 19780 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_268
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_280
timestamp 1676037725
transform 1 0 26864 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1676037725
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1676037725
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1676037725
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1676037725
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1676037725
transform 1 0 9016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1676037725
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_131
timestamp 1676037725
transform 1 0 13156 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_143
timestamp 1676037725
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_147
timestamp 1676037725
transform 1 0 14628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1676037725
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1676037725
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_202
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_252
timestamp 1676037725
transform 1 0 24288 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_260
timestamp 1676037725
transform 1 0 25024 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1676037725
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_36
timestamp 1676037725
transform 1 0 4416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_44
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1676037725
transform 1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1676037725
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_63
timestamp 1676037725
transform 1 0 6900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1676037725
transform 1 0 9752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_105
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1676037725
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_279
timestamp 1676037725
transform 1 0 26772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1676037725
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_12
timestamp 1676037725
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_67
timestamp 1676037725
transform 1 0 7268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_94
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_122
timestamp 1676037725
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_183
timestamp 1676037725
transform 1 0 17940 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_13
timestamp 1676037725
transform 1 0 2300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1676037725
transform 1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1676037725
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1676037725
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_66
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_94
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_100
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1676037725
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_220
timestamp 1676037725
transform 1 0 21344 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1676037725
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_279
timestamp 1676037725
transform 1 0 26772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1676037725
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_9
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1676037725
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1676037725
transform 1 0 3864 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1676037725
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_122
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_198
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1676037725
transform 1 0 19872 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_40
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1676037725
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1676037725
transform 1 0 6808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_92
timestamp 1676037725
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1676037725
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1676037725
transform 1 0 10672 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_126
timestamp 1676037725
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_149
timestamp 1676037725
transform 1 0 14812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_161
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_227
timestamp 1676037725
transform 1 0 21988 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_240
timestamp 1676037725
transform 1 0 23184 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1676037725
transform 1 0 26496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_280
timestamp 1676037725
transform 1 0 26864 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1676037725
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_19
timestamp 1676037725
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_31
timestamp 1676037725
transform 1 0 3956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1676037725
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_74
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_90
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1676037725
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_183
timestamp 1676037725
transform 1 0 17940 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_201
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_232
timestamp 1676037725
transform 1 0 22448 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_36
timestamp 1676037725
transform 1 0 4416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1676037725
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 1676037725
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1676037725
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_211
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1676037725
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1676037725
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_67
timestamp 1676037725
transform 1 0 7268 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_83
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_101
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1676037725
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_131
timestamp 1676037725
transform 1 0 13156 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1676037725
transform 1 0 19872 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_247
timestamp 1676037725
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_259
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_36
timestamp 1676037725
transform 1 0 4416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_45
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_55
timestamp 1676037725
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_64
timestamp 1676037725
transform 1 0 6992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_72
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_100
timestamp 1676037725
transform 1 0 10304 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_116
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1676037725
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1676037725
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp 1676037725
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_238
timestamp 1676037725
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_261
timestamp 1676037725
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_278
timestamp 1676037725
transform 1 0 26680 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_290
timestamp 1676037725
transform 1 0 27784 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_298
timestamp 1676037725
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1676037725
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_63
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_70
timestamp 1676037725
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_76
timestamp 1676037725
transform 1 0 8096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_92
timestamp 1676037725
transform 1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_122
timestamp 1676037725
transform 1 0 12328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_134
timestamp 1676037725
transform 1 0 13432 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_140
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_263
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_55
timestamp 1676037725
transform 1 0 6164 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_69
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1676037725
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_148
timestamp 1676037725
transform 1 0 14720 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_172
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1676037725
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_26
timestamp 1676037725
transform 1 0 3496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_36
timestamp 1676037725
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1676037725
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1676037725
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_67
timestamp 1676037725
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1676037725
transform 1 0 13616 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_155
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_185
timestamp 1676037725
transform 1 0 18124 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_256
timestamp 1676037725
transform 1 0 24656 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_49
timestamp 1676037725
transform 1 0 5612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_71
timestamp 1676037725
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_110
timestamp 1676037725
transform 1 0 11224 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_129
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1676037725
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_162
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1676037725
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_271
timestamp 1676037725
transform 1 0 26036 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_65
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_72
timestamp 1676037725
transform 1 0 7728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_84
timestamp 1676037725
transform 1 0 8832 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_92
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1676037725
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_144
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_156
timestamp 1676037725
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1676037725
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_243
timestamp 1676037725
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_263
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1676037725
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_52
timestamp 1676037725
transform 1 0 5888 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_64
timestamp 1676037725
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_76
timestamp 1676037725
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_93
timestamp 1676037725
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_99
timestamp 1676037725
transform 1 0 10212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_128
timestamp 1676037725
transform 1 0 12880 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_217
timestamp 1676037725
transform 1 0 21068 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_223
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_235
timestamp 1676037725
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_285
timestamp 1676037725
transform 1 0 27324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1676037725
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_8
timestamp 1676037725
transform 1 0 1840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_36
timestamp 1676037725
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_48
timestamp 1676037725
transform 1 0 5520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_64
timestamp 1676037725
transform 1 0 6992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_68
timestamp 1676037725
transform 1 0 7360 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_74
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_86
timestamp 1676037725
transform 1 0 9016 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_92
timestamp 1676037725
transform 1 0 9568 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1676037725
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_122
timestamp 1676037725
transform 1 0 12328 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_134
timestamp 1676037725
transform 1 0 13432 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1676037725
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_14
timestamp 1676037725
transform 1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_48
timestamp 1676037725
transform 1 0 5520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_56
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_74
timestamp 1676037725
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_103
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_115
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_128
timestamp 1676037725
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_170
timestamp 1676037725
transform 1 0 16744 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_215
timestamp 1676037725
transform 1 0 20884 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_232
timestamp 1676037725
transform 1 0 22448 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1676037725
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_12
timestamp 1676037725
transform 1 0 2208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_25
timestamp 1676037725
transform 1 0 3404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_32
timestamp 1676037725
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_45
timestamp 1676037725
transform 1 0 5244 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1676037725
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1676037725
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1676037725
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_132
timestamp 1676037725
transform 1 0 13248 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1676037725
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_176
timestamp 1676037725
transform 1 0 17296 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_188
timestamp 1676037725
transform 1 0 18400 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_200
timestamp 1676037725
transform 1 0 19504 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_212
timestamp 1676037725
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1676037725
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_40
timestamp 1676037725
transform 1 0 4784 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_48
timestamp 1676037725
transform 1 0 5520 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_57
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1676037725
transform 1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1676037725
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_96
timestamp 1676037725
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_108
timestamp 1676037725
transform 1 0 11040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_122
timestamp 1676037725
transform 1 0 12328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_126
timestamp 1676037725
transform 1 0 12696 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1676037725
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_261
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_272
timestamp 1676037725
transform 1 0 26128 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_280
timestamp 1676037725
transform 1 0 26864 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1676037725
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_10
timestamp 1676037725
transform 1 0 2024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_31
timestamp 1676037725
transform 1 0 3956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1676037725
transform 1 0 5152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_66
timestamp 1676037725
transform 1 0 7176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_87
timestamp 1676037725
transform 1 0 9108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_99
timestamp 1676037725
transform 1 0 10212 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1676037725
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_124
timestamp 1676037725
transform 1 0 12512 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_130
timestamp 1676037725
transform 1 0 13064 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_136
timestamp 1676037725
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1676037725
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_203
timestamp 1676037725
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1676037725
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1676037725
transform 1 0 5428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_54
timestamp 1676037725
transform 1 0 6072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_58
timestamp 1676037725
transform 1 0 6440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_64
timestamp 1676037725
transform 1 0 6992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_71
timestamp 1676037725
transform 1 0 7636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1676037725
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1676037725
transform 1 0 9476 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_101
timestamp 1676037725
transform 1 0 10396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_113
timestamp 1676037725
transform 1 0 11500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1676037725
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1676037725
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_161
timestamp 1676037725
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_180
timestamp 1676037725
transform 1 0 17664 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1676037725
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_241
timestamp 1676037725
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_282
timestamp 1676037725
transform 1 0 27048 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1676037725
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_298
timestamp 1676037725
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_14
timestamp 1676037725
transform 1 0 2392 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_35
timestamp 1676037725
transform 1 0 4324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1676037725
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_64
timestamp 1676037725
transform 1 0 6992 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_71
timestamp 1676037725
transform 1 0 7636 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_78
timestamp 1676037725
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_90
timestamp 1676037725
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1676037725
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_124
timestamp 1676037725
transform 1 0 12512 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_130
timestamp 1676037725
transform 1 0 13064 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1676037725
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_145
timestamp 1676037725
transform 1 0 14444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_157
timestamp 1676037725
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1676037725
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_188
timestamp 1676037725
transform 1 0 18400 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_212
timestamp 1676037725
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_254
timestamp 1676037725
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_266
timestamp 1676037725
transform 1 0 25576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1676037725
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_35
timestamp 1676037725
transform 1 0 4324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_59
timestamp 1676037725
transform 1 0 6532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_73
timestamp 1676037725
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1676037725
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_90
timestamp 1676037725
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_98
timestamp 1676037725
transform 1 0 10120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_104
timestamp 1676037725
transform 1 0 10672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_113
timestamp 1676037725
transform 1 0 11500 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_120
timestamp 1676037725
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1676037725
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_146
timestamp 1676037725
transform 1 0 14536 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_158
timestamp 1676037725
transform 1 0 15640 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_170
timestamp 1676037725
transform 1 0 16744 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_182
timestamp 1676037725
transform 1 0 17848 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_229
timestamp 1676037725
transform 1 0 22172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1676037725
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1676037725
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1676037725
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_12
timestamp 1676037725
transform 1 0 2208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_36
timestamp 1676037725
transform 1 0 4416 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_45
timestamp 1676037725
transform 1 0 5244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1676037725
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_64
timestamp 1676037725
transform 1 0 6992 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_77
timestamp 1676037725
transform 1 0 8188 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_86
timestamp 1676037725
transform 1 0 9016 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_94
timestamp 1676037725
transform 1 0 9752 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_106
timestamp 1676037725
transform 1 0 10856 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_132
timestamp 1676037725
transform 1 0 13248 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_144
timestamp 1676037725
transform 1 0 14352 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_9
timestamp 1676037725
transform 1 0 1932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1676037725
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_47
timestamp 1676037725
transform 1 0 5428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_56
timestamp 1676037725
transform 1 0 6256 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1676037725
transform 1 0 6992 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_71
timestamp 1676037725
transform 1 0 7636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1676037725
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_90
timestamp 1676037725
transform 1 0 9384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_104
timestamp 1676037725
transform 1 0 10672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_112
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_118
timestamp 1676037725
transform 1 0 11960 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_127
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_148
timestamp 1676037725
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_160
timestamp 1676037725
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_172
timestamp 1676037725
transform 1 0 16928 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_184
timestamp 1676037725
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1676037725
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_12
timestamp 1676037725
transform 1 0 2208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_36
timestamp 1676037725
transform 1 0 4416 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_44
timestamp 1676037725
transform 1 0 5152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_68
timestamp 1676037725
transform 1 0 7360 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_72
timestamp 1676037725
transform 1 0 7728 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_76
timestamp 1676037725
transform 1 0 8096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_83
timestamp 1676037725
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_90
timestamp 1676037725
transform 1 0 9384 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_97
timestamp 1676037725
transform 1 0 10028 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_103
timestamp 1676037725
transform 1 0 10580 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1676037725
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_127
timestamp 1676037725
transform 1 0 12788 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_138
timestamp 1676037725
transform 1 0 13800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_147
timestamp 1676037725
transform 1 0 14628 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_155
timestamp 1676037725
transform 1 0 15364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1676037725
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_51
timestamp 1676037725
transform 1 0 5796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_60
timestamp 1676037725
transform 1 0 6624 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_68
timestamp 1676037725
transform 1 0 7360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_74
timestamp 1676037725
transform 1 0 7912 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1676037725
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_90
timestamp 1676037725
transform 1 0 9384 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_101
timestamp 1676037725
transform 1 0 10396 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_110
timestamp 1676037725
transform 1 0 11224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_118
timestamp 1676037725
transform 1 0 11960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_129
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_154
timestamp 1676037725
transform 1 0 15272 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_163
timestamp 1676037725
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_175
timestamp 1676037725
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1676037725
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1676037725
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_64
timestamp 1676037725
transform 1 0 6992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_73
timestamp 1676037725
transform 1 0 7820 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_88
timestamp 1676037725
transform 1 0 9200 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_127
timestamp 1676037725
transform 1 0 12788 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1676037725
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1676037725
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1676037725
transform 1 0 15272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1676037725
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1676037725
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_38
timestamp 1676037725
transform 1 0 4600 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_62
timestamp 1676037725
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_66
timestamp 1676037725
transform 1 0 7176 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_72
timestamp 1676037725
transform 1 0 7728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_76
timestamp 1676037725
transform 1 0 8096 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_94
timestamp 1676037725
transform 1 0 9752 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_103
timestamp 1676037725
transform 1 0 10580 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_112
timestamp 1676037725
transform 1 0 11408 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_129
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1676037725
transform 1 0 15272 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_162
timestamp 1676037725
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_174
timestamp 1676037725
transform 1 0 17112 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 1676037725
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_297
timestamp 1676037725
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_12
timestamp 1676037725
transform 1 0 2208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_36
timestamp 1676037725
transform 1 0 4416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_70
timestamp 1676037725
transform 1 0 7544 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_79
timestamp 1676037725
transform 1 0 8372 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_88
timestamp 1676037725
transform 1 0 9200 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_101
timestamp 1676037725
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_120
timestamp 1676037725
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_128
timestamp 1676037725
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_133
timestamp 1676037725
transform 1 0 13340 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_142
timestamp 1676037725
transform 1 0 14168 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_151
timestamp 1676037725
transform 1 0 14996 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1676037725
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1676037725
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_39
timestamp 1676037725
transform 1 0 4692 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_47
timestamp 1676037725
transform 1 0 5428 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_62
timestamp 1676037725
transform 1 0 6808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_69
timestamp 1676037725
transform 1 0 7452 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1676037725
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_90
timestamp 1676037725
transform 1 0 9384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_94
timestamp 1676037725
transform 1 0 9752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_100
timestamp 1676037725
transform 1 0 10304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_118
timestamp 1676037725
transform 1 0 11960 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_126
timestamp 1676037725
transform 1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_146
timestamp 1676037725
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1676037725
transform 1 0 15824 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_167
timestamp 1676037725
transform 1 0 16468 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_179
timestamp 1676037725
transform 1 0 17572 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_191
timestamp 1676037725
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_297
timestamp 1676037725
transform 1 0 28428 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_25
timestamp 1676037725
transform 1 0 3404 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_29
timestamp 1676037725
transform 1 0 3772 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_36
timestamp 1676037725
transform 1 0 4416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1676037725
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1676037725
transform 1 0 6808 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_82
timestamp 1676037725
transform 1 0 8648 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1676037725
transform 1 0 8924 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 1676037725
transform 1 0 9568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1676037725
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_103
timestamp 1676037725
transform 1 0 10580 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 1676037725
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1676037725
transform 1 0 11960 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_132
timestamp 1676037725
transform 1 0 13248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1676037725
transform 1 0 14076 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_146
timestamp 1676037725
transform 1 0 14536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1676037725
transform 1 0 15180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1676037725
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_197
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1676037725
transform 1 0 20332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1676037725
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_253
timestamp 1676037725
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_265
timestamp 1676037725
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1676037725
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 28888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 28888 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[0\].cap
timestamp 1676037725
transform 1 0 16192 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[0\].cap_39 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[1\].cap_46
timestamp 1676037725
transform 1 0 6532 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[1\].cap
timestamp 1676037725
transform 1 0 4416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[2\].cap_47
timestamp 1676037725
transform 1 0 7820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[2\].cap
timestamp 1676037725
transform 1 0 8004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[3\].cap
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[3\].cap_48
timestamp 1676037725
transform 1 0 13064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[4\].cap
timestamp 1676037725
transform 1 0 15548 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[4\].cap_49
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[5\].cap_50
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[5\].cap
timestamp 1676037725
transform 1 0 10396 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[6\].cap_51
timestamp 1676037725
transform 1 0 7176 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[6\].cap
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[7\].cap
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[7\].cap_52
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[8\].cap
timestamp 1676037725
transform 1 0 12328 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[8\].cap_53
timestamp 1676037725
transform 1 0 7176 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[9\].cap_54
timestamp 1676037725
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[9\].cap
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[10\].cap
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[10\].cap_40
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[11\].cap_41
timestamp 1676037725
transform 1 0 9108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[11\].cap
timestamp 1676037725
transform 1 0 3772 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[12\].cap_42
timestamp 1676037725
transform 1 0 6532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[12\].cap
timestamp 1676037725
transform 1 0 9752 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[13\].cap
timestamp 1676037725
transform 1 0 14904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[13\].cap_43
timestamp 1676037725
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[14\].cap_44
timestamp 1676037725
transform 1 0 9936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[14\].cap
timestamp 1676037725
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  temp1.capload\[15\].cap_45
timestamp 1676037725
transform 1 0 12972 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  temp1.capload\[15\].cap
timestamp 1676037725
transform 1 0 14904 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 9844 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 7728 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 11040 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 10212 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 13156 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 12328 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 13156 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 12328 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 12328 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 13156 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 13156 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 11500 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 6164 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 8188 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 7360 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 8740 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 6532 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 8740 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 5612 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 7912 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1676037725
transform 1 0 7268 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1676037725
transform 1 0 4784 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1676037725
transform 1 0 5520 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1676037725
transform 1 0 4784 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1676037725
transform 1 0 7084 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 11500 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1676037725
transform 1 0 15640 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1676037725
transform 1 0 10672 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1676037725
transform 1 0 13156 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1676037725
transform 1 0 11776 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1676037725
transform 1 0 12512 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1676037725
transform 1 0 9292 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1676037725
transform 1 0 10672 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1676037725
transform 1 0 14812 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1676037725
transform 1 0 10120 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1676037725
transform 1 0 10948 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1676037725
transform 1 0 12328 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1676037725
transform 1 0 9936 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1676037725
transform 1 0 14168 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1676037725
transform 1 0 9844 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1676037725
transform 1 0 14812 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1676037725
transform 1 0 9936 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1676037725
transform 1 0 14536 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1676037725
transform 1 0 10672 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1676037725
transform 1 0 10764 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1676037725
transform 1 0 11684 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1676037725
transform 1 0 15640 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1676037725
transform 1 0 9936 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd_56
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1676037725
transform 1 0 13984 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  temp1.dac.vdac_single.einvp_batch\[0\].vref
timestamp 1676037725
transform 1 0 18032 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  temp1.dac.vdac_single.einvp_batch\[0\].vref_55
timestamp 1676037725
transform 1 0 18124 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  temp1.dcdc
timestamp 1676037725
transform 1 0 3956 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  temp1.inv1_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_2
timestamp 1676037725
transform 1 0 2760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_3
timestamp 1676037725
transform 1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  temp1.inv2_4
timestamp 1676037725
transform 1 0 9108 0 1 27200
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 1640 400 1760 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 3680 400 3800 0 FreeSans 480 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 0 5720 400 5840 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal3 s 0 7760 400 7880 0 FreeSans 480 0 0 0 io_in[3]
port 3 nsew signal input
flabel metal3 s 0 9800 400 9920 0 FreeSans 480 0 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 0 11840 400 11960 0 FreeSans 480 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal3 s 0 13880 400 14000 0 FreeSans 480 0 0 0 io_in[6]
port 6 nsew signal input
flabel metal3 s 0 15920 400 16040 0 FreeSans 480 0 0 0 io_in[7]
port 7 nsew signal input
flabel metal3 s 0 17960 400 18080 0 FreeSans 480 0 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal3 s 0 20000 400 20120 0 FreeSans 480 0 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal3 s 0 22040 400 22160 0 FreeSans 480 0 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal3 s 0 24080 400 24200 0 FreeSans 480 0 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal3 s 0 26120 400 26240 0 FreeSans 480 0 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal3 s 0 28160 400 28280 0 FreeSans 480 0 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal3 s 0 30200 400 30320 0 FreeSans 480 0 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal3 s 0 32240 400 32360 0 FreeSans 480 0 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 4417 1040 4737 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 11363 1040 11683 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 18309 1040 18629 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 25255 1040 25575 32688 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7890 1040 8210 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 14836 1040 15156 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 21782 1040 22102 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 28728 1040 29048 32688 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 14996 32096 14996 32096 0 vccd1
rlabel via1 15076 32640 15076 32640 0 vssd1
rlabel metal1 3951 26962 3951 26962 0 _0000_
rlabel metal1 4002 27472 4002 27472 0 _0001_
rlabel metal2 4278 25500 4278 25500 0 _0002_
rlabel metal1 2336 25874 2336 25874 0 _0003_
rlabel metal2 4278 27166 4278 27166 0 _0004_
rlabel metal2 3450 29002 3450 29002 0 _0005_
rlabel metal2 4370 29274 4370 29274 0 _0006_
rlabel metal1 8050 1190 8050 1190 0 _0007_
rlabel metal2 2530 12784 2530 12784 0 _0008_
rlabel metal2 1886 9316 1886 9316 0 _0009_
rlabel metal1 1962 2346 1962 2346 0 _0010_
rlabel metal3 14513 25228 14513 25228 0 _0011_
rlabel via1 2249 1258 2249 1258 0 _0012_
rlabel metal1 12926 19210 12926 19210 0 _0013_
rlabel metal1 1824 3434 1824 3434 0 _0014_
rlabel metal1 1784 4590 1784 4590 0 _0015_
rlabel metal1 3496 19482 3496 19482 0 _0016_
rlabel metal1 2162 16966 2162 16966 0 _0017_
rlabel metal2 2714 6817 2714 6817 0 _0018_
rlabel metal1 3588 5882 3588 5882 0 _0019_
rlabel metal1 11914 16626 11914 16626 0 _0020_
rlabel metal1 6440 20026 6440 20026 0 _0021_
rlabel metal1 6532 17306 6532 17306 0 _0022_
rlabel metal2 7728 18564 7728 18564 0 _0023_
rlabel metal2 14766 24276 14766 24276 0 _0024_
rlabel metal1 11546 23698 11546 23698 0 _0025_
rlabel metal1 2254 24072 2254 24072 0 _0026_
rlabel metal1 4830 29478 4830 29478 0 _0027_
rlabel metal1 9798 29172 9798 29172 0 _0028_
rlabel metal2 2438 26724 2438 26724 0 _0029_
rlabel metal1 12834 24208 12834 24208 0 _0030_
rlabel metal2 8326 24718 8326 24718 0 _0031_
rlabel metal1 8602 20026 8602 20026 0 _0032_
rlabel metal1 5658 19890 5658 19890 0 _0033_
rlabel metal2 2806 16796 2806 16796 0 _0034_
rlabel metal1 14674 17646 14674 17646 0 _0035_
rlabel metal1 1978 30294 1978 30294 0 _0036_
rlabel metal1 9936 20230 9936 20230 0 _0037_
rlabel metal1 4186 18904 4186 18904 0 _0038_
rlabel metal1 11040 19346 11040 19346 0 _0039_
rlabel metal1 8004 18666 8004 18666 0 _0040_
rlabel metal1 7774 15028 7774 15028 0 _0041_
rlabel metal1 9108 14382 9108 14382 0 _0042_
rlabel metal1 7130 13940 7130 13940 0 _0043_
rlabel metal1 7038 13770 7038 13770 0 _0044_
rlabel metal2 2438 14348 2438 14348 0 _0045_
rlabel metal1 5244 13838 5244 13838 0 _0046_
rlabel metal1 8766 13906 8766 13906 0 _0047_
rlabel metal1 13570 12818 13570 12818 0 _0048_
rlabel metal2 17250 19346 17250 19346 0 _0049_
rlabel metal1 17066 6800 17066 6800 0 _0050_
rlabel metal1 21528 15402 21528 15402 0 _0051_
rlabel metal1 14904 13430 14904 13430 0 _0052_
rlabel metal1 12834 12682 12834 12682 0 _0053_
rlabel metal1 1886 29172 1886 29172 0 _0054_
rlabel metal1 11776 12206 11776 12206 0 _0055_
rlabel metal2 9246 10336 9246 10336 0 _0056_
rlabel metal1 11546 13226 11546 13226 0 _0057_
rlabel metal1 18224 17238 18224 17238 0 _0058_
rlabel metal1 18676 7990 18676 7990 0 _0059_
rlabel metal1 13800 8466 13800 8466 0 _0060_
rlabel metal3 17825 16660 17825 16660 0 _0061_
rlabel metal1 19626 8262 19626 8262 0 _0062_
rlabel metal2 20930 16626 20930 16626 0 _0063_
rlabel metal1 20976 9554 20976 9554 0 _0064_
rlabel metal1 24242 1972 24242 1972 0 _0065_
rlabel metal1 15870 13226 15870 13226 0 _0066_
rlabel metal1 17296 14994 17296 14994 0 _0067_
rlabel metal1 18538 14858 18538 14858 0 _0068_
rlabel metal1 19550 11662 19550 11662 0 _0069_
rlabel metal2 19734 10234 19734 10234 0 _0070_
rlabel metal1 13754 9384 13754 9384 0 _0071_
rlabel via1 19920 4590 19920 4590 0 _0072_
rlabel metal1 17434 12172 17434 12172 0 _0073_
rlabel metal1 16392 13974 16392 13974 0 _0074_
rlabel metal1 18906 13872 18906 13872 0 _0075_
rlabel metal1 25875 9554 25875 9554 0 _0076_
rlabel metal2 20700 9860 20700 9860 0 _0077_
rlabel metal1 19826 4726 19826 4726 0 _0078_
rlabel metal1 20056 16150 20056 16150 0 _0079_
rlabel via1 20666 6766 20666 6766 0 _0080_
rlabel metal1 22180 18326 22180 18326 0 _0081_
rlabel metal1 21965 14246 21965 14246 0 _0082_
rlabel metal1 13478 12614 13478 12614 0 _0083_
rlabel metal1 22126 1428 22126 1428 0 _0084_
rlabel metal1 25392 14382 25392 14382 0 _0085_
rlabel metal2 22678 11322 22678 11322 0 _0086_
rlabel metal1 19550 9044 19550 9044 0 _0087_
rlabel metal1 14168 12750 14168 12750 0 _0088_
rlabel metal2 12696 13702 12696 13702 0 _0089_
rlabel metal1 15410 12954 15410 12954 0 _0090_
rlabel metal1 20378 7480 20378 7480 0 _0091_
rlabel metal1 17066 16592 17066 16592 0 _0092_
rlabel metal1 18883 18258 18883 18258 0 _0093_
rlabel metal1 11776 11322 11776 11322 0 _0094_
rlabel via1 21116 1938 21116 1938 0 _0095_
rlabel metal1 20792 7854 20792 7854 0 _0096_
rlabel metal2 22310 8143 22310 8143 0 _0097_
rlabel metal1 11546 9996 11546 9996 0 _0098_
rlabel metal1 16054 15470 16054 15470 0 _0099_
rlabel metal1 20470 18700 20470 18700 0 _0100_
rlabel metal1 20424 7378 20424 7378 0 _0101_
rlabel metal1 14260 7786 14260 7786 0 _0102_
rlabel metal2 17710 16762 17710 16762 0 _0103_
rlabel metal3 18147 15300 18147 15300 0 _0104_
rlabel metal1 21298 12240 21298 12240 0 _0105_
rlabel metal1 13363 6766 13363 6766 0 _0106_
rlabel metal1 17112 11118 17112 11118 0 _0107_
rlabel metal1 16614 15130 16614 15130 0 _0108_
rlabel metal1 23140 7854 23140 7854 0 _0109_
rlabel metal2 10902 15793 10902 15793 0 _0110_
rlabel metal1 21436 10710 21436 10710 0 _0111_
rlabel metal2 15042 7021 15042 7021 0 _0112_
rlabel metal1 14398 6970 14398 6970 0 _0113_
rlabel metal1 17434 12614 17434 12614 0 _0114_
rlabel via1 16148 12818 16148 12818 0 _0115_
rlabel metal1 12328 5270 12328 5270 0 _0116_
rlabel metal2 18538 9044 18538 9044 0 _0117_
rlabel metal2 13570 6086 13570 6086 0 _0118_
rlabel metal2 14214 6698 14214 6698 0 _0119_
rlabel metal2 14812 2380 14812 2380 0 _0120_
rlabel metal1 20930 1904 20930 1904 0 _0121_
rlabel via1 24127 14994 24127 14994 0 _0122_
rlabel metal3 17687 15436 17687 15436 0 _0123_
rlabel metal1 15456 5882 15456 5882 0 _0124_
rlabel metal2 14398 7038 14398 7038 0 _0125_
rlabel metal2 10534 14637 10534 14637 0 _0126_
rlabel metal2 8602 12070 8602 12070 0 _0127_
rlabel metal2 9614 13872 9614 13872 0 _0128_
rlabel metal2 16146 7378 16146 7378 0 _0129_
rlabel metal1 15594 5202 15594 5202 0 _0130_
rlabel metal1 21068 1190 21068 1190 0 _0131_
rlabel metal1 15410 5032 15410 5032 0 _0132_
rlabel metal1 18262 8874 18262 8874 0 _0133_
rlabel metal1 15824 5134 15824 5134 0 _0134_
rlabel metal1 12788 2414 12788 2414 0 _0135_
rlabel metal1 13754 2618 13754 2618 0 _0136_
rlabel metal1 15410 5338 15410 5338 0 _0137_
rlabel metal2 17158 14586 17158 14586 0 _0138_
rlabel metal2 21114 17408 21114 17408 0 _0139_
rlabel metal2 20838 17816 20838 17816 0 _0140_
rlabel metal2 22402 15946 22402 15946 0 _0141_
rlabel metal1 20930 16660 20930 16660 0 _0142_
rlabel metal1 23736 12954 23736 12954 0 _0143_
rlabel metal1 22632 12614 22632 12614 0 _0144_
rlabel metal1 17020 12410 17020 12410 0 _0145_
rlabel via1 13662 8245 13662 8245 0 _0146_
rlabel metal1 9798 7446 9798 7446 0 _0147_
rlabel metal1 5704 14382 5704 14382 0 _0148_
rlabel metal1 4646 9452 4646 9452 0 _0149_
rlabel metal1 23276 13430 23276 13430 0 _0150_
rlabel metal2 23690 13600 23690 13600 0 _0151_
rlabel metal1 23644 12410 23644 12410 0 _0152_
rlabel metal1 19826 12818 19826 12818 0 _0153_
rlabel metal1 24426 10778 24426 10778 0 _0154_
rlabel metal1 23828 12750 23828 12750 0 _0155_
rlabel metal1 23506 6426 23506 6426 0 _0156_
rlabel metal1 19780 12614 19780 12614 0 _0157_
rlabel metal1 17250 15674 17250 15674 0 _0158_
rlabel metal1 16698 13498 16698 13498 0 _0159_
rlabel metal2 16790 17578 16790 17578 0 _0160_
rlabel metal1 18722 12750 18722 12750 0 _0161_
rlabel metal2 21482 16660 21482 16660 0 _0162_
rlabel metal2 20102 18564 20102 18564 0 _0163_
rlabel metal1 20240 18938 20240 18938 0 _0164_
rlabel metal2 19458 14569 19458 14569 0 _0165_
rlabel metal3 18216 11220 18216 11220 0 _0166_
rlabel metal1 14352 3706 14352 3706 0 _0167_
rlabel metal1 17388 8602 17388 8602 0 _0168_
rlabel metal2 19458 10948 19458 10948 0 _0169_
rlabel metal1 17664 9010 17664 9010 0 _0170_
rlabel metal1 18952 2414 18952 2414 0 _0171_
rlabel metal1 18308 2618 18308 2618 0 _0172_
rlabel metal1 16974 1190 16974 1190 0 _0173_
rlabel metal1 19872 1190 19872 1190 0 _0174_
rlabel metal1 18538 3094 18538 3094 0 _0175_
rlabel metal2 16238 10030 16238 10030 0 _0176_
rlabel metal1 9292 10778 9292 10778 0 _0177_
rlabel metal1 6716 12614 6716 12614 0 _0178_
rlabel metal1 14904 4726 14904 4726 0 _0179_
rlabel metal1 14812 9078 14812 9078 0 _0180_
rlabel metal1 15456 14042 15456 14042 0 _0181_
rlabel metal1 14996 8806 14996 8806 0 _0182_
rlabel metal1 17664 13498 17664 13498 0 _0183_
rlabel metal1 17894 12954 17894 12954 0 _0184_
rlabel metal3 17273 12988 17273 12988 0 _0185_
rlabel metal1 15778 11288 15778 11288 0 _0186_
rlabel metal1 18078 13923 18078 13923 0 _0187_
rlabel metal2 19458 12716 19458 12716 0 _0188_
rlabel metal1 18216 13770 18216 13770 0 _0189_
rlabel metal1 17480 13702 17480 13702 0 _0190_
rlabel metal2 13938 13061 13938 13061 0 _0191_
rlabel metal1 13846 7242 13846 7242 0 _0192_
rlabel metal1 16790 10438 16790 10438 0 _0193_
rlabel metal1 15134 10778 15134 10778 0 _0194_
rlabel metal2 18262 10676 18262 10676 0 _0195_
rlabel metal1 17158 9146 17158 9146 0 _0196_
rlabel metal1 16928 11050 16928 11050 0 _0197_
rlabel metal1 22678 5882 22678 5882 0 _0198_
rlabel metal1 23322 8058 23322 8058 0 _0199_
rlabel via2 22770 9571 22770 9571 0 _0200_
rlabel metal1 22862 9418 22862 9418 0 _0201_
rlabel metal1 22632 9486 22632 9486 0 _0202_
rlabel metal1 21206 5814 21206 5814 0 _0203_
rlabel metal2 17802 9826 17802 9826 0 _0204_
rlabel metal1 18308 10234 18308 10234 0 _0205_
rlabel metal1 7958 13906 7958 13906 0 _0206_
rlabel viali 6862 12886 6862 12886 0 _0207_
rlabel metal1 19596 14586 19596 14586 0 _0208_
rlabel metal2 17802 15232 17802 15232 0 _0209_
rlabel metal1 17894 14518 17894 14518 0 _0210_
rlabel metal1 17250 14246 17250 14246 0 _0211_
rlabel metal2 18906 6902 18906 6902 0 _0212_
rlabel metal2 20378 6358 20378 6358 0 _0213_
rlabel metal1 19504 8058 19504 8058 0 _0214_
rlabel metal1 15962 7208 15962 7208 0 _0215_
rlabel metal1 4876 18326 4876 18326 0 _0216_
rlabel metal1 8924 15878 8924 15878 0 _0217_
rlabel metal1 15778 7446 15778 7446 0 _0218_
rlabel metal1 15732 1530 15732 1530 0 _0219_
rlabel metal1 14398 1462 14398 1462 0 _0220_
rlabel metal2 14582 1632 14582 1632 0 _0221_
rlabel metal1 15226 1326 15226 1326 0 _0222_
rlabel metal1 16100 7514 16100 7514 0 _0223_
rlabel via2 15686 12835 15686 12835 0 _0224_
rlabel metal1 15916 9418 15916 9418 0 _0225_
rlabel metal1 16146 6970 16146 6970 0 _0226_
rlabel metal1 13340 7990 13340 7990 0 _0227_
rlabel metal1 22678 10642 22678 10642 0 _0228_
rlabel metal2 23828 16524 23828 16524 0 _0229_
rlabel metal2 22402 9044 22402 9044 0 _0230_
rlabel metal2 22218 10761 22218 10761 0 _0231_
rlabel metal1 16284 9554 16284 9554 0 _0232_
rlabel metal2 15226 9418 15226 9418 0 _0233_
rlabel metal1 8096 12682 8096 12682 0 _0234_
rlabel metal1 8234 12750 8234 12750 0 _0235_
rlabel metal2 7130 11356 7130 11356 0 _0236_
rlabel metal1 6578 9010 6578 9010 0 _0237_
rlabel metal2 6762 9418 6762 9418 0 _0238_
rlabel metal1 19596 15878 19596 15878 0 _0239_
rlabel metal1 22218 10030 22218 10030 0 _0240_
rlabel metal1 20654 1836 20654 1836 0 _0241_
rlabel metal1 21574 10234 21574 10234 0 _0242_
rlabel metal2 23598 16932 23598 16932 0 _0243_
rlabel metal1 21804 10098 21804 10098 0 _0244_
rlabel metal1 26634 14042 26634 14042 0 _0245_
rlabel metal1 25668 9690 25668 9690 0 _0246_
rlabel metal1 16330 10098 16330 10098 0 _0247_
rlabel metal1 18032 18258 18032 18258 0 _0248_
rlabel metal3 16859 18020 16859 18020 0 _0249_
rlabel metal1 16330 6324 16330 6324 0 _0250_
rlabel metal1 15732 6426 15732 6426 0 _0251_
rlabel metal2 15318 6868 15318 6868 0 _0252_
rlabel metal2 17526 7956 17526 7956 0 _0253_
rlabel metal2 12558 6018 12558 6018 0 _0254_
rlabel metal2 12190 7582 12190 7582 0 _0255_
rlabel metal1 16008 8602 16008 8602 0 _0256_
rlabel metal2 8418 10370 8418 10370 0 _0257_
rlabel metal1 8142 9418 8142 9418 0 _0258_
rlabel metal1 8556 10710 8556 10710 0 _0259_
rlabel metal1 8924 10574 8924 10574 0 _0260_
rlabel metal1 6946 8908 6946 8908 0 _0261_
rlabel metal1 6210 7854 6210 7854 0 _0262_
rlabel metal1 6118 9146 6118 9146 0 _0263_
rlabel metal1 7222 9146 7222 9146 0 _0264_
rlabel metal1 7820 12954 7820 12954 0 _0265_
rlabel metal1 7130 12614 7130 12614 0 _0266_
rlabel metal1 6026 7378 6026 7378 0 _0267_
rlabel metal1 5474 6630 5474 6630 0 _0268_
rlabel via1 4830 7174 4830 7174 0 _0269_
rlabel metal1 6624 8466 6624 8466 0 _0270_
rlabel metal1 5520 6426 5520 6426 0 _0271_
rlabel metal2 5566 6970 5566 6970 0 _0272_
rlabel metal1 5704 8466 5704 8466 0 _0273_
rlabel metal2 5934 7446 5934 7446 0 _0274_
rlabel metal2 5290 9231 5290 9231 0 _0275_
rlabel metal1 4508 9146 4508 9146 0 _0276_
rlabel metal1 4094 10234 4094 10234 0 _0277_
rlabel metal2 3542 10642 3542 10642 0 _0278_
rlabel metal1 6762 12240 6762 12240 0 _0279_
rlabel metal1 4738 13362 4738 13362 0 _0280_
rlabel metal1 5888 10438 5888 10438 0 _0281_
rlabel metal1 5244 8874 5244 8874 0 _0282_
rlabel metal1 5014 9622 5014 9622 0 _0283_
rlabel metal1 5428 8806 5428 8806 0 _0284_
rlabel metal1 4692 7854 4692 7854 0 _0285_
rlabel metal1 4876 8058 4876 8058 0 _0286_
rlabel metal1 6118 11152 6118 11152 0 _0287_
rlabel metal2 5290 11492 5290 11492 0 _0288_
rlabel metal1 4140 11526 4140 11526 0 _0289_
rlabel metal2 5934 11764 5934 11764 0 _0290_
rlabel metal1 5290 12376 5290 12376 0 _0291_
rlabel metal1 5704 13294 5704 13294 0 _0292_
rlabel metal2 6946 12274 6946 12274 0 _0293_
rlabel metal1 7452 13430 7452 13430 0 _0294_
rlabel metal2 7682 16082 7682 16082 0 _0295_
rlabel metal1 1794 15436 1794 15436 0 _0296_
rlabel metal1 2369 15606 2369 15606 0 _0297_
rlabel metal1 7268 17850 7268 17850 0 _0298_
rlabel metal2 14490 16864 14490 16864 0 _0299_
rlabel metal1 8556 18938 8556 18938 0 _0300_
rlabel metal1 3266 17850 3266 17850 0 _0301_
rlabel metal2 5290 21624 5290 21624 0 _0302_
rlabel metal2 6762 21148 6762 21148 0 _0303_
rlabel metal1 5474 21998 5474 21998 0 _0304_
rlabel metal2 4370 20230 4370 20230 0 _0305_
rlabel metal2 2346 21828 2346 21828 0 _0306_
rlabel metal1 6256 21930 6256 21930 0 _0307_
rlabel metal2 8878 26078 8878 26078 0 _0308_
rlabel metal1 4324 13158 4324 13158 0 _0309_
rlabel metal1 5152 12614 5152 12614 0 _0310_
rlabel metal1 7038 12172 7038 12172 0 _0311_
rlabel metal1 5152 12954 5152 12954 0 _0312_
rlabel metal2 5566 15300 5566 15300 0 _0313_
rlabel metal1 6744 16082 6744 16082 0 _0314_
rlabel metal2 7222 17068 7222 17068 0 _0315_
rlabel metal1 7498 18156 7498 18156 0 _0316_
rlabel metal2 12742 17748 12742 17748 0 _0317_
rlabel metal1 6762 18394 6762 18394 0 _0318_
rlabel metal1 4922 23120 4922 23120 0 _0319_
rlabel metal1 5796 24922 5796 24922 0 _0320_
rlabel metal1 10626 16558 10626 16558 0 _0321_
rlabel metal1 11362 14416 11362 14416 0 _0322_
rlabel via1 11252 14382 11252 14382 0 _0323_
rlabel metal1 11178 14586 11178 14586 0 _0324_
rlabel via1 10442 18258 10442 18258 0 _0325_
rlabel metal1 10442 18394 10442 18394 0 _0326_
rlabel metal2 12466 18904 12466 18904 0 _0327_
rlabel metal2 2162 21794 2162 21794 0 _0328_
rlabel metal1 2714 21964 2714 21964 0 _0329_
rlabel metal1 7222 29002 7222 29002 0 _0330_
rlabel metal1 6026 12954 6026 12954 0 _0331_
rlabel metal1 7130 15538 7130 15538 0 _0332_
rlabel metal1 7130 15402 7130 15402 0 _0333_
rlabel metal1 11822 14552 11822 14552 0 _0334_
rlabel metal1 8372 15674 8372 15674 0 _0335_
rlabel metal1 8326 19244 8326 19244 0 _0336_
rlabel metal1 14030 16150 14030 16150 0 _0337_
rlabel metal1 2152 24174 2152 24174 0 _0338_
rlabel metal2 1794 26724 1794 26724 0 _0339_
rlabel metal1 7406 14314 7406 14314 0 _0340_
rlabel metal1 9154 14586 9154 14586 0 _0341_
rlabel viali 10258 14994 10258 14994 0 _0342_
rlabel metal1 10994 19482 10994 19482 0 _0343_
rlabel metal2 10534 19924 10534 19924 0 _0344_
rlabel metal1 14260 17850 14260 17850 0 _0345_
rlabel metal2 4922 23460 4922 23460 0 _0346_
rlabel metal1 11316 17306 11316 17306 0 _0347_
rlabel metal1 4876 13498 4876 13498 0 _0348_
rlabel via1 6946 14909 6946 14909 0 _0349_
rlabel metal2 5842 14552 5842 14552 0 _0350_
rlabel metal2 6026 14042 6026 14042 0 _0351_
rlabel metal1 5980 14042 5980 14042 0 _0352_
rlabel metal1 5934 18734 5934 18734 0 _0353_
rlabel metal1 5750 18802 5750 18802 0 _0354_
rlabel metal1 6532 18666 6532 18666 0 _0355_
rlabel metal1 6946 20570 6946 20570 0 _0356_
rlabel metal1 7406 25398 7406 25398 0 _0357_
rlabel metal1 6762 28118 6762 28118 0 _0358_
rlabel metal1 6854 25874 6854 25874 0 _0359_
rlabel metal1 6716 25466 6716 25466 0 _0360_
rlabel metal1 4600 13906 4600 13906 0 _0361_
rlabel metal1 5014 14042 5014 14042 0 _0362_
rlabel metal1 6118 11866 6118 11866 0 _0363_
rlabel metal1 7314 14926 7314 14926 0 _0364_
rlabel metal1 6624 15130 6624 15130 0 _0365_
rlabel metal2 6486 20468 6486 20468 0 _0366_
rlabel metal1 6900 21658 6900 21658 0 _0367_
rlabel metal1 5612 22066 5612 22066 0 _0368_
rlabel metal2 5658 30464 5658 30464 0 _0369_
rlabel metal1 14904 24174 14904 24174 0 _0370_
rlabel metal2 16238 20502 16238 20502 0 _0371_
rlabel metal1 13662 18326 13662 18326 0 _0372_
rlabel metal2 13018 20128 13018 20128 0 _0373_
rlabel metal1 5428 20910 5428 20910 0 _0374_
rlabel metal1 4784 19346 4784 19346 0 _0375_
rlabel viali 3542 19333 3542 19333 0 _0376_
rlabel metal1 6394 16762 6394 16762 0 _0377_
rlabel metal1 7084 20026 7084 20026 0 _0378_
rlabel metal2 13202 27744 13202 27744 0 _0379_
rlabel metal1 4462 31722 4462 31722 0 _0380_
rlabel metal2 3266 18904 3266 18904 0 _0381_
rlabel metal1 5428 20570 5428 20570 0 _0382_
rlabel metal1 4094 31790 4094 31790 0 _0383_
rlabel metal1 8832 25398 8832 25398 0 _0384_
rlabel metal2 9614 27540 9614 27540 0 _0385_
rlabel metal2 11730 27540 11730 27540 0 _0386_
rlabel metal2 6670 28730 6670 28730 0 _0387_
rlabel metal2 12282 25500 12282 25500 0 _0388_
rlabel metal2 4094 27268 4094 27268 0 _0389_
rlabel metal1 4738 27336 4738 27336 0 _0390_
rlabel metal1 5014 26996 5014 26996 0 _0391_
rlabel metal2 12558 19992 12558 19992 0 _0392_
rlabel metal2 4002 28220 4002 28220 0 _0393_
rlabel metal2 4094 25262 4094 25262 0 _0394_
rlabel metal1 1886 25908 1886 25908 0 _0395_
rlabel metal1 2070 28084 2070 28084 0 _0396_
rlabel metal1 4600 28186 4600 28186 0 _0397_
rlabel metal2 2254 29988 2254 29988 0 _0398_
rlabel metal2 12834 22508 12834 22508 0 _0399_
rlabel metal2 13202 25007 13202 25007 0 _0400_
rlabel metal1 2576 17170 2576 17170 0 _0401_
rlabel metal1 22402 2516 22402 2516 0 _0402_
rlabel metal3 10143 6868 10143 6868 0 _0403_
rlabel metal2 13386 22848 13386 22848 0 _0404_
rlabel metal1 11960 20570 11960 20570 0 _0405_
rlabel metal2 16606 25160 16606 25160 0 _0406_
rlabel metal2 17250 25330 17250 25330 0 _0407_
rlabel metal2 15962 20910 15962 20910 0 _0408_
rlabel metal1 12834 19414 12834 19414 0 _0409_
rlabel metal1 7268 22678 7268 22678 0 _0410_
rlabel metal1 7314 22202 7314 22202 0 _0411_
rlabel metal1 5198 20944 5198 20944 0 _0412_
rlabel metal2 3358 19516 3358 19516 0 _0413_
rlabel metal2 3082 17680 3082 17680 0 _0414_
rlabel metal1 2806 17204 2806 17204 0 _0415_
rlabel metal1 4646 16524 4646 16524 0 _0416_
rlabel metal2 9706 16167 9706 16167 0 _0417_
rlabel metal1 7176 16218 7176 16218 0 _0418_
rlabel metal2 11914 15810 11914 15810 0 _0419_
rlabel metal1 7263 5610 7263 5610 0 cal_lut\[0\]
rlabel metal1 18262 10744 18262 10744 0 cal_lut\[100\]
rlabel metal1 14536 10438 14536 10438 0 cal_lut\[101\]
rlabel metal2 10902 13396 10902 13396 0 cal_lut\[102\]
rlabel metal3 17871 9044 17871 9044 0 cal_lut\[103\]
rlabel metal1 12742 21080 12742 21080 0 cal_lut\[104\]
rlabel metal3 14467 11764 14467 11764 0 cal_lut\[105\]
rlabel metal1 15589 16490 15589 16490 0 cal_lut\[106\]
rlabel metal1 16376 16422 16376 16422 0 cal_lut\[107\]
rlabel metal1 22264 18598 22264 18598 0 cal_lut\[108\]
rlabel metal1 25760 21318 25760 21318 0 cal_lut\[109\]
rlabel metal1 27922 15334 27922 15334 0 cal_lut\[10\]
rlabel metal1 24242 18802 24242 18802 0 cal_lut\[110\]
rlabel metal1 22908 17850 22908 17850 0 cal_lut\[111\]
rlabel metal1 21160 15878 21160 15878 0 cal_lut\[112\]
rlabel metal1 25760 14314 25760 14314 0 cal_lut\[113\]
rlabel via2 21942 15555 21942 15555 0 cal_lut\[114\]
rlabel metal1 27078 21930 27078 21930 0 cal_lut\[115\]
rlabel metal1 25847 17238 25847 17238 0 cal_lut\[116\]
rlabel metal1 25985 12818 25985 12818 0 cal_lut\[117\]
rlabel metal2 20194 4964 20194 4964 0 cal_lut\[118\]
rlabel metal1 26128 9146 26128 9146 0 cal_lut\[119\]
rlabel metal1 25806 9350 25806 9350 0 cal_lut\[11\]
rlabel metal1 24242 7718 24242 7718 0 cal_lut\[120\]
rlabel metal1 26618 6698 26618 6698 0 cal_lut\[121\]
rlabel metal1 25428 10642 25428 10642 0 cal_lut\[122\]
rlabel metal1 24932 13158 24932 13158 0 cal_lut\[123\]
rlabel metal1 27600 10234 27600 10234 0 cal_lut\[124\]
rlabel metal1 26624 4590 26624 4590 0 cal_lut\[125\]
rlabel metal2 21390 10455 21390 10455 0 cal_lut\[126\]
rlabel via1 24973 13226 24973 13226 0 cal_lut\[127\]
rlabel metal2 26266 15232 26266 15232 0 cal_lut\[128\]
rlabel metal1 27170 14314 27170 14314 0 cal_lut\[129\]
rlabel metal2 23138 9690 23138 9690 0 cal_lut\[12\]
rlabel metal1 26388 12138 26388 12138 0 cal_lut\[130\]
rlabel metal1 24559 11798 24559 11798 0 cal_lut\[131\]
rlabel via3 23437 19380 23437 19380 0 cal_lut\[132\]
rlabel metal1 20654 17204 20654 17204 0 cal_lut\[133\]
rlabel metal1 20051 26962 20051 26962 0 cal_lut\[134\]
rlabel metal1 20424 26758 20424 26758 0 cal_lut\[135\]
rlabel metal1 22586 16626 22586 16626 0 cal_lut\[136\]
rlabel metal1 20224 24106 20224 24106 0 cal_lut\[137\]
rlabel metal1 21696 21930 21696 21930 0 cal_lut\[138\]
rlabel metal1 20286 17272 20286 17272 0 cal_lut\[139\]
rlabel metal2 18630 8993 18630 8993 0 cal_lut\[13\]
rlabel metal1 20086 19754 20086 19754 0 cal_lut\[140\]
rlabel metal2 22218 19533 22218 19533 0 cal_lut\[141\]
rlabel via2 21206 14773 21206 14773 0 cal_lut\[142\]
rlabel via2 17986 12597 17986 12597 0 cal_lut\[143\]
rlabel metal1 14480 7854 14480 7854 0 cal_lut\[144\]
rlabel metal1 17751 11118 17751 11118 0 cal_lut\[145\]
rlabel via1 20097 7786 20097 7786 0 cal_lut\[146\]
rlabel metal1 21022 8058 21022 8058 0 cal_lut\[147\]
rlabel metal1 18860 7718 18860 7718 0 cal_lut\[148\]
rlabel metal1 25341 8466 25341 8466 0 cal_lut\[149\]
rlabel metal1 18354 11526 18354 11526 0 cal_lut\[14\]
rlabel via1 25898 8602 25898 8602 0 cal_lut\[150\]
rlabel metal1 22632 1258 22632 1258 0 cal_lut\[151\]
rlabel via1 24881 2346 24881 2346 0 cal_lut\[152\]
rlabel metal1 23230 2312 23230 2312 0 cal_lut\[153\]
rlabel metal2 18584 1428 18584 1428 0 cal_lut\[154\]
rlabel metal1 18400 1190 18400 1190 0 cal_lut\[155\]
rlabel via1 18441 5270 18441 5270 0 cal_lut\[156\]
rlabel metal2 20930 2043 20930 2043 0 cal_lut\[157\]
rlabel via1 20746 1938 20746 1938 0 cal_lut\[158\]
rlabel via1 15773 2006 15773 2006 0 cal_lut\[159\]
rlabel metal2 15318 11679 15318 11679 0 cal_lut\[15\]
rlabel metal1 16606 1802 16606 1802 0 cal_lut\[160\]
rlabel metal1 20194 2040 20194 2040 0 cal_lut\[161\]
rlabel metal1 21206 11186 21206 11186 0 cal_lut\[162\]
rlabel metal1 25668 14042 25668 14042 0 cal_lut\[163\]
rlabel via1 23501 21522 23501 21522 0 cal_lut\[164\]
rlabel metal1 21500 20910 21500 20910 0 cal_lut\[165\]
rlabel metal1 18344 20434 18344 20434 0 cal_lut\[166\]
rlabel metal1 16728 19754 16728 19754 0 cal_lut\[167\]
rlabel metal1 16969 26282 16969 26282 0 cal_lut\[168\]
rlabel metal2 17618 27302 17618 27302 0 cal_lut\[169\]
rlabel metal1 12052 11254 12052 11254 0 cal_lut\[16\]
rlabel metal1 15589 23698 15589 23698 0 cal_lut\[170\]
rlabel metal1 16008 23494 16008 23494 0 cal_lut\[171\]
rlabel metal1 15042 22406 15042 22406 0 cal_lut\[172\]
rlabel metal1 14428 18326 14428 18326 0 cal_lut\[173\]
rlabel metal1 15911 14314 15911 14314 0 cal_lut\[174\]
rlabel metal1 16790 14586 16790 14586 0 cal_lut\[175\]
rlabel metal1 18584 17850 18584 17850 0 cal_lut\[176\]
rlabel metal1 18947 25942 18947 25942 0 cal_lut\[177\]
rlabel metal2 19734 23875 19734 23875 0 cal_lut\[178\]
rlabel metal1 22995 17170 22995 17170 0 cal_lut\[179\]
rlabel metal2 13938 10166 13938 10166 0 cal_lut\[17\]
rlabel metal1 22310 11186 22310 11186 0 cal_lut\[180\]
rlabel metal1 26894 7786 26894 7786 0 cal_lut\[181\]
rlabel metal1 27319 13226 27319 13226 0 cal_lut\[182\]
rlabel metal1 24150 12784 24150 12784 0 cal_lut\[183\]
rlabel metal1 26434 18666 26434 18666 0 cal_lut\[184\]
rlabel metal1 27416 18598 27416 18598 0 cal_lut\[185\]
rlabel metal1 27084 3502 27084 3502 0 cal_lut\[186\]
rlabel metal1 25284 1258 25284 1258 0 cal_lut\[187\]
rlabel metal1 25760 1938 25760 1938 0 cal_lut\[188\]
rlabel metal1 25709 7378 25709 7378 0 cal_lut\[189\]
rlabel metal1 14766 6800 14766 6800 0 cal_lut\[18\]
rlabel metal1 26894 8874 26894 8874 0 cal_lut\[190\]
rlabel metal1 27232 11730 27232 11730 0 cal_lut\[191\]
rlabel metal1 11546 2414 11546 2414 0 cal_lut\[19\]
rlabel metal1 8234 5882 8234 5882 0 cal_lut\[1\]
rlabel metal1 8919 2006 8919 2006 0 cal_lut\[20\]
rlabel metal1 6987 3026 6987 3026 0 cal_lut\[21\]
rlabel metal1 4917 1938 4917 1938 0 cal_lut\[22\]
rlabel metal1 12650 7208 12650 7208 0 cal_lut\[23\]
rlabel metal1 11454 5678 11454 5678 0 cal_lut\[24\]
rlabel via1 13110 2414 13110 2414 0 cal_lut\[25\]
rlabel metal2 5198 4760 5198 4760 0 cal_lut\[26\]
rlabel metal1 12834 3468 12834 3468 0 cal_lut\[27\]
rlabel metal2 13018 6749 13018 6749 0 cal_lut\[28\]
rlabel metal1 14950 4488 14950 4488 0 cal_lut\[29\]
rlabel metal2 6854 4607 6854 4607 0 cal_lut\[2\]
rlabel metal1 13662 6358 13662 6358 0 cal_lut\[30\]
rlabel metal1 16238 7956 16238 7956 0 cal_lut\[31\]
rlabel metal1 11254 8534 11254 8534 0 cal_lut\[32\]
rlabel metal1 12788 8602 12788 8602 0 cal_lut\[33\]
rlabel metal1 12972 14042 12972 14042 0 cal_lut\[34\]
rlabel metal1 13340 18598 13340 18598 0 cal_lut\[35\]
rlabel metal2 15502 19312 15502 19312 0 cal_lut\[36\]
rlabel metal1 17480 20774 17480 20774 0 cal_lut\[37\]
rlabel metal2 13846 15198 13846 15198 0 cal_lut\[38\]
rlabel metal1 17066 15504 17066 15504 0 cal_lut\[39\]
rlabel metal1 7125 6698 7125 6698 0 cal_lut\[3\]
rlabel metal1 14060 15062 14060 15062 0 cal_lut\[40\]
rlabel metal2 21022 14909 21022 14909 0 cal_lut\[41\]
rlabel metal1 23230 15878 23230 15878 0 cal_lut\[42\]
rlabel metal2 26450 16592 26450 16592 0 cal_lut\[43\]
rlabel metal1 27968 17510 27968 17510 0 cal_lut\[44\]
rlabel via1 24145 22678 24145 22678 0 cal_lut\[45\]
rlabel metal1 24686 21930 24686 21930 0 cal_lut\[46\]
rlabel via1 20373 21522 20373 21522 0 cal_lut\[47\]
rlabel metal1 20184 22610 20184 22610 0 cal_lut\[48\]
rlabel metal1 17751 23018 17751 23018 0 cal_lut\[49\]
rlabel metal1 8873 7446 8873 7446 0 cal_lut\[4\]
rlabel metal1 18400 22950 18400 22950 0 cal_lut\[50\]
rlabel metal1 18998 21862 18998 21862 0 cal_lut\[51\]
rlabel metal1 9885 21590 9885 21590 0 cal_lut\[52\]
rlabel metal1 13928 19346 13928 19346 0 cal_lut\[53\]
rlabel metal1 18614 17578 18614 17578 0 cal_lut\[54\]
rlabel via1 24881 16490 24881 16490 0 cal_lut\[55\]
rlabel metal1 22995 14314 22995 14314 0 cal_lut\[56\]
rlabel via1 21109 8874 21109 8874 0 cal_lut\[57\]
rlabel metal2 20470 6868 20470 6868 0 cal_lut\[58\]
rlabel via1 17613 6290 17613 6290 0 cal_lut\[59\]
rlabel metal1 10120 10574 10120 10574 0 cal_lut\[5\]
rlabel metal1 17383 2006 17383 2006 0 cal_lut\[60\]
rlabel metal1 15221 2346 15221 2346 0 cal_lut\[61\]
rlabel metal2 21022 2108 21022 2108 0 cal_lut\[62\]
rlabel metal1 15686 3366 15686 3366 0 cal_lut\[63\]
rlabel metal1 13248 3162 13248 3162 0 cal_lut\[64\]
rlabel metal1 13151 2006 13151 2006 0 cal_lut\[65\]
rlabel metal1 13984 2074 13984 2074 0 cal_lut\[66\]
rlabel metal1 13018 3400 13018 3400 0 cal_lut\[67\]
rlabel metal1 13933 5270 13933 5270 0 cal_lut\[68\]
rlabel metal1 14628 3026 14628 3026 0 cal_lut\[69\]
rlabel metal2 20792 13124 20792 13124 0 cal_lut\[6\]
rlabel metal1 14858 1292 14858 1292 0 cal_lut\[70\]
rlabel metal1 14766 4794 14766 4794 0 cal_lut\[71\]
rlabel metal1 17199 4590 17199 4590 0 cal_lut\[72\]
rlabel metal2 17710 2587 17710 2587 0 cal_lut\[73\]
rlabel metal2 11730 3502 11730 3502 0 cal_lut\[74\]
rlabel metal1 13386 2856 13386 2856 0 cal_lut\[75\]
rlabel metal1 12466 7344 12466 7344 0 cal_lut\[76\]
rlabel metal1 15134 8908 15134 8908 0 cal_lut\[77\]
rlabel metal1 19688 15334 19688 15334 0 cal_lut\[78\]
rlabel metal1 20792 15674 20792 15674 0 cal_lut\[79\]
rlabel metal1 22586 13158 22586 13158 0 cal_lut\[7\]
rlabel metal1 23593 18326 23593 18326 0 cal_lut\[80\]
rlabel via2 24426 18037 24426 18037 0 cal_lut\[81\]
rlabel metal1 25208 20230 25208 20230 0 cal_lut\[82\]
rlabel metal1 26031 15062 26031 15062 0 cal_lut\[83\]
rlabel metal1 23041 1326 23041 1326 0 cal_lut\[84\]
rlabel metal2 23782 1088 23782 1088 0 cal_lut\[85\]
rlabel metal2 20562 3808 20562 3808 0 cal_lut\[86\]
rlabel metal1 19734 1326 19734 1326 0 cal_lut\[87\]
rlabel metal1 20838 3162 20838 3162 0 cal_lut\[88\]
rlabel metal2 21574 6868 21574 6868 0 cal_lut\[89\]
rlabel metal1 25806 15334 25806 15334 0 cal_lut\[8\]
rlabel metal1 25054 6358 25054 6358 0 cal_lut\[90\]
rlabel metal1 26496 6426 26496 6426 0 cal_lut\[91\]
rlabel metal2 25990 7140 25990 7140 0 cal_lut\[92\]
rlabel metal1 23904 2006 23904 2006 0 cal_lut\[93\]
rlabel metal1 23092 2006 23092 2006 0 cal_lut\[94\]
rlabel metal1 22673 1938 22673 1938 0 cal_lut\[95\]
rlabel metal1 23368 2074 23368 2074 0 cal_lut\[96\]
rlabel metal2 20286 6460 20286 6460 0 cal_lut\[97\]
rlabel metal1 20925 5610 20925 5610 0 cal_lut\[98\]
rlabel metal1 21528 5882 21528 5882 0 cal_lut\[99\]
rlabel metal2 26634 14552 26634 14552 0 cal_lut\[9\]
rlabel metal2 2622 25704 2622 25704 0 clknet_0__0390_
rlabel metal2 2622 13396 2622 13396 0 clknet_0_io_in[0]
rlabel metal1 1656 32402 1656 32402 0 clknet_0_net57
rlabel metal1 1702 30804 1702 30804 0 clknet_0_temp1.dcdel_capnode_notouch_
rlabel metal1 2576 28050 2576 28050 0 clknet_0_temp1.i_precharge_n
rlabel metal2 5014 26928 5014 26928 0 clknet_1_0__leaf__0390_
rlabel metal2 1610 6562 1610 6562 0 clknet_1_0__leaf_io_in[0]
rlabel metal2 2714 25194 2714 25194 0 clknet_1_0__leaf_net57
rlabel metal1 15778 31722 15778 31722 0 clknet_1_0__leaf_temp1.dcdel_capnode_notouch_
rlabel metal2 3358 32062 3358 32062 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal1 2070 29070 2070 29070 0 clknet_1_1__leaf__0390_
rlabel metal2 1886 19108 1886 19108 0 clknet_1_1__leaf_io_in[0]
rlabel metal1 5934 32470 5934 32470 0 clknet_1_1__leaf_net57
rlabel metal1 10350 32402 10350 32402 0 clknet_1_1__leaf_temp1.dcdel_capnode_notouch_
rlabel metal1 4140 28186 4140 28186 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal2 5382 969 5382 969 0 ctr\[0\]
rlabel metal1 4600 17170 4600 17170 0 ctr\[10\]
rlabel metal2 5658 16218 5658 16218 0 ctr\[11\]
rlabel metal1 6072 16082 6072 16082 0 ctr\[12\]
rlabel metal1 13018 25330 13018 25330 0 ctr\[1\]
rlabel metal1 10856 1258 10856 1258 0 ctr\[2\]
rlabel via2 3358 2635 3358 2635 0 ctr\[3\]
rlabel metal1 16882 24174 16882 24174 0 ctr\[4\]
rlabel metal2 15594 19584 15594 19584 0 ctr\[5\]
rlabel metal1 13110 24820 13110 24820 0 ctr\[6\]
rlabel metal2 7406 14450 7406 14450 0 ctr\[7\]
rlabel via2 7498 17629 7498 17629 0 ctr\[8\]
rlabel metal2 6946 16031 6946 16031 0 ctr\[9\]
rlabel metal1 13708 17510 13708 17510 0 dbg3\[0\]
rlabel metal1 13018 17646 13018 17646 0 dbg3\[1\]
rlabel metal2 9982 17986 9982 17986 0 dbg3\[2\]
rlabel metal2 13478 17884 13478 17884 0 dbg3\[3\]
rlabel metal3 6417 26316 6417 26316 0 dbg3\[4\]
rlabel metal1 12098 17136 12098 17136 0 dbg3\[5\]
rlabel via2 8234 11067 8234 11067 0 dec1.i_ones
rlabel metal3 1602 1700 1602 1700 0 io_in[0]
rlabel metal3 820 3740 820 3740 0 io_in[1]
rlabel metal3 1050 5780 1050 5780 0 io_in[2]
rlabel metal3 636 7820 636 7820 0 io_in[3]
rlabel metal3 590 9860 590 9860 0 io_in[4]
rlabel metal3 544 11900 544 11900 0 io_in[5]
rlabel metal3 452 13940 452 13940 0 io_in[6]
rlabel metal3 498 15980 498 15980 0 io_in[7]
rlabel metal2 3910 19975 3910 19975 0 io_out[0]
rlabel metal2 4140 20060 4140 20060 0 io_out[1]
rlabel metal3 1142 22100 1142 22100 0 io_out[2]
rlabel metal3 590 24140 590 24140 0 io_out[3]
rlabel metal1 4784 24310 4784 24310 0 io_out[4]
rlabel metal2 6578 26792 6578 26792 0 io_out[5]
rlabel via2 4002 30277 4002 30277 0 io_out[6]
rlabel metal3 1556 32300 1556 32300 0 io_out[7]
rlabel metal2 17710 25840 17710 25840 0 net1
rlabel metal1 11132 31790 11132 31790 0 net10
rlabel metal1 10442 31858 10442 31858 0 net11
rlabel metal1 13800 29614 13800 29614 0 net12
rlabel metal2 14398 30464 14398 30464 0 net13
rlabel metal1 7958 1802 7958 1802 0 net14
rlabel metal1 2714 5236 2714 5236 0 net15
rlabel metal1 14812 2482 14812 2482 0 net16
rlabel metal2 13294 5508 13294 5508 0 net17
rlabel metal2 14306 11152 14306 11152 0 net18
rlabel metal1 1978 5270 1978 5270 0 net19
rlabel metal2 2806 6732 2806 6732 0 net2
rlabel metal1 16974 1802 16974 1802 0 net20
rlabel metal1 16974 1326 16974 1326 0 net21
rlabel metal1 24288 2482 24288 2482 0 net22
rlabel metal2 27002 1904 27002 1904 0 net23
rlabel metal2 25254 5406 25254 5406 0 net24
rlabel metal1 17572 5542 17572 5542 0 net25
rlabel metal1 26864 7854 26864 7854 0 net26
rlabel metal1 25806 14994 25806 14994 0 net27
rlabel metal1 19688 14926 19688 14926 0 net28
rlabel metal1 14904 16626 14904 16626 0 net29
rlabel metal2 4278 6120 4278 6120 0 net3
rlabel metal2 12926 22814 12926 22814 0 net30
rlabel metal2 16790 20400 16790 20400 0 net31
rlabel metal1 22034 20468 22034 20468 0 net32
rlabel metal1 21850 16082 21850 16082 0 net33
rlabel metal2 19734 15317 19734 15317 0 net34
rlabel metal1 22034 22644 22034 22644 0 net35
rlabel metal1 20884 24242 20884 24242 0 net36
rlabel metal2 21850 26656 21850 26656 0 net37
rlabel metal2 16882 11407 16882 11407 0 net38
rlabel metal1 13846 29240 13846 29240 0 net39
rlabel metal2 1794 10914 1794 10914 0 net4
rlabel metal1 2277 23494 2277 23494 0 net40
rlabel viali 4002 24785 4002 24785 0 net41
rlabel metal1 6831 31994 6831 31994 0 net42
rlabel metal1 15134 32334 15134 32334 0 net43
rlabel metal1 11040 29002 11040 29002 0 net44
rlabel metal2 15134 31994 15134 31994 0 net45
rlabel metal1 5842 32198 5842 32198 0 net46
rlabel metal1 8234 26996 8234 26996 0 net47
rlabel metal1 15778 31858 15778 31858 0 net48
rlabel metal2 15778 30566 15778 30566 0 net49
rlabel metal2 1886 13328 1886 13328 0 net5
rlabel metal1 7222 32266 7222 32266 0 net50
rlabel metal1 14306 31722 14306 31722 0 net51
rlabel metal2 14490 31110 14490 31110 0 net52
rlabel metal2 12558 32198 12558 32198 0 net53
rlabel metal1 10626 31926 10626 31926 0 net54
rlabel metal2 18354 27200 18354 27200 0 net55
rlabel metal2 14398 27132 14398 27132 0 net56
rlabel metal1 1702 29648 1702 29648 0 net57
rlabel metal2 2162 27302 2162 27302 0 net58
rlabel metal1 2001 24718 2001 24718 0 net59
rlabel metal2 2714 17442 2714 17442 0 net6
rlabel metal1 4278 31824 4278 31824 0 net60
rlabel metal2 1702 17442 1702 17442 0 net7
rlabel metal2 14214 29308 14214 29308 0 net8
rlabel metal2 12650 30906 12650 30906 0 net9
rlabel metal2 8234 26588 8234 26588 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal1 7406 26928 7406 26928 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal1 8510 25466 8510 25466 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal1 7636 28050 7636 28050 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal1 10672 27506 10672 27506 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 8970 26962 8970 26962 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal1 13110 25874 13110 25874 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal1 13202 28492 13202 28492 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal1 13110 25738 13110 25738 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 5198 31790 5198 31790 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal1 7912 31790 7912 31790 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal1 5566 31926 5566 31926 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 12006 29410 12006 29410 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal2 11914 26452 11914 26452 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal2 12742 25228 12742 25228 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal1 13892 26962 13892 26962 0 temp1.dac.vdac_single.en_pupd
rlabel metal2 5198 32470 5198 32470 0 temp1.dac_vout_notouch_
rlabel metal1 4692 30702 4692 30702 0 temp1.dcdel_capnode_notouch_
rlabel metal1 6440 29274 6440 29274 0 temp1.i_precharge_n
rlabel metal1 1610 26826 1610 26826 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>
